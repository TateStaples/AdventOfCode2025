module day8_opt_a (
    x0_value,
    edge_j,
    edge_i,
    n_nodes,
    clear,
    clock,
    edge_last,
    edge_valid,
    edge_phase,
    x0_last,
    x0_valid,
    load,
    x0_ready,
    edge_ready,
    done_,
    part1_result,
    part2_result,
    state
);

    input [31:0] x0_value;
    input [7:0] edge_j;
    input [7:0] edge_i;
    input [7:0] n_nodes;
    input clear;
    input clock;
    input edge_last;
    input edge_valid;
    input edge_phase;
    input x0_last;
    input x0_valid;
    input load;
    output x0_ready;
    output edge_ready;
    output done_;
    output [63:0] part1_result;
    output [63:0] part2_result;
    output [2:0] state;

    wire [63:0] _4700;
    reg [31:0] _4708;
    wire [31:0] _4707;
    wire [63:0] _4709;
    wire [7:0] _818;
    wire _819;
    wire _820;
    wire [31:0] _824;
    wire [31:0] _826;
    wire [31:0] _2;
    reg [31:0] _823;
    wire [7:0] _827;
    wire _828;
    wire _829;
    wire [31:0] _833;
    wire [31:0] _835;
    wire [31:0] _3;
    reg [31:0] _832;
    wire [7:0] _836;
    wire _837;
    wire _838;
    wire [31:0] _842;
    wire [31:0] _844;
    wire [31:0] _4;
    reg [31:0] _841;
    wire [7:0] _845;
    wire _846;
    wire _847;
    wire [31:0] _851;
    wire [31:0] _853;
    wire [31:0] _5;
    reg [31:0] _850;
    wire [7:0] _854;
    wire _855;
    wire _856;
    wire [31:0] _860;
    wire [31:0] _862;
    wire [31:0] _6;
    reg [31:0] _859;
    wire [7:0] _863;
    wire _864;
    wire _865;
    wire [31:0] _869;
    wire [31:0] _871;
    wire [31:0] _7;
    reg [31:0] _868;
    wire [7:0] _872;
    wire _873;
    wire _874;
    wire [31:0] _878;
    wire [31:0] _880;
    wire [31:0] _8;
    reg [31:0] _877;
    wire [7:0] _881;
    wire _882;
    wire _883;
    wire [31:0] _887;
    wire [31:0] _889;
    wire [31:0] _9;
    reg [31:0] _886;
    wire [7:0] _890;
    wire _891;
    wire _892;
    wire [31:0] _896;
    wire [31:0] _898;
    wire [31:0] _10;
    reg [31:0] _895;
    wire [7:0] _899;
    wire _900;
    wire _901;
    wire [31:0] _905;
    wire [31:0] _907;
    wire [31:0] _11;
    reg [31:0] _904;
    wire [7:0] _908;
    wire _909;
    wire _910;
    wire [31:0] _914;
    wire [31:0] _916;
    wire [31:0] _12;
    reg [31:0] _913;
    wire [7:0] _917;
    wire _918;
    wire _919;
    wire [31:0] _923;
    wire [31:0] _925;
    wire [31:0] _13;
    reg [31:0] _922;
    wire [7:0] _926;
    wire _927;
    wire _928;
    wire [31:0] _932;
    wire [31:0] _934;
    wire [31:0] _14;
    reg [31:0] _931;
    wire [7:0] _935;
    wire _936;
    wire _937;
    wire [31:0] _941;
    wire [31:0] _943;
    wire [31:0] _15;
    reg [31:0] _940;
    wire [7:0] _944;
    wire _945;
    wire _946;
    wire [31:0] _950;
    wire [31:0] _952;
    wire [31:0] _16;
    reg [31:0] _949;
    wire [7:0] _953;
    wire _954;
    wire _955;
    wire [31:0] _959;
    wire [31:0] _961;
    wire [31:0] _17;
    reg [31:0] _958;
    wire [7:0] _962;
    wire _963;
    wire _964;
    wire [31:0] _968;
    wire [31:0] _970;
    wire [31:0] _18;
    reg [31:0] _967;
    wire [7:0] _971;
    wire _972;
    wire _973;
    wire [31:0] _977;
    wire [31:0] _979;
    wire [31:0] _19;
    reg [31:0] _976;
    wire [7:0] _980;
    wire _981;
    wire _982;
    wire [31:0] _986;
    wire [31:0] _988;
    wire [31:0] _20;
    reg [31:0] _985;
    wire [7:0] _989;
    wire _990;
    wire _991;
    wire [31:0] _995;
    wire [31:0] _997;
    wire [31:0] _21;
    reg [31:0] _994;
    wire [7:0] _998;
    wire _999;
    wire _1000;
    wire [31:0] _1004;
    wire [31:0] _1006;
    wire [31:0] _22;
    reg [31:0] _1003;
    wire [7:0] _1007;
    wire _1008;
    wire _1009;
    wire [31:0] _1013;
    wire [31:0] _1015;
    wire [31:0] _23;
    reg [31:0] _1012;
    wire [7:0] _1016;
    wire _1017;
    wire _1018;
    wire [31:0] _1022;
    wire [31:0] _1024;
    wire [31:0] _24;
    reg [31:0] _1021;
    wire [7:0] _1025;
    wire _1026;
    wire _1027;
    wire [31:0] _1031;
    wire [31:0] _1033;
    wire [31:0] _25;
    reg [31:0] _1030;
    wire [7:0] _1034;
    wire _1035;
    wire _1036;
    wire [31:0] _1040;
    wire [31:0] _1042;
    wire [31:0] _26;
    reg [31:0] _1039;
    wire [7:0] _1043;
    wire _1044;
    wire _1045;
    wire [31:0] _1049;
    wire [31:0] _1051;
    wire [31:0] _27;
    reg [31:0] _1048;
    wire [7:0] _1052;
    wire _1053;
    wire _1054;
    wire [31:0] _1058;
    wire [31:0] _1060;
    wire [31:0] _28;
    reg [31:0] _1057;
    wire [7:0] _1061;
    wire _1062;
    wire _1063;
    wire [31:0] _1067;
    wire [31:0] _1069;
    wire [31:0] _29;
    reg [31:0] _1066;
    wire [7:0] _1070;
    wire _1071;
    wire _1072;
    wire [31:0] _1076;
    wire [31:0] _1078;
    wire [31:0] _30;
    reg [31:0] _1075;
    wire [7:0] _1079;
    wire _1080;
    wire _1081;
    wire [31:0] _1085;
    wire [31:0] _1087;
    wire [31:0] _31;
    reg [31:0] _1084;
    wire [7:0] _1088;
    wire _1089;
    wire _1090;
    wire [31:0] _1094;
    wire [31:0] _1096;
    wire [31:0] _32;
    reg [31:0] _1093;
    wire [7:0] _1097;
    wire _1098;
    wire _1099;
    wire [31:0] _1103;
    wire [31:0] _1105;
    wire [31:0] _33;
    reg [31:0] _1102;
    wire [7:0] _1106;
    wire _1107;
    wire _1108;
    wire [31:0] _1112;
    wire [31:0] _1114;
    wire [31:0] _34;
    reg [31:0] _1111;
    wire [7:0] _1115;
    wire _1116;
    wire _1117;
    wire [31:0] _1121;
    wire [31:0] _1123;
    wire [31:0] _35;
    reg [31:0] _1120;
    wire [7:0] _1124;
    wire _1125;
    wire _1126;
    wire [31:0] _1130;
    wire [31:0] _1132;
    wire [31:0] _36;
    reg [31:0] _1129;
    wire [7:0] _1133;
    wire _1134;
    wire _1135;
    wire [31:0] _1139;
    wire [31:0] _1141;
    wire [31:0] _37;
    reg [31:0] _1138;
    wire [7:0] _1142;
    wire _1143;
    wire _1144;
    wire [31:0] _1148;
    wire [31:0] _1150;
    wire [31:0] _38;
    reg [31:0] _1147;
    wire [7:0] _1151;
    wire _1152;
    wire _1153;
    wire [31:0] _1157;
    wire [31:0] _1159;
    wire [31:0] _39;
    reg [31:0] _1156;
    wire [7:0] _1160;
    wire _1161;
    wire _1162;
    wire [31:0] _1166;
    wire [31:0] _1168;
    wire [31:0] _40;
    reg [31:0] _1165;
    wire [7:0] _1169;
    wire _1170;
    wire _1171;
    wire [31:0] _1175;
    wire [31:0] _1177;
    wire [31:0] _41;
    reg [31:0] _1174;
    wire [7:0] _1178;
    wire _1179;
    wire _1180;
    wire [31:0] _1184;
    wire [31:0] _1186;
    wire [31:0] _42;
    reg [31:0] _1183;
    wire [7:0] _1187;
    wire _1188;
    wire _1189;
    wire [31:0] _1193;
    wire [31:0] _1195;
    wire [31:0] _43;
    reg [31:0] _1192;
    wire [7:0] _1196;
    wire _1197;
    wire _1198;
    wire [31:0] _1202;
    wire [31:0] _1204;
    wire [31:0] _44;
    reg [31:0] _1201;
    wire [7:0] _1205;
    wire _1206;
    wire _1207;
    wire [31:0] _1211;
    wire [31:0] _1213;
    wire [31:0] _45;
    reg [31:0] _1210;
    wire [7:0] _1214;
    wire _1215;
    wire _1216;
    wire [31:0] _1220;
    wire [31:0] _1222;
    wire [31:0] _46;
    reg [31:0] _1219;
    wire [7:0] _1223;
    wire _1224;
    wire _1225;
    wire [31:0] _1229;
    wire [31:0] _1231;
    wire [31:0] _47;
    reg [31:0] _1228;
    wire [7:0] _1232;
    wire _1233;
    wire _1234;
    wire [31:0] _1238;
    wire [31:0] _1240;
    wire [31:0] _48;
    reg [31:0] _1237;
    wire [7:0] _1241;
    wire _1242;
    wire _1243;
    wire [31:0] _1247;
    wire [31:0] _1249;
    wire [31:0] _49;
    reg [31:0] _1246;
    wire [7:0] _1250;
    wire _1251;
    wire _1252;
    wire [31:0] _1256;
    wire [31:0] _1258;
    wire [31:0] _50;
    reg [31:0] _1255;
    wire [7:0] _1259;
    wire _1260;
    wire _1261;
    wire [31:0] _1265;
    wire [31:0] _1267;
    wire [31:0] _51;
    reg [31:0] _1264;
    wire [7:0] _1268;
    wire _1269;
    wire _1270;
    wire [31:0] _1274;
    wire [31:0] _1276;
    wire [31:0] _52;
    reg [31:0] _1273;
    wire [7:0] _1277;
    wire _1278;
    wire _1279;
    wire [31:0] _1283;
    wire [31:0] _1285;
    wire [31:0] _53;
    reg [31:0] _1282;
    wire [7:0] _1286;
    wire _1287;
    wire _1288;
    wire [31:0] _1292;
    wire [31:0] _1294;
    wire [31:0] _54;
    reg [31:0] _1291;
    wire [7:0] _1295;
    wire _1296;
    wire _1297;
    wire [31:0] _1301;
    wire [31:0] _1303;
    wire [31:0] _55;
    reg [31:0] _1300;
    wire [7:0] _1304;
    wire _1305;
    wire _1306;
    wire [31:0] _1310;
    wire [31:0] _1312;
    wire [31:0] _56;
    reg [31:0] _1309;
    wire [7:0] _1313;
    wire _1314;
    wire _1315;
    wire [31:0] _1319;
    wire [31:0] _1321;
    wire [31:0] _57;
    reg [31:0] _1318;
    wire [7:0] _1322;
    wire _1323;
    wire _1324;
    wire [31:0] _1328;
    wire [31:0] _1330;
    wire [31:0] _58;
    reg [31:0] _1327;
    wire [7:0] _1331;
    wire _1332;
    wire _1333;
    wire [31:0] _1337;
    wire [31:0] _1339;
    wire [31:0] _59;
    reg [31:0] _1336;
    wire [7:0] _1340;
    wire _1341;
    wire _1342;
    wire [31:0] _1346;
    wire [31:0] _1348;
    wire [31:0] _60;
    reg [31:0] _1345;
    wire [7:0] _1349;
    wire _1350;
    wire _1351;
    wire [31:0] _1355;
    wire [31:0] _1357;
    wire [31:0] _61;
    reg [31:0] _1354;
    wire [7:0] _1358;
    wire _1359;
    wire _1360;
    wire [31:0] _1364;
    wire [31:0] _1366;
    wire [31:0] _62;
    reg [31:0] _1363;
    wire [7:0] _1367;
    wire _1368;
    wire _1369;
    wire [31:0] _1373;
    wire [31:0] _1375;
    wire [31:0] _63;
    reg [31:0] _1372;
    wire [7:0] _1376;
    wire _1377;
    wire _1378;
    wire [31:0] _1382;
    wire [31:0] _1384;
    wire [31:0] _64;
    reg [31:0] _1381;
    wire [7:0] _1385;
    wire _1386;
    wire _1387;
    wire [31:0] _1391;
    wire [31:0] _1393;
    wire [31:0] _65;
    reg [31:0] _1390;
    wire [7:0] _1394;
    wire _1395;
    wire _1396;
    wire [31:0] _1400;
    wire [31:0] _1402;
    wire [31:0] _66;
    reg [31:0] _1399;
    wire [7:0] _1403;
    wire _1404;
    wire _1405;
    wire [31:0] _1409;
    wire [31:0] _1411;
    wire [31:0] _67;
    reg [31:0] _1408;
    wire [7:0] _1412;
    wire _1413;
    wire _1414;
    wire [31:0] _1418;
    wire [31:0] _1420;
    wire [31:0] _68;
    reg [31:0] _1417;
    wire [7:0] _1421;
    wire _1422;
    wire _1423;
    wire [31:0] _1427;
    wire [31:0] _1429;
    wire [31:0] _69;
    reg [31:0] _1426;
    wire [7:0] _1430;
    wire _1431;
    wire _1432;
    wire [31:0] _1436;
    wire [31:0] _1438;
    wire [31:0] _70;
    reg [31:0] _1435;
    wire [7:0] _1439;
    wire _1440;
    wire _1441;
    wire [31:0] _1445;
    wire [31:0] _1447;
    wire [31:0] _71;
    reg [31:0] _1444;
    wire [7:0] _1448;
    wire _1449;
    wire _1450;
    wire [31:0] _1454;
    wire [31:0] _1456;
    wire [31:0] _72;
    reg [31:0] _1453;
    wire [7:0] _1457;
    wire _1458;
    wire _1459;
    wire [31:0] _1463;
    wire [31:0] _1465;
    wire [31:0] _73;
    reg [31:0] _1462;
    wire [7:0] _1466;
    wire _1467;
    wire _1468;
    wire [31:0] _1472;
    wire [31:0] _1474;
    wire [31:0] _74;
    reg [31:0] _1471;
    wire [7:0] _1475;
    wire _1476;
    wire _1477;
    wire [31:0] _1481;
    wire [31:0] _1483;
    wire [31:0] _75;
    reg [31:0] _1480;
    wire [7:0] _1484;
    wire _1485;
    wire _1486;
    wire [31:0] _1490;
    wire [31:0] _1492;
    wire [31:0] _76;
    reg [31:0] _1489;
    wire [7:0] _1493;
    wire _1494;
    wire _1495;
    wire [31:0] _1499;
    wire [31:0] _1501;
    wire [31:0] _77;
    reg [31:0] _1498;
    wire [7:0] _1502;
    wire _1503;
    wire _1504;
    wire [31:0] _1508;
    wire [31:0] _1510;
    wire [31:0] _78;
    reg [31:0] _1507;
    wire [7:0] _1511;
    wire _1512;
    wire _1513;
    wire [31:0] _1517;
    wire [31:0] _1519;
    wire [31:0] _79;
    reg [31:0] _1516;
    wire [7:0] _1520;
    wire _1521;
    wire _1522;
    wire [31:0] _1526;
    wire [31:0] _1528;
    wire [31:0] _80;
    reg [31:0] _1525;
    wire [7:0] _1529;
    wire _1530;
    wire _1531;
    wire [31:0] _1535;
    wire [31:0] _1537;
    wire [31:0] _81;
    reg [31:0] _1534;
    wire [7:0] _1538;
    wire _1539;
    wire _1540;
    wire [31:0] _1544;
    wire [31:0] _1546;
    wire [31:0] _82;
    reg [31:0] _1543;
    wire [7:0] _1547;
    wire _1548;
    wire _1549;
    wire [31:0] _1553;
    wire [31:0] _1555;
    wire [31:0] _83;
    reg [31:0] _1552;
    wire [7:0] _1556;
    wire _1557;
    wire _1558;
    wire [31:0] _1562;
    wire [31:0] _1564;
    wire [31:0] _84;
    reg [31:0] _1561;
    wire [7:0] _1565;
    wire _1566;
    wire _1567;
    wire [31:0] _1571;
    wire [31:0] _1573;
    wire [31:0] _85;
    reg [31:0] _1570;
    wire [7:0] _1574;
    wire _1575;
    wire _1576;
    wire [31:0] _1580;
    wire [31:0] _1582;
    wire [31:0] _86;
    reg [31:0] _1579;
    wire [7:0] _1583;
    wire _1584;
    wire _1585;
    wire [31:0] _1589;
    wire [31:0] _1591;
    wire [31:0] _87;
    reg [31:0] _1588;
    wire [7:0] _1592;
    wire _1593;
    wire _1594;
    wire [31:0] _1598;
    wire [31:0] _1600;
    wire [31:0] _88;
    reg [31:0] _1597;
    wire [7:0] _1601;
    wire _1602;
    wire _1603;
    wire [31:0] _1607;
    wire [31:0] _1609;
    wire [31:0] _89;
    reg [31:0] _1606;
    wire [7:0] _1610;
    wire _1611;
    wire _1612;
    wire [31:0] _1616;
    wire [31:0] _1618;
    wire [31:0] _90;
    reg [31:0] _1615;
    wire [7:0] _1619;
    wire _1620;
    wire _1621;
    wire [31:0] _1625;
    wire [31:0] _1627;
    wire [31:0] _91;
    reg [31:0] _1624;
    wire [7:0] _1628;
    wire _1629;
    wire _1630;
    wire [31:0] _1634;
    wire [31:0] _1636;
    wire [31:0] _92;
    reg [31:0] _1633;
    wire [7:0] _1637;
    wire _1638;
    wire _1639;
    wire [31:0] _1643;
    wire [31:0] _1645;
    wire [31:0] _93;
    reg [31:0] _1642;
    wire [7:0] _1646;
    wire _1647;
    wire _1648;
    wire [31:0] _1652;
    wire [31:0] _1654;
    wire [31:0] _94;
    reg [31:0] _1651;
    wire [7:0] _1655;
    wire _1656;
    wire _1657;
    wire [31:0] _1661;
    wire [31:0] _1663;
    wire [31:0] _95;
    reg [31:0] _1660;
    wire [7:0] _1664;
    wire _1665;
    wire _1666;
    wire [31:0] _1670;
    wire [31:0] _1672;
    wire [31:0] _96;
    reg [31:0] _1669;
    wire [7:0] _1673;
    wire _1674;
    wire _1675;
    wire [31:0] _1679;
    wire [31:0] _1681;
    wire [31:0] _97;
    reg [31:0] _1678;
    wire [7:0] _1682;
    wire _1683;
    wire _1684;
    wire [31:0] _1688;
    wire [31:0] _1690;
    wire [31:0] _98;
    reg [31:0] _1687;
    wire [7:0] _1691;
    wire _1692;
    wire _1693;
    wire [31:0] _1697;
    wire [31:0] _1699;
    wire [31:0] _99;
    reg [31:0] _1696;
    wire [7:0] _1700;
    wire _1701;
    wire _1702;
    wire [31:0] _1706;
    wire [31:0] _1708;
    wire [31:0] _100;
    reg [31:0] _1705;
    wire [7:0] _1709;
    wire _1710;
    wire _1711;
    wire [31:0] _1715;
    wire [31:0] _1717;
    wire [31:0] _101;
    reg [31:0] _1714;
    wire [7:0] _1718;
    wire _1719;
    wire _1720;
    wire [31:0] _1724;
    wire [31:0] _1726;
    wire [31:0] _102;
    reg [31:0] _1723;
    wire [7:0] _1727;
    wire _1728;
    wire _1729;
    wire [31:0] _1733;
    wire [31:0] _1735;
    wire [31:0] _103;
    reg [31:0] _1732;
    wire [7:0] _1736;
    wire _1737;
    wire _1738;
    wire [31:0] _1742;
    wire [31:0] _1744;
    wire [31:0] _104;
    reg [31:0] _1741;
    wire [7:0] _1745;
    wire _1746;
    wire _1747;
    wire [31:0] _1751;
    wire [31:0] _1753;
    wire [31:0] _105;
    reg [31:0] _1750;
    wire [7:0] _1754;
    wire _1755;
    wire _1756;
    wire [31:0] _1760;
    wire [31:0] _1762;
    wire [31:0] _106;
    reg [31:0] _1759;
    wire [7:0] _1763;
    wire _1764;
    wire _1765;
    wire [31:0] _1769;
    wire [31:0] _1771;
    wire [31:0] _107;
    reg [31:0] _1768;
    wire [7:0] _1772;
    wire _1773;
    wire _1774;
    wire [31:0] _1778;
    wire [31:0] _1780;
    wire [31:0] _108;
    reg [31:0] _1777;
    wire [7:0] _1781;
    wire _1782;
    wire _1783;
    wire [31:0] _1787;
    wire [31:0] _1789;
    wire [31:0] _109;
    reg [31:0] _1786;
    wire [7:0] _1790;
    wire _1791;
    wire _1792;
    wire [31:0] _1796;
    wire [31:0] _1798;
    wire [31:0] _110;
    reg [31:0] _1795;
    wire [7:0] _1799;
    wire _1800;
    wire _1801;
    wire [31:0] _1805;
    wire [31:0] _1807;
    wire [31:0] _111;
    reg [31:0] _1804;
    wire [7:0] _1808;
    wire _1809;
    wire _1810;
    wire [31:0] _1814;
    wire [31:0] _1816;
    wire [31:0] _112;
    reg [31:0] _1813;
    wire [7:0] _1817;
    wire _1818;
    wire _1819;
    wire [31:0] _1823;
    wire [31:0] _1825;
    wire [31:0] _113;
    reg [31:0] _1822;
    wire [7:0] _1826;
    wire _1827;
    wire _1828;
    wire [31:0] _1832;
    wire [31:0] _1834;
    wire [31:0] _114;
    reg [31:0] _1831;
    wire [7:0] _1835;
    wire _1836;
    wire _1837;
    wire [31:0] _1841;
    wire [31:0] _1843;
    wire [31:0] _115;
    reg [31:0] _1840;
    wire [7:0] _1844;
    wire _1845;
    wire _1846;
    wire [31:0] _1850;
    wire [31:0] _1852;
    wire [31:0] _116;
    reg [31:0] _1849;
    wire [7:0] _1853;
    wire _1854;
    wire _1855;
    wire [31:0] _1859;
    wire [31:0] _1861;
    wire [31:0] _117;
    reg [31:0] _1858;
    wire [7:0] _1862;
    wire _1863;
    wire _1864;
    wire [31:0] _1868;
    wire [31:0] _1870;
    wire [31:0] _118;
    reg [31:0] _1867;
    wire [7:0] _1871;
    wire _1872;
    wire _1873;
    wire [31:0] _1877;
    wire [31:0] _1879;
    wire [31:0] _119;
    reg [31:0] _1876;
    wire [7:0] _1880;
    wire _1881;
    wire _1882;
    wire [31:0] _1886;
    wire [31:0] _1888;
    wire [31:0] _120;
    reg [31:0] _1885;
    wire [7:0] _1889;
    wire _1890;
    wire _1891;
    wire [31:0] _1895;
    wire [31:0] _1897;
    wire [31:0] _121;
    reg [31:0] _1894;
    wire [7:0] _1898;
    wire _1899;
    wire _1900;
    wire [31:0] _1904;
    wire [31:0] _1906;
    wire [31:0] _122;
    reg [31:0] _1903;
    wire [7:0] _1907;
    wire _1908;
    wire _1909;
    wire [31:0] _1913;
    wire [31:0] _1915;
    wire [31:0] _123;
    reg [31:0] _1912;
    wire [7:0] _1916;
    wire _1917;
    wire _1918;
    wire [31:0] _1922;
    wire [31:0] _1924;
    wire [31:0] _124;
    reg [31:0] _1921;
    wire [7:0] _1925;
    wire _1926;
    wire _1927;
    wire [31:0] _1931;
    wire [31:0] _1933;
    wire [31:0] _125;
    reg [31:0] _1930;
    wire [7:0] _1934;
    wire _1935;
    wire _1936;
    wire [31:0] _1940;
    wire [31:0] _1942;
    wire [31:0] _126;
    reg [31:0] _1939;
    wire [7:0] _1943;
    wire _1944;
    wire _1945;
    wire [31:0] _1949;
    wire [31:0] _1951;
    wire [31:0] _127;
    reg [31:0] _1948;
    wire [7:0] _1952;
    wire _1953;
    wire _1954;
    wire [31:0] _1958;
    wire [31:0] _1960;
    wire [31:0] _128;
    reg [31:0] _1957;
    wire [7:0] _1961;
    wire _1962;
    wire _1963;
    wire [31:0] _1967;
    wire [31:0] _1969;
    wire [31:0] _129;
    reg [31:0] _1966;
    wire [7:0] _1970;
    wire _1971;
    wire _1972;
    wire [31:0] _1976;
    wire [31:0] _1978;
    wire [31:0] _130;
    reg [31:0] _1975;
    wire [7:0] _1979;
    wire _1980;
    wire _1981;
    wire [31:0] _1985;
    wire [31:0] _1987;
    wire [31:0] _131;
    reg [31:0] _1984;
    wire [7:0] _1988;
    wire _1989;
    wire _1990;
    wire [31:0] _1994;
    wire [31:0] _1996;
    wire [31:0] _132;
    reg [31:0] _1993;
    wire [7:0] _1997;
    wire _1998;
    wire _1999;
    wire [31:0] _2003;
    wire [31:0] _2005;
    wire [31:0] _133;
    reg [31:0] _2002;
    wire [7:0] _2006;
    wire _2007;
    wire _2008;
    wire [31:0] _2012;
    wire [31:0] _2014;
    wire [31:0] _134;
    reg [31:0] _2011;
    wire [7:0] _2015;
    wire _2016;
    wire _2017;
    wire [31:0] _2021;
    wire [31:0] _2023;
    wire [31:0] _135;
    reg [31:0] _2020;
    wire [7:0] _2024;
    wire _2025;
    wire _2026;
    wire [31:0] _2030;
    wire [31:0] _2032;
    wire [31:0] _136;
    reg [31:0] _2029;
    wire [7:0] _2033;
    wire _2034;
    wire _2035;
    wire [31:0] _2039;
    wire [31:0] _2041;
    wire [31:0] _137;
    reg [31:0] _2038;
    wire [7:0] _2042;
    wire _2043;
    wire _2044;
    wire [31:0] _2048;
    wire [31:0] _2050;
    wire [31:0] _138;
    reg [31:0] _2047;
    wire [7:0] _2051;
    wire _2052;
    wire _2053;
    wire [31:0] _2057;
    wire [31:0] _2059;
    wire [31:0] _139;
    reg [31:0] _2056;
    wire [7:0] _2060;
    wire _2061;
    wire _2062;
    wire [31:0] _2066;
    wire [31:0] _2068;
    wire [31:0] _140;
    reg [31:0] _2065;
    wire [7:0] _2069;
    wire _2070;
    wire _2071;
    wire [31:0] _2075;
    wire [31:0] _2077;
    wire [31:0] _141;
    reg [31:0] _2074;
    wire [7:0] _2078;
    wire _2079;
    wire _2080;
    wire [31:0] _2084;
    wire [31:0] _2086;
    wire [31:0] _142;
    reg [31:0] _2083;
    wire [7:0] _2087;
    wire _2088;
    wire _2089;
    wire [31:0] _2093;
    wire [31:0] _2095;
    wire [31:0] _143;
    reg [31:0] _2092;
    wire [7:0] _2096;
    wire _2097;
    wire _2098;
    wire [31:0] _2102;
    wire [31:0] _2104;
    wire [31:0] _144;
    reg [31:0] _2101;
    wire [7:0] _2105;
    wire _2106;
    wire _2107;
    wire [31:0] _2111;
    wire [31:0] _2113;
    wire [31:0] _145;
    reg [31:0] _2110;
    wire [7:0] _2114;
    wire _2115;
    wire _2116;
    wire [31:0] _2120;
    wire [31:0] _2122;
    wire [31:0] _146;
    reg [31:0] _2119;
    wire [7:0] _2123;
    wire _2124;
    wire _2125;
    wire [31:0] _2129;
    wire [31:0] _2131;
    wire [31:0] _147;
    reg [31:0] _2128;
    wire [7:0] _2132;
    wire _2133;
    wire _2134;
    wire [31:0] _2138;
    wire [31:0] _2140;
    wire [31:0] _148;
    reg [31:0] _2137;
    wire [7:0] _2141;
    wire _2142;
    wire _2143;
    wire [31:0] _2147;
    wire [31:0] _2149;
    wire [31:0] _149;
    reg [31:0] _2146;
    wire [7:0] _2150;
    wire _2151;
    wire _2152;
    wire [31:0] _2156;
    wire [31:0] _2158;
    wire [31:0] _150;
    reg [31:0] _2155;
    wire [7:0] _2159;
    wire _2160;
    wire _2161;
    wire [31:0] _2165;
    wire [31:0] _2167;
    wire [31:0] _151;
    reg [31:0] _2164;
    wire [7:0] _2168;
    wire _2169;
    wire _2170;
    wire [31:0] _2174;
    wire [31:0] _2176;
    wire [31:0] _152;
    reg [31:0] _2173;
    wire [7:0] _2177;
    wire _2178;
    wire _2179;
    wire [31:0] _2183;
    wire [31:0] _2185;
    wire [31:0] _153;
    reg [31:0] _2182;
    wire [7:0] _2186;
    wire _2187;
    wire _2188;
    wire [31:0] _2192;
    wire [31:0] _2194;
    wire [31:0] _154;
    reg [31:0] _2191;
    wire [7:0] _2195;
    wire _2196;
    wire _2197;
    wire [31:0] _2201;
    wire [31:0] _2203;
    wire [31:0] _155;
    reg [31:0] _2200;
    wire [7:0] _2204;
    wire _2205;
    wire _2206;
    wire [31:0] _2210;
    wire [31:0] _2212;
    wire [31:0] _156;
    reg [31:0] _2209;
    wire [7:0] _2213;
    wire _2214;
    wire _2215;
    wire [31:0] _2219;
    wire [31:0] _2221;
    wire [31:0] _157;
    reg [31:0] _2218;
    wire [7:0] _2222;
    wire _2223;
    wire _2224;
    wire [31:0] _2228;
    wire [31:0] _2230;
    wire [31:0] _158;
    reg [31:0] _2227;
    wire [7:0] _2231;
    wire _2232;
    wire _2233;
    wire [31:0] _2237;
    wire [31:0] _2239;
    wire [31:0] _159;
    reg [31:0] _2236;
    wire [7:0] _2240;
    wire _2241;
    wire _2242;
    wire [31:0] _2246;
    wire [31:0] _2248;
    wire [31:0] _160;
    reg [31:0] _2245;
    wire [7:0] _2249;
    wire _2250;
    wire _2251;
    wire [31:0] _2255;
    wire [31:0] _2257;
    wire [31:0] _161;
    reg [31:0] _2254;
    wire [7:0] _2258;
    wire _2259;
    wire _2260;
    wire [31:0] _2264;
    wire [31:0] _2266;
    wire [31:0] _162;
    reg [31:0] _2263;
    wire [7:0] _2267;
    wire _2268;
    wire _2269;
    wire [31:0] _2273;
    wire [31:0] _2275;
    wire [31:0] _163;
    reg [31:0] _2272;
    wire [7:0] _2276;
    wire _2277;
    wire _2278;
    wire [31:0] _2282;
    wire [31:0] _2284;
    wire [31:0] _164;
    reg [31:0] _2281;
    wire [7:0] _2285;
    wire _2286;
    wire _2287;
    wire [31:0] _2291;
    wire [31:0] _2293;
    wire [31:0] _165;
    reg [31:0] _2290;
    wire [7:0] _2294;
    wire _2295;
    wire _2296;
    wire [31:0] _2300;
    wire [31:0] _2302;
    wire [31:0] _166;
    reg [31:0] _2299;
    wire [7:0] _2303;
    wire _2304;
    wire _2305;
    wire [31:0] _2309;
    wire [31:0] _2311;
    wire [31:0] _167;
    reg [31:0] _2308;
    wire [7:0] _2312;
    wire _2313;
    wire _2314;
    wire [31:0] _2318;
    wire [31:0] _2320;
    wire [31:0] _168;
    reg [31:0] _2317;
    wire [7:0] _2321;
    wire _2322;
    wire _2323;
    wire [31:0] _2327;
    wire [31:0] _2329;
    wire [31:0] _169;
    reg [31:0] _2326;
    wire [7:0] _2330;
    wire _2331;
    wire _2332;
    wire [31:0] _2336;
    wire [31:0] _2338;
    wire [31:0] _170;
    reg [31:0] _2335;
    wire [7:0] _2339;
    wire _2340;
    wire _2341;
    wire [31:0] _2345;
    wire [31:0] _2347;
    wire [31:0] _171;
    reg [31:0] _2344;
    wire [7:0] _2348;
    wire _2349;
    wire _2350;
    wire [31:0] _2354;
    wire [31:0] _2356;
    wire [31:0] _172;
    reg [31:0] _2353;
    wire [7:0] _2357;
    wire _2358;
    wire _2359;
    wire [31:0] _2363;
    wire [31:0] _2365;
    wire [31:0] _173;
    reg [31:0] _2362;
    wire [7:0] _2366;
    wire _2367;
    wire _2368;
    wire [31:0] _2372;
    wire [31:0] _2374;
    wire [31:0] _174;
    reg [31:0] _2371;
    wire [7:0] _2375;
    wire _2376;
    wire _2377;
    wire [31:0] _2381;
    wire [31:0] _2383;
    wire [31:0] _175;
    reg [31:0] _2380;
    wire [7:0] _2384;
    wire _2385;
    wire _2386;
    wire [31:0] _2390;
    wire [31:0] _2392;
    wire [31:0] _176;
    reg [31:0] _2389;
    wire [7:0] _2393;
    wire _2394;
    wire _2395;
    wire [31:0] _2399;
    wire [31:0] _2401;
    wire [31:0] _177;
    reg [31:0] _2398;
    wire [7:0] _2402;
    wire _2403;
    wire _2404;
    wire [31:0] _2408;
    wire [31:0] _2410;
    wire [31:0] _178;
    reg [31:0] _2407;
    wire [7:0] _2411;
    wire _2412;
    wire _2413;
    wire [31:0] _2417;
    wire [31:0] _2419;
    wire [31:0] _179;
    reg [31:0] _2416;
    wire [7:0] _2420;
    wire _2421;
    wire _2422;
    wire [31:0] _2426;
    wire [31:0] _2428;
    wire [31:0] _180;
    reg [31:0] _2425;
    wire [7:0] _2429;
    wire _2430;
    wire _2431;
    wire [31:0] _2435;
    wire [31:0] _2437;
    wire [31:0] _181;
    reg [31:0] _2434;
    wire [7:0] _2438;
    wire _2439;
    wire _2440;
    wire [31:0] _2444;
    wire [31:0] _2446;
    wire [31:0] _182;
    reg [31:0] _2443;
    wire [7:0] _2447;
    wire _2448;
    wire _2449;
    wire [31:0] _2453;
    wire [31:0] _2455;
    wire [31:0] _183;
    reg [31:0] _2452;
    wire [7:0] _2456;
    wire _2457;
    wire _2458;
    wire [31:0] _2462;
    wire [31:0] _2464;
    wire [31:0] _184;
    reg [31:0] _2461;
    wire [7:0] _2465;
    wire _2466;
    wire _2467;
    wire [31:0] _2471;
    wire [31:0] _2473;
    wire [31:0] _185;
    reg [31:0] _2470;
    wire [7:0] _2474;
    wire _2475;
    wire _2476;
    wire [31:0] _2480;
    wire [31:0] _2482;
    wire [31:0] _186;
    reg [31:0] _2479;
    wire [7:0] _2483;
    wire _2484;
    wire _2485;
    wire [31:0] _2489;
    wire [31:0] _2491;
    wire [31:0] _187;
    reg [31:0] _2488;
    wire [7:0] _2492;
    wire _2493;
    wire _2494;
    wire [31:0] _2498;
    wire [31:0] _2500;
    wire [31:0] _188;
    reg [31:0] _2497;
    wire [7:0] _2501;
    wire _2502;
    wire _2503;
    wire [31:0] _2507;
    wire [31:0] _2509;
    wire [31:0] _189;
    reg [31:0] _2506;
    wire [7:0] _2510;
    wire _2511;
    wire _2512;
    wire [31:0] _2516;
    wire [31:0] _2518;
    wire [31:0] _190;
    reg [31:0] _2515;
    wire [7:0] _2519;
    wire _2520;
    wire _2521;
    wire [31:0] _2525;
    wire [31:0] _2527;
    wire [31:0] _191;
    reg [31:0] _2524;
    wire [7:0] _2528;
    wire _2529;
    wire _2530;
    wire [31:0] _2534;
    wire [31:0] _2536;
    wire [31:0] _192;
    reg [31:0] _2533;
    wire [7:0] _2537;
    wire _2538;
    wire _2539;
    wire [31:0] _2543;
    wire [31:0] _2545;
    wire [31:0] _193;
    reg [31:0] _2542;
    wire [7:0] _2546;
    wire _2547;
    wire _2548;
    wire [31:0] _2552;
    wire [31:0] _2554;
    wire [31:0] _194;
    reg [31:0] _2551;
    wire [7:0] _2555;
    wire _2556;
    wire _2557;
    wire [31:0] _2561;
    wire [31:0] _2563;
    wire [31:0] _195;
    reg [31:0] _2560;
    wire [7:0] _2564;
    wire _2565;
    wire _2566;
    wire [31:0] _2570;
    wire [31:0] _2572;
    wire [31:0] _196;
    reg [31:0] _2569;
    wire [7:0] _2573;
    wire _2574;
    wire _2575;
    wire [31:0] _2579;
    wire [31:0] _2581;
    wire [31:0] _197;
    reg [31:0] _2578;
    wire [7:0] _2582;
    wire _2583;
    wire _2584;
    wire [31:0] _2588;
    wire [31:0] _2590;
    wire [31:0] _198;
    reg [31:0] _2587;
    wire [7:0] _2591;
    wire _2592;
    wire _2593;
    wire [31:0] _2597;
    wire [31:0] _2599;
    wire [31:0] _199;
    reg [31:0] _2596;
    wire [7:0] _2600;
    wire _2601;
    wire _2602;
    wire [31:0] _2606;
    wire [31:0] _2608;
    wire [31:0] _200;
    reg [31:0] _2605;
    wire [7:0] _2609;
    wire _2610;
    wire _2611;
    wire [31:0] _2615;
    wire [31:0] _2617;
    wire [31:0] _201;
    reg [31:0] _2614;
    wire [7:0] _2618;
    wire _2619;
    wire _2620;
    wire [31:0] _2624;
    wire [31:0] _2626;
    wire [31:0] _202;
    reg [31:0] _2623;
    wire [7:0] _2627;
    wire _2628;
    wire _2629;
    wire [31:0] _2633;
    wire [31:0] _2635;
    wire [31:0] _203;
    reg [31:0] _2632;
    wire [7:0] _2636;
    wire _2637;
    wire _2638;
    wire [31:0] _2642;
    wire [31:0] _2644;
    wire [31:0] _204;
    reg [31:0] _2641;
    wire [7:0] _2645;
    wire _2646;
    wire _2647;
    wire [31:0] _2651;
    wire [31:0] _2653;
    wire [31:0] _205;
    reg [31:0] _2650;
    wire [7:0] _2654;
    wire _2655;
    wire _2656;
    wire [31:0] _2660;
    wire [31:0] _2662;
    wire [31:0] _206;
    reg [31:0] _2659;
    wire [7:0] _2663;
    wire _2664;
    wire _2665;
    wire [31:0] _2669;
    wire [31:0] _2671;
    wire [31:0] _207;
    reg [31:0] _2668;
    wire [7:0] _2672;
    wire _2673;
    wire _2674;
    wire [31:0] _2678;
    wire [31:0] _2680;
    wire [31:0] _208;
    reg [31:0] _2677;
    wire [7:0] _2681;
    wire _2682;
    wire _2683;
    wire [31:0] _2687;
    wire [31:0] _2689;
    wire [31:0] _209;
    reg [31:0] _2686;
    wire [7:0] _2690;
    wire _2691;
    wire _2692;
    wire [31:0] _2696;
    wire [31:0] _2698;
    wire [31:0] _210;
    reg [31:0] _2695;
    wire [7:0] _2699;
    wire _2700;
    wire _2701;
    wire [31:0] _2705;
    wire [31:0] _2707;
    wire [31:0] _211;
    reg [31:0] _2704;
    wire [7:0] _2708;
    wire _2709;
    wire _2710;
    wire [31:0] _2714;
    wire [31:0] _2716;
    wire [31:0] _212;
    reg [31:0] _2713;
    wire [7:0] _2717;
    wire _2718;
    wire _2719;
    wire [31:0] _2723;
    wire [31:0] _2725;
    wire [31:0] _213;
    reg [31:0] _2722;
    wire [7:0] _2726;
    wire _2727;
    wire _2728;
    wire [31:0] _2732;
    wire [31:0] _2734;
    wire [31:0] _214;
    reg [31:0] _2731;
    wire [7:0] _2735;
    wire _2736;
    wire _2737;
    wire [31:0] _2741;
    wire [31:0] _2743;
    wire [31:0] _215;
    reg [31:0] _2740;
    wire [7:0] _2744;
    wire _2745;
    wire _2746;
    wire [31:0] _2750;
    wire [31:0] _2752;
    wire [31:0] _216;
    reg [31:0] _2749;
    wire [7:0] _2753;
    wire _2754;
    wire _2755;
    wire [31:0] _2759;
    wire [31:0] _2761;
    wire [31:0] _217;
    reg [31:0] _2758;
    wire [7:0] _2762;
    wire _2763;
    wire _2764;
    wire [31:0] _2768;
    wire [31:0] _2770;
    wire [31:0] _218;
    reg [31:0] _2767;
    wire [7:0] _2771;
    wire _2772;
    wire _2773;
    wire [31:0] _2777;
    wire [31:0] _2779;
    wire [31:0] _219;
    reg [31:0] _2776;
    wire [7:0] _2780;
    wire _2781;
    wire _2782;
    wire [31:0] _2786;
    wire [31:0] _2788;
    wire [31:0] _220;
    reg [31:0] _2785;
    wire [7:0] _2789;
    wire _2790;
    wire _2791;
    wire [31:0] _2795;
    wire [31:0] _2797;
    wire [31:0] _221;
    reg [31:0] _2794;
    wire [7:0] _2798;
    wire _2799;
    wire _2800;
    wire [31:0] _2804;
    wire [31:0] _2806;
    wire [31:0] _222;
    reg [31:0] _2803;
    wire [7:0] _2807;
    wire _2808;
    wire _2809;
    wire [31:0] _2813;
    wire [31:0] _2815;
    wire [31:0] _223;
    reg [31:0] _2812;
    wire [7:0] _2816;
    wire _2817;
    wire _2818;
    wire [31:0] _2822;
    wire [31:0] _2824;
    wire [31:0] _224;
    reg [31:0] _2821;
    wire [7:0] _2825;
    wire _2826;
    wire _2827;
    wire [31:0] _2831;
    wire [31:0] _2833;
    wire [31:0] _225;
    reg [31:0] _2830;
    wire [7:0] _2834;
    wire _2835;
    wire _2836;
    wire [31:0] _2840;
    wire [31:0] _2842;
    wire [31:0] _226;
    reg [31:0] _2839;
    wire [7:0] _2843;
    wire _2844;
    wire _2845;
    wire [31:0] _2849;
    wire [31:0] _2851;
    wire [31:0] _227;
    reg [31:0] _2848;
    wire [7:0] _2852;
    wire _2853;
    wire _2854;
    wire [31:0] _2858;
    wire [31:0] _2860;
    wire [31:0] _228;
    reg [31:0] _2857;
    wire [7:0] _2861;
    wire _2862;
    wire _2863;
    wire [31:0] _2867;
    wire [31:0] _2869;
    wire [31:0] _229;
    reg [31:0] _2866;
    wire [7:0] _2870;
    wire _2871;
    wire _2872;
    wire [31:0] _2876;
    wire [31:0] _2878;
    wire [31:0] _230;
    reg [31:0] _2875;
    wire [7:0] _2879;
    wire _2880;
    wire _2881;
    wire [31:0] _2885;
    wire [31:0] _2887;
    wire [31:0] _231;
    reg [31:0] _2884;
    wire [7:0] _2888;
    wire _2889;
    wire _2890;
    wire [31:0] _2894;
    wire [31:0] _2896;
    wire [31:0] _232;
    reg [31:0] _2893;
    wire [7:0] _2897;
    wire _2898;
    wire _2899;
    wire [31:0] _2903;
    wire [31:0] _2905;
    wire [31:0] _233;
    reg [31:0] _2902;
    wire [7:0] _2906;
    wire _2907;
    wire _2908;
    wire [31:0] _2912;
    wire [31:0] _2914;
    wire [31:0] _234;
    reg [31:0] _2911;
    wire [7:0] _2915;
    wire _2916;
    wire _2917;
    wire [31:0] _2921;
    wire [31:0] _2923;
    wire [31:0] _235;
    reg [31:0] _2920;
    wire [7:0] _2924;
    wire _2925;
    wire _2926;
    wire [31:0] _2930;
    wire [31:0] _2932;
    wire [31:0] _236;
    reg [31:0] _2929;
    wire [7:0] _2933;
    wire _2934;
    wire _2935;
    wire [31:0] _2939;
    wire [31:0] _2941;
    wire [31:0] _237;
    reg [31:0] _2938;
    wire [7:0] _2942;
    wire _2943;
    wire _2944;
    wire [31:0] _2948;
    wire [31:0] _2950;
    wire [31:0] _238;
    reg [31:0] _2947;
    wire [7:0] _2951;
    wire _2952;
    wire _2953;
    wire [31:0] _2957;
    wire [31:0] _2959;
    wire [31:0] _239;
    reg [31:0] _2956;
    wire [7:0] _2960;
    wire _2961;
    wire _2962;
    wire [31:0] _2966;
    wire [31:0] _2968;
    wire [31:0] _240;
    reg [31:0] _2965;
    wire [7:0] _2969;
    wire _2970;
    wire _2971;
    wire [31:0] _2975;
    wire [31:0] _2977;
    wire [31:0] _241;
    reg [31:0] _2974;
    wire [7:0] _2978;
    wire _2979;
    wire _2980;
    wire [31:0] _2984;
    wire [31:0] _2986;
    wire [31:0] _242;
    reg [31:0] _2983;
    wire [7:0] _2987;
    wire _2988;
    wire _2989;
    wire [31:0] _2993;
    wire [31:0] _2995;
    wire [31:0] _243;
    reg [31:0] _2992;
    wire [7:0] _2996;
    wire _2997;
    wire _2998;
    wire [31:0] _3002;
    wire [31:0] _3004;
    wire [31:0] _244;
    reg [31:0] _3001;
    wire [7:0] _3005;
    wire _3006;
    wire _3007;
    wire [31:0] _3011;
    wire [31:0] _3013;
    wire [31:0] _245;
    reg [31:0] _3010;
    wire [7:0] _3014;
    wire _3015;
    wire _3016;
    wire [31:0] _3020;
    wire [31:0] _3022;
    wire [31:0] _246;
    reg [31:0] _3019;
    wire [7:0] _3023;
    wire _3024;
    wire _3025;
    wire [31:0] _3029;
    wire [31:0] _3031;
    wire [31:0] _247;
    reg [31:0] _3028;
    wire [7:0] _3032;
    wire _3033;
    wire _3034;
    wire [31:0] _3038;
    wire [31:0] _3040;
    wire [31:0] _248;
    reg [31:0] _3037;
    wire [7:0] _3041;
    wire _3042;
    wire _3043;
    wire [31:0] _3047;
    wire [31:0] _3049;
    wire [31:0] _249;
    reg [31:0] _3046;
    wire [7:0] _3050;
    wire _3051;
    wire _3052;
    wire [31:0] _3056;
    wire [31:0] _3058;
    wire [31:0] _250;
    reg [31:0] _3055;
    wire [7:0] _3059;
    wire _3060;
    wire _3061;
    wire [31:0] _3065;
    wire [31:0] _3067;
    wire [31:0] _251;
    reg [31:0] _3064;
    wire [7:0] _3068;
    wire _3069;
    wire _3070;
    wire [31:0] _3074;
    wire [31:0] _3076;
    wire [31:0] _252;
    reg [31:0] _3073;
    wire [7:0] _3077;
    wire _3078;
    wire _3079;
    wire [31:0] _3083;
    wire [31:0] _3085;
    wire [31:0] _253;
    reg [31:0] _3082;
    wire [7:0] _3086;
    wire _3087;
    wire _3088;
    wire [31:0] _3092;
    wire [31:0] _3094;
    wire [31:0] _254;
    reg [31:0] _3091;
    wire [7:0] _3095;
    wire _3096;
    wire _3097;
    wire [31:0] _3101;
    wire [31:0] _3103;
    wire [31:0] _255;
    reg [31:0] _3100;
    wire [7:0] _3104;
    wire _3105;
    wire _3106;
    wire [31:0] _3110;
    wire [31:0] _3112;
    wire [31:0] _256;
    reg [31:0] _3109;
    wire [31:0] _258;
    wire [7:0] _3118;
    wire [7:0] _3116;
    wire [7:0] _3114;
    wire [7:0] _3117;
    wire [7:0] _259;
    reg [7:0] _817;
    wire _3119;
    wire _3120;
    wire [31:0] _3124;
    wire [31:0] _3126;
    wire [31:0] _260;
    reg [31:0] _3123;
    reg [31:0] _4705;
    wire [63:0] _4706;
    wire [127:0] _4710;
    wire [63:0] _4711;
    wire [63:0] _4703;
    wire [63:0] _4712;
    wire [63:0] _261;
    reg [63:0] _4701;
    wire [15:0] _4718;
    wire _5251;
    wire [15:0] _5252;
    wire [15:0] _5253;
    wire [15:0] _5254;
    wire [15:0] _4721;
    wire [15:0] _4723;
    wire [15:0] _5255;
    wire [15:0] _263;
    reg [15:0] _4719;
    wire [47:0] _5282;
    wire [63:0] _5283;
    wire _5250;
    wire [15:0] _5260;
    wire [15:0] _5261;
    wire [15:0] _5257;
    wire [15:0] _5259;
    wire [15:0] _5262;
    wire [15:0] _264;
    reg [15:0] _5249;
    wire [63:0] _5279;
    reg [15:0] _5244;
    wire _5241;
    wire _5239;
    wire _5237;
    wire _5235;
    wire _5233;
    wire _5231;
    wire _5229;
    wire _5227;
    wire _5225;
    wire _5223;
    wire _5221;
    wire _5219;
    wire _5217;
    wire _5215;
    wire _5213;
    wire _5211;
    wire _5209;
    wire _5207;
    wire _5205;
    wire _5203;
    wire _5201;
    wire _5199;
    wire _5197;
    wire _5195;
    wire _5193;
    wire _5191;
    wire _5189;
    wire _5187;
    wire _5185;
    wire _5183;
    wire _5181;
    wire _5179;
    wire _5177;
    wire _5175;
    wire _5173;
    wire _5171;
    wire _5169;
    wire _5167;
    wire _5165;
    wire _5163;
    wire _5161;
    wire _5159;
    wire _5157;
    wire _5155;
    wire _5153;
    wire _5151;
    wire _5149;
    wire _5147;
    wire _5145;
    wire _5143;
    wire _5141;
    wire _5139;
    wire _5137;
    wire _5135;
    wire _5133;
    wire _5131;
    wire _5129;
    wire _5127;
    wire _5125;
    wire _5123;
    wire _5121;
    wire _5119;
    wire _5117;
    wire _5115;
    wire _5113;
    wire _5111;
    wire _5109;
    wire _5107;
    wire _5105;
    wire _5103;
    wire _5101;
    wire _5099;
    wire _5097;
    wire _5095;
    wire _5093;
    wire _5091;
    wire _5089;
    wire _5087;
    wire _5085;
    wire _5083;
    wire _5081;
    wire _5079;
    wire _5077;
    wire _5075;
    wire _5073;
    wire _5071;
    wire _5069;
    wire _5067;
    wire _5065;
    wire _5063;
    wire _5061;
    wire _5059;
    wire _5057;
    wire _5055;
    wire _5053;
    wire _5051;
    wire _5049;
    wire _5047;
    wire _5045;
    wire _5043;
    wire _5041;
    wire _5039;
    wire _5037;
    wire _5035;
    wire _5033;
    wire _5031;
    wire _5029;
    wire _5027;
    wire _5025;
    wire _5023;
    wire _5021;
    wire _5019;
    wire _5017;
    wire _5015;
    wire _5013;
    wire _5011;
    wire _5009;
    wire _5007;
    wire _5005;
    wire _5003;
    wire _5001;
    wire _4999;
    wire _4997;
    wire _4995;
    wire _4993;
    wire _4991;
    wire _4989;
    wire _4987;
    wire _4985;
    wire _4983;
    wire _4981;
    wire _4979;
    wire _4977;
    wire _4975;
    wire _4973;
    wire _4971;
    wire _4969;
    wire _4967;
    wire _4965;
    wire _4963;
    wire _4961;
    wire _4959;
    wire _4957;
    wire _4955;
    wire _4953;
    wire _4951;
    wire _4949;
    wire _4947;
    wire _4945;
    wire _4943;
    wire _4941;
    wire _4939;
    wire _4937;
    wire _4935;
    wire _4933;
    wire _4931;
    wire _4929;
    wire _4927;
    wire _4925;
    wire _4923;
    wire _4921;
    wire _4919;
    wire _4917;
    wire _4915;
    wire _4913;
    wire _4911;
    wire _4909;
    wire _4907;
    wire _4905;
    wire _4903;
    wire _4901;
    wire _4899;
    wire _4897;
    wire _4895;
    wire _4893;
    wire _4891;
    wire _4889;
    wire _4887;
    wire _4885;
    wire _4883;
    wire _4881;
    wire _4879;
    wire _4877;
    wire _4875;
    wire _4873;
    wire _4871;
    wire _4869;
    wire _4867;
    wire _4865;
    wire _4863;
    wire _4861;
    wire _4859;
    wire _4857;
    wire _4855;
    wire _4853;
    wire _4851;
    wire _4849;
    wire _4847;
    wire _4845;
    wire _4843;
    wire _4841;
    wire _4839;
    wire _4837;
    wire _4835;
    wire _4833;
    wire _4831;
    wire _4829;
    wire _4827;
    wire _4825;
    wire _4823;
    wire _4821;
    wire _4819;
    wire _4817;
    wire _4815;
    wire _4813;
    wire _4811;
    wire _4809;
    wire _4807;
    wire _4805;
    wire _4803;
    wire _4801;
    wire _4799;
    wire _4797;
    wire _4795;
    wire _4793;
    wire _4791;
    wire _4789;
    wire _4787;
    wire _4785;
    wire _4783;
    wire _4781;
    wire _4779;
    wire _4777;
    wire _4775;
    wire _4773;
    wire _4771;
    wire _4769;
    wire _4767;
    wire _4765;
    wire _4763;
    wire _4761;
    wire _4759;
    wire _4757;
    wire _4755;
    wire _4753;
    wire _4751;
    wire _4749;
    wire _4747;
    wire _4745;
    wire _4743;
    wire _4741;
    wire _4739;
    wire _4737;
    wire _4735;
    wire _4733;
    wire _4731;
    reg _5242;
    wire [15:0] _5245;
    wire _5246;
    wire [15:0] _5267;
    wire [15:0] _5264;
    wire [15:0] _5266;
    wire [15:0] _5268;
    wire [15:0] _265;
    reg [15:0] _4726;
    wire [63:0] _5277;
    wire [127:0] _5280;
    wire [63:0] _5281;
    wire [127:0] _5284;
    wire [63:0] _5285;
    wire [63:0] _5275;
    wire [63:0] _5286;
    wire [63:0] _266;
    reg [63:0] _5273;
    wire _5288;
    wire [2:0] _809;
    wire [2:0] _5287;
    wire _11990;
    wire _11991;
    wire [2:0] _11992;
    wire [15:0] _4696;
    wire [15:0] _4694;
    wire _4697;
    wire [15:0] _11940;
    wire _5306;
    wire _5300;
    wire _5301;
    wire _5307;
    wire [15:0] _5308;
    wire _5298;
    wire _5299;
    wire [15:0] _5310;
    wire [15:0] _5312;
    wire [15:0] _270;
    reg [15:0] _4690;
    wire _5319;
    wire _5316;
    wire _5317;
    wire _5320;
    wire [15:0] _5321;
    wire _5314;
    wire _5315;
    wire [15:0] _5323;
    wire [15:0] _5325;
    wire [15:0] _271;
    reg [15:0] _4687;
    wire _5332;
    wire _5329;
    wire _5330;
    wire _5333;
    wire [15:0] _5334;
    wire _5327;
    wire _5328;
    wire [15:0] _5336;
    wire [15:0] _5338;
    wire [15:0] _272;
    reg [15:0] _4684;
    wire _5345;
    wire _5342;
    wire _5343;
    wire _5346;
    wire [15:0] _5347;
    wire _5340;
    wire _5341;
    wire [15:0] _5349;
    wire [15:0] _5351;
    wire [15:0] _273;
    reg [15:0] _4681;
    wire _5358;
    wire _5355;
    wire _5356;
    wire _5359;
    wire [15:0] _5360;
    wire _5353;
    wire _5354;
    wire [15:0] _5362;
    wire [15:0] _5364;
    wire [15:0] _274;
    reg [15:0] _4678;
    wire _5371;
    wire _5368;
    wire _5369;
    wire _5372;
    wire [15:0] _5373;
    wire _5366;
    wire _5367;
    wire [15:0] _5375;
    wire [15:0] _5377;
    wire [15:0] _275;
    reg [15:0] _4675;
    wire _5384;
    wire _5381;
    wire _5382;
    wire _5385;
    wire [15:0] _5386;
    wire _5379;
    wire _5380;
    wire [15:0] _5388;
    wire [15:0] _5390;
    wire [15:0] _276;
    reg [15:0] _4672;
    wire _5397;
    wire _5394;
    wire _5395;
    wire _5398;
    wire [15:0] _5399;
    wire _5392;
    wire _5393;
    wire [15:0] _5401;
    wire [15:0] _5403;
    wire [15:0] _277;
    reg [15:0] _4669;
    wire _5410;
    wire _5407;
    wire _5408;
    wire _5411;
    wire [15:0] _5412;
    wire _5405;
    wire _5406;
    wire [15:0] _5414;
    wire [15:0] _5416;
    wire [15:0] _278;
    reg [15:0] _4666;
    wire _5423;
    wire _5420;
    wire _5421;
    wire _5424;
    wire [15:0] _5425;
    wire _5418;
    wire _5419;
    wire [15:0] _5427;
    wire [15:0] _5429;
    wire [15:0] _279;
    reg [15:0] _4663;
    wire _5436;
    wire _5433;
    wire _5434;
    wire _5437;
    wire [15:0] _5438;
    wire _5431;
    wire _5432;
    wire [15:0] _5440;
    wire [15:0] _5442;
    wire [15:0] _280;
    reg [15:0] _4660;
    wire _5449;
    wire _5446;
    wire _5447;
    wire _5450;
    wire [15:0] _5451;
    wire _5444;
    wire _5445;
    wire [15:0] _5453;
    wire [15:0] _5455;
    wire [15:0] _281;
    reg [15:0] _4657;
    wire _5462;
    wire _5459;
    wire _5460;
    wire _5463;
    wire [15:0] _5464;
    wire _5457;
    wire _5458;
    wire [15:0] _5466;
    wire [15:0] _5468;
    wire [15:0] _282;
    reg [15:0] _4654;
    wire _5475;
    wire _5472;
    wire _5473;
    wire _5476;
    wire [15:0] _5477;
    wire _5470;
    wire _5471;
    wire [15:0] _5479;
    wire [15:0] _5481;
    wire [15:0] _283;
    reg [15:0] _4651;
    wire _5488;
    wire _5485;
    wire _5486;
    wire _5489;
    wire [15:0] _5490;
    wire _5483;
    wire _5484;
    wire [15:0] _5492;
    wire [15:0] _5494;
    wire [15:0] _284;
    reg [15:0] _4648;
    wire _5501;
    wire _5498;
    wire _5499;
    wire _5502;
    wire [15:0] _5503;
    wire _5496;
    wire _5497;
    wire [15:0] _5505;
    wire [15:0] _5507;
    wire [15:0] _285;
    reg [15:0] _4645;
    wire _5514;
    wire _5511;
    wire _5512;
    wire _5515;
    wire [15:0] _5516;
    wire _5509;
    wire _5510;
    wire [15:0] _5518;
    wire [15:0] _5520;
    wire [15:0] _286;
    reg [15:0] _4642;
    wire _5527;
    wire _5524;
    wire _5525;
    wire _5528;
    wire [15:0] _5529;
    wire _5522;
    wire _5523;
    wire [15:0] _5531;
    wire [15:0] _5533;
    wire [15:0] _287;
    reg [15:0] _4639;
    wire _5540;
    wire _5537;
    wire _5538;
    wire _5541;
    wire [15:0] _5542;
    wire _5535;
    wire _5536;
    wire [15:0] _5544;
    wire [15:0] _5546;
    wire [15:0] _288;
    reg [15:0] _4636;
    wire _5553;
    wire _5550;
    wire _5551;
    wire _5554;
    wire [15:0] _5555;
    wire _5548;
    wire _5549;
    wire [15:0] _5557;
    wire [15:0] _5559;
    wire [15:0] _289;
    reg [15:0] _4633;
    wire _5566;
    wire _5563;
    wire _5564;
    wire _5567;
    wire [15:0] _5568;
    wire _5561;
    wire _5562;
    wire [15:0] _5570;
    wire [15:0] _5572;
    wire [15:0] _290;
    reg [15:0] _4630;
    wire _5579;
    wire _5576;
    wire _5577;
    wire _5580;
    wire [15:0] _5581;
    wire _5574;
    wire _5575;
    wire [15:0] _5583;
    wire [15:0] _5585;
    wire [15:0] _291;
    reg [15:0] _4627;
    wire _5592;
    wire _5589;
    wire _5590;
    wire _5593;
    wire [15:0] _5594;
    wire _5587;
    wire _5588;
    wire [15:0] _5596;
    wire [15:0] _5598;
    wire [15:0] _292;
    reg [15:0] _4624;
    wire _5605;
    wire _5602;
    wire _5603;
    wire _5606;
    wire [15:0] _5607;
    wire _5600;
    wire _5601;
    wire [15:0] _5609;
    wire [15:0] _5611;
    wire [15:0] _293;
    reg [15:0] _4621;
    wire _5618;
    wire _5615;
    wire _5616;
    wire _5619;
    wire [15:0] _5620;
    wire _5613;
    wire _5614;
    wire [15:0] _5622;
    wire [15:0] _5624;
    wire [15:0] _294;
    reg [15:0] _4618;
    wire _5631;
    wire _5628;
    wire _5629;
    wire _5632;
    wire [15:0] _5633;
    wire _5626;
    wire _5627;
    wire [15:0] _5635;
    wire [15:0] _5637;
    wire [15:0] _295;
    reg [15:0] _4615;
    wire _5644;
    wire _5641;
    wire _5642;
    wire _5645;
    wire [15:0] _5646;
    wire _5639;
    wire _5640;
    wire [15:0] _5648;
    wire [15:0] _5650;
    wire [15:0] _296;
    reg [15:0] _4612;
    wire _5657;
    wire _5654;
    wire _5655;
    wire _5658;
    wire [15:0] _5659;
    wire _5652;
    wire _5653;
    wire [15:0] _5661;
    wire [15:0] _5663;
    wire [15:0] _297;
    reg [15:0] _4609;
    wire _5670;
    wire _5667;
    wire _5668;
    wire _5671;
    wire [15:0] _5672;
    wire _5665;
    wire _5666;
    wire [15:0] _5674;
    wire [15:0] _5676;
    wire [15:0] _298;
    reg [15:0] _4606;
    wire _5683;
    wire _5680;
    wire _5681;
    wire _5684;
    wire [15:0] _5685;
    wire _5678;
    wire _5679;
    wire [15:0] _5687;
    wire [15:0] _5689;
    wire [15:0] _299;
    reg [15:0] _4603;
    wire _5696;
    wire _5693;
    wire _5694;
    wire _5697;
    wire [15:0] _5698;
    wire _5691;
    wire _5692;
    wire [15:0] _5700;
    wire [15:0] _5702;
    wire [15:0] _300;
    reg [15:0] _4600;
    wire _5709;
    wire _5706;
    wire _5707;
    wire _5710;
    wire [15:0] _5711;
    wire _5704;
    wire _5705;
    wire [15:0] _5713;
    wire [15:0] _5715;
    wire [15:0] _301;
    reg [15:0] _4597;
    wire _5722;
    wire _5719;
    wire _5720;
    wire _5723;
    wire [15:0] _5724;
    wire _5717;
    wire _5718;
    wire [15:0] _5726;
    wire [15:0] _5728;
    wire [15:0] _302;
    reg [15:0] _4594;
    wire _5735;
    wire _5732;
    wire _5733;
    wire _5736;
    wire [15:0] _5737;
    wire _5730;
    wire _5731;
    wire [15:0] _5739;
    wire [15:0] _5741;
    wire [15:0] _303;
    reg [15:0] _4591;
    wire _5748;
    wire _5745;
    wire _5746;
    wire _5749;
    wire [15:0] _5750;
    wire _5743;
    wire _5744;
    wire [15:0] _5752;
    wire [15:0] _5754;
    wire [15:0] _304;
    reg [15:0] _4588;
    wire _5761;
    wire _5758;
    wire _5759;
    wire _5762;
    wire [15:0] _5763;
    wire _5756;
    wire _5757;
    wire [15:0] _5765;
    wire [15:0] _5767;
    wire [15:0] _305;
    reg [15:0] _4585;
    wire _5774;
    wire _5771;
    wire _5772;
    wire _5775;
    wire [15:0] _5776;
    wire _5769;
    wire _5770;
    wire [15:0] _5778;
    wire [15:0] _5780;
    wire [15:0] _306;
    reg [15:0] _4582;
    wire _5787;
    wire _5784;
    wire _5785;
    wire _5788;
    wire [15:0] _5789;
    wire _5782;
    wire _5783;
    wire [15:0] _5791;
    wire [15:0] _5793;
    wire [15:0] _307;
    reg [15:0] _4579;
    wire _5800;
    wire _5797;
    wire _5798;
    wire _5801;
    wire [15:0] _5802;
    wire _5795;
    wire _5796;
    wire [15:0] _5804;
    wire [15:0] _5806;
    wire [15:0] _308;
    reg [15:0] _4576;
    wire _5813;
    wire _5810;
    wire _5811;
    wire _5814;
    wire [15:0] _5815;
    wire _5808;
    wire _5809;
    wire [15:0] _5817;
    wire [15:0] _5819;
    wire [15:0] _309;
    reg [15:0] _4573;
    wire _5826;
    wire _5823;
    wire _5824;
    wire _5827;
    wire [15:0] _5828;
    wire _5821;
    wire _5822;
    wire [15:0] _5830;
    wire [15:0] _5832;
    wire [15:0] _310;
    reg [15:0] _4570;
    wire _5839;
    wire _5836;
    wire _5837;
    wire _5840;
    wire [15:0] _5841;
    wire _5834;
    wire _5835;
    wire [15:0] _5843;
    wire [15:0] _5845;
    wire [15:0] _311;
    reg [15:0] _4567;
    wire _5852;
    wire _5849;
    wire _5850;
    wire _5853;
    wire [15:0] _5854;
    wire _5847;
    wire _5848;
    wire [15:0] _5856;
    wire [15:0] _5858;
    wire [15:0] _312;
    reg [15:0] _4564;
    wire _5865;
    wire _5862;
    wire _5863;
    wire _5866;
    wire [15:0] _5867;
    wire _5860;
    wire _5861;
    wire [15:0] _5869;
    wire [15:0] _5871;
    wire [15:0] _313;
    reg [15:0] _4561;
    wire _5878;
    wire _5875;
    wire _5876;
    wire _5879;
    wire [15:0] _5880;
    wire _5873;
    wire _5874;
    wire [15:0] _5882;
    wire [15:0] _5884;
    wire [15:0] _314;
    reg [15:0] _4558;
    wire _5891;
    wire _5888;
    wire _5889;
    wire _5892;
    wire [15:0] _5893;
    wire _5886;
    wire _5887;
    wire [15:0] _5895;
    wire [15:0] _5897;
    wire [15:0] _315;
    reg [15:0] _4555;
    wire _5904;
    wire _5901;
    wire _5902;
    wire _5905;
    wire [15:0] _5906;
    wire _5899;
    wire _5900;
    wire [15:0] _5908;
    wire [15:0] _5910;
    wire [15:0] _316;
    reg [15:0] _4552;
    wire _5917;
    wire _5914;
    wire _5915;
    wire _5918;
    wire [15:0] _5919;
    wire _5912;
    wire _5913;
    wire [15:0] _5921;
    wire [15:0] _5923;
    wire [15:0] _317;
    reg [15:0] _4549;
    wire _5930;
    wire _5927;
    wire _5928;
    wire _5931;
    wire [15:0] _5932;
    wire _5925;
    wire _5926;
    wire [15:0] _5934;
    wire [15:0] _5936;
    wire [15:0] _318;
    reg [15:0] _4546;
    wire _5943;
    wire _5940;
    wire _5941;
    wire _5944;
    wire [15:0] _5945;
    wire _5938;
    wire _5939;
    wire [15:0] _5947;
    wire [15:0] _5949;
    wire [15:0] _319;
    reg [15:0] _4543;
    wire _5956;
    wire _5953;
    wire _5954;
    wire _5957;
    wire [15:0] _5958;
    wire _5951;
    wire _5952;
    wire [15:0] _5960;
    wire [15:0] _5962;
    wire [15:0] _320;
    reg [15:0] _4540;
    wire _5969;
    wire _5966;
    wire _5967;
    wire _5970;
    wire [15:0] _5971;
    wire _5964;
    wire _5965;
    wire [15:0] _5973;
    wire [15:0] _5975;
    wire [15:0] _321;
    reg [15:0] _4537;
    wire _5982;
    wire _5979;
    wire _5980;
    wire _5983;
    wire [15:0] _5984;
    wire _5977;
    wire _5978;
    wire [15:0] _5986;
    wire [15:0] _5988;
    wire [15:0] _322;
    reg [15:0] _4534;
    wire _5995;
    wire _5992;
    wire _5993;
    wire _5996;
    wire [15:0] _5997;
    wire _5990;
    wire _5991;
    wire [15:0] _5999;
    wire [15:0] _6001;
    wire [15:0] _323;
    reg [15:0] _4531;
    wire _6008;
    wire _6005;
    wire _6006;
    wire _6009;
    wire [15:0] _6010;
    wire _6003;
    wire _6004;
    wire [15:0] _6012;
    wire [15:0] _6014;
    wire [15:0] _324;
    reg [15:0] _4528;
    wire _6021;
    wire _6018;
    wire _6019;
    wire _6022;
    wire [15:0] _6023;
    wire _6016;
    wire _6017;
    wire [15:0] _6025;
    wire [15:0] _6027;
    wire [15:0] _325;
    reg [15:0] _4525;
    wire _6034;
    wire _6031;
    wire _6032;
    wire _6035;
    wire [15:0] _6036;
    wire _6029;
    wire _6030;
    wire [15:0] _6038;
    wire [15:0] _6040;
    wire [15:0] _326;
    reg [15:0] _4522;
    wire _6047;
    wire _6044;
    wire _6045;
    wire _6048;
    wire [15:0] _6049;
    wire _6042;
    wire _6043;
    wire [15:0] _6051;
    wire [15:0] _6053;
    wire [15:0] _327;
    reg [15:0] _4519;
    wire _6060;
    wire _6057;
    wire _6058;
    wire _6061;
    wire [15:0] _6062;
    wire _6055;
    wire _6056;
    wire [15:0] _6064;
    wire [15:0] _6066;
    wire [15:0] _328;
    reg [15:0] _4516;
    wire _6073;
    wire _6070;
    wire _6071;
    wire _6074;
    wire [15:0] _6075;
    wire _6068;
    wire _6069;
    wire [15:0] _6077;
    wire [15:0] _6079;
    wire [15:0] _329;
    reg [15:0] _4513;
    wire _6086;
    wire _6083;
    wire _6084;
    wire _6087;
    wire [15:0] _6088;
    wire _6081;
    wire _6082;
    wire [15:0] _6090;
    wire [15:0] _6092;
    wire [15:0] _330;
    reg [15:0] _4510;
    wire _6099;
    wire _6096;
    wire _6097;
    wire _6100;
    wire [15:0] _6101;
    wire _6094;
    wire _6095;
    wire [15:0] _6103;
    wire [15:0] _6105;
    wire [15:0] _331;
    reg [15:0] _4507;
    wire _6112;
    wire _6109;
    wire _6110;
    wire _6113;
    wire [15:0] _6114;
    wire _6107;
    wire _6108;
    wire [15:0] _6116;
    wire [15:0] _6118;
    wire [15:0] _332;
    reg [15:0] _4504;
    wire _6125;
    wire _6122;
    wire _6123;
    wire _6126;
    wire [15:0] _6127;
    wire _6120;
    wire _6121;
    wire [15:0] _6129;
    wire [15:0] _6131;
    wire [15:0] _333;
    reg [15:0] _4501;
    wire _6138;
    wire _6135;
    wire _6136;
    wire _6139;
    wire [15:0] _6140;
    wire _6133;
    wire _6134;
    wire [15:0] _6142;
    wire [15:0] _6144;
    wire [15:0] _334;
    reg [15:0] _4498;
    wire _6151;
    wire _6148;
    wire _6149;
    wire _6152;
    wire [15:0] _6153;
    wire _6146;
    wire _6147;
    wire [15:0] _6155;
    wire [15:0] _6157;
    wire [15:0] _335;
    reg [15:0] _4495;
    wire _6164;
    wire _6161;
    wire _6162;
    wire _6165;
    wire [15:0] _6166;
    wire _6159;
    wire _6160;
    wire [15:0] _6168;
    wire [15:0] _6170;
    wire [15:0] _336;
    reg [15:0] _4492;
    wire _6177;
    wire _6174;
    wire _6175;
    wire _6178;
    wire [15:0] _6179;
    wire _6172;
    wire _6173;
    wire [15:0] _6181;
    wire [15:0] _6183;
    wire [15:0] _337;
    reg [15:0] _4489;
    wire _6190;
    wire _6187;
    wire _6188;
    wire _6191;
    wire [15:0] _6192;
    wire _6185;
    wire _6186;
    wire [15:0] _6194;
    wire [15:0] _6196;
    wire [15:0] _338;
    reg [15:0] _4486;
    wire _6203;
    wire _6200;
    wire _6201;
    wire _6204;
    wire [15:0] _6205;
    wire _6198;
    wire _6199;
    wire [15:0] _6207;
    wire [15:0] _6209;
    wire [15:0] _339;
    reg [15:0] _4483;
    wire _6216;
    wire _6213;
    wire _6214;
    wire _6217;
    wire [15:0] _6218;
    wire _6211;
    wire _6212;
    wire [15:0] _6220;
    wire [15:0] _6222;
    wire [15:0] _340;
    reg [15:0] _4480;
    wire _6229;
    wire _6226;
    wire _6227;
    wire _6230;
    wire [15:0] _6231;
    wire _6224;
    wire _6225;
    wire [15:0] _6233;
    wire [15:0] _6235;
    wire [15:0] _341;
    reg [15:0] _4477;
    wire _6242;
    wire _6239;
    wire _6240;
    wire _6243;
    wire [15:0] _6244;
    wire _6237;
    wire _6238;
    wire [15:0] _6246;
    wire [15:0] _6248;
    wire [15:0] _342;
    reg [15:0] _4474;
    wire _6255;
    wire _6252;
    wire _6253;
    wire _6256;
    wire [15:0] _6257;
    wire _6250;
    wire _6251;
    wire [15:0] _6259;
    wire [15:0] _6261;
    wire [15:0] _343;
    reg [15:0] _4471;
    wire _6268;
    wire _6265;
    wire _6266;
    wire _6269;
    wire [15:0] _6270;
    wire _6263;
    wire _6264;
    wire [15:0] _6272;
    wire [15:0] _6274;
    wire [15:0] _344;
    reg [15:0] _4468;
    wire _6281;
    wire _6278;
    wire _6279;
    wire _6282;
    wire [15:0] _6283;
    wire _6276;
    wire _6277;
    wire [15:0] _6285;
    wire [15:0] _6287;
    wire [15:0] _345;
    reg [15:0] _4465;
    wire _6294;
    wire _6291;
    wire _6292;
    wire _6295;
    wire [15:0] _6296;
    wire _6289;
    wire _6290;
    wire [15:0] _6298;
    wire [15:0] _6300;
    wire [15:0] _346;
    reg [15:0] _4462;
    wire _6307;
    wire _6304;
    wire _6305;
    wire _6308;
    wire [15:0] _6309;
    wire _6302;
    wire _6303;
    wire [15:0] _6311;
    wire [15:0] _6313;
    wire [15:0] _347;
    reg [15:0] _4459;
    wire _6320;
    wire _6317;
    wire _6318;
    wire _6321;
    wire [15:0] _6322;
    wire _6315;
    wire _6316;
    wire [15:0] _6324;
    wire [15:0] _6326;
    wire [15:0] _348;
    reg [15:0] _4456;
    wire _6333;
    wire _6330;
    wire _6331;
    wire _6334;
    wire [15:0] _6335;
    wire _6328;
    wire _6329;
    wire [15:0] _6337;
    wire [15:0] _6339;
    wire [15:0] _349;
    reg [15:0] _4453;
    wire _6346;
    wire _6343;
    wire _6344;
    wire _6347;
    wire [15:0] _6348;
    wire _6341;
    wire _6342;
    wire [15:0] _6350;
    wire [15:0] _6352;
    wire [15:0] _350;
    reg [15:0] _4450;
    wire _6359;
    wire _6356;
    wire _6357;
    wire _6360;
    wire [15:0] _6361;
    wire _6354;
    wire _6355;
    wire [15:0] _6363;
    wire [15:0] _6365;
    wire [15:0] _351;
    reg [15:0] _4447;
    wire _6372;
    wire _6369;
    wire _6370;
    wire _6373;
    wire [15:0] _6374;
    wire _6367;
    wire _6368;
    wire [15:0] _6376;
    wire [15:0] _6378;
    wire [15:0] _352;
    reg [15:0] _4444;
    wire _6385;
    wire _6382;
    wire _6383;
    wire _6386;
    wire [15:0] _6387;
    wire _6380;
    wire _6381;
    wire [15:0] _6389;
    wire [15:0] _6391;
    wire [15:0] _353;
    reg [15:0] _4441;
    wire _6398;
    wire _6395;
    wire _6396;
    wire _6399;
    wire [15:0] _6400;
    wire _6393;
    wire _6394;
    wire [15:0] _6402;
    wire [15:0] _6404;
    wire [15:0] _354;
    reg [15:0] _4438;
    wire _6411;
    wire _6408;
    wire _6409;
    wire _6412;
    wire [15:0] _6413;
    wire _6406;
    wire _6407;
    wire [15:0] _6415;
    wire [15:0] _6417;
    wire [15:0] _355;
    reg [15:0] _4435;
    wire _6424;
    wire _6421;
    wire _6422;
    wire _6425;
    wire [15:0] _6426;
    wire _6419;
    wire _6420;
    wire [15:0] _6428;
    wire [15:0] _6430;
    wire [15:0] _356;
    reg [15:0] _4432;
    wire _6437;
    wire _6434;
    wire _6435;
    wire _6438;
    wire [15:0] _6439;
    wire _6432;
    wire _6433;
    wire [15:0] _6441;
    wire [15:0] _6443;
    wire [15:0] _357;
    reg [15:0] _4429;
    wire _6450;
    wire _6447;
    wire _6448;
    wire _6451;
    wire [15:0] _6452;
    wire _6445;
    wire _6446;
    wire [15:0] _6454;
    wire [15:0] _6456;
    wire [15:0] _358;
    reg [15:0] _4426;
    wire _6463;
    wire _6460;
    wire _6461;
    wire _6464;
    wire [15:0] _6465;
    wire _6458;
    wire _6459;
    wire [15:0] _6467;
    wire [15:0] _6469;
    wire [15:0] _359;
    reg [15:0] _4423;
    wire _6476;
    wire _6473;
    wire _6474;
    wire _6477;
    wire [15:0] _6478;
    wire _6471;
    wire _6472;
    wire [15:0] _6480;
    wire [15:0] _6482;
    wire [15:0] _360;
    reg [15:0] _4420;
    wire _6489;
    wire _6486;
    wire _6487;
    wire _6490;
    wire [15:0] _6491;
    wire _6484;
    wire _6485;
    wire [15:0] _6493;
    wire [15:0] _6495;
    wire [15:0] _361;
    reg [15:0] _4417;
    wire _6502;
    wire _6499;
    wire _6500;
    wire _6503;
    wire [15:0] _6504;
    wire _6497;
    wire _6498;
    wire [15:0] _6506;
    wire [15:0] _6508;
    wire [15:0] _362;
    reg [15:0] _4414;
    wire _6515;
    wire _6512;
    wire _6513;
    wire _6516;
    wire [15:0] _6517;
    wire _6510;
    wire _6511;
    wire [15:0] _6519;
    wire [15:0] _6521;
    wire [15:0] _363;
    reg [15:0] _4411;
    wire _6528;
    wire _6525;
    wire _6526;
    wire _6529;
    wire [15:0] _6530;
    wire _6523;
    wire _6524;
    wire [15:0] _6532;
    wire [15:0] _6534;
    wire [15:0] _364;
    reg [15:0] _4408;
    wire _6541;
    wire _6538;
    wire _6539;
    wire _6542;
    wire [15:0] _6543;
    wire _6536;
    wire _6537;
    wire [15:0] _6545;
    wire [15:0] _6547;
    wire [15:0] _365;
    reg [15:0] _4405;
    wire _6554;
    wire _6551;
    wire _6552;
    wire _6555;
    wire [15:0] _6556;
    wire _6549;
    wire _6550;
    wire [15:0] _6558;
    wire [15:0] _6560;
    wire [15:0] _366;
    reg [15:0] _4402;
    wire _6567;
    wire _6564;
    wire _6565;
    wire _6568;
    wire [15:0] _6569;
    wire _6562;
    wire _6563;
    wire [15:0] _6571;
    wire [15:0] _6573;
    wire [15:0] _367;
    reg [15:0] _4399;
    wire _6580;
    wire _6577;
    wire _6578;
    wire _6581;
    wire [15:0] _6582;
    wire _6575;
    wire _6576;
    wire [15:0] _6584;
    wire [15:0] _6586;
    wire [15:0] _368;
    reg [15:0] _4396;
    wire _6593;
    wire _6590;
    wire _6591;
    wire _6594;
    wire [15:0] _6595;
    wire _6588;
    wire _6589;
    wire [15:0] _6597;
    wire [15:0] _6599;
    wire [15:0] _369;
    reg [15:0] _4393;
    wire _6606;
    wire _6603;
    wire _6604;
    wire _6607;
    wire [15:0] _6608;
    wire _6601;
    wire _6602;
    wire [15:0] _6610;
    wire [15:0] _6612;
    wire [15:0] _370;
    reg [15:0] _4390;
    wire _6619;
    wire _6616;
    wire _6617;
    wire _6620;
    wire [15:0] _6621;
    wire _6614;
    wire _6615;
    wire [15:0] _6623;
    wire [15:0] _6625;
    wire [15:0] _371;
    reg [15:0] _4387;
    wire _6632;
    wire _6629;
    wire _6630;
    wire _6633;
    wire [15:0] _6634;
    wire _6627;
    wire _6628;
    wire [15:0] _6636;
    wire [15:0] _6638;
    wire [15:0] _372;
    reg [15:0] _4384;
    wire _6645;
    wire _6642;
    wire _6643;
    wire _6646;
    wire [15:0] _6647;
    wire _6640;
    wire _6641;
    wire [15:0] _6649;
    wire [15:0] _6651;
    wire [15:0] _373;
    reg [15:0] _4381;
    wire _6658;
    wire _6655;
    wire _6656;
    wire _6659;
    wire [15:0] _6660;
    wire _6653;
    wire _6654;
    wire [15:0] _6662;
    wire [15:0] _6664;
    wire [15:0] _374;
    reg [15:0] _4378;
    wire _6671;
    wire _6668;
    wire _6669;
    wire _6672;
    wire [15:0] _6673;
    wire _6666;
    wire _6667;
    wire [15:0] _6675;
    wire [15:0] _6677;
    wire [15:0] _375;
    reg [15:0] _4375;
    wire _6684;
    wire _6681;
    wire _6682;
    wire _6685;
    wire [15:0] _6686;
    wire _6679;
    wire _6680;
    wire [15:0] _6688;
    wire [15:0] _6690;
    wire [15:0] _376;
    reg [15:0] _4372;
    wire _6697;
    wire _6694;
    wire _6695;
    wire _6698;
    wire [15:0] _6699;
    wire _6692;
    wire _6693;
    wire [15:0] _6701;
    wire [15:0] _6703;
    wire [15:0] _377;
    reg [15:0] _4369;
    wire _6710;
    wire _6707;
    wire _6708;
    wire _6711;
    wire [15:0] _6712;
    wire _6705;
    wire _6706;
    wire [15:0] _6714;
    wire [15:0] _6716;
    wire [15:0] _378;
    reg [15:0] _4366;
    wire _6723;
    wire _6720;
    wire _6721;
    wire _6724;
    wire [15:0] _6725;
    wire _6718;
    wire _6719;
    wire [15:0] _6727;
    wire [15:0] _6729;
    wire [15:0] _379;
    reg [15:0] _4363;
    wire _6736;
    wire _6733;
    wire _6734;
    wire _6737;
    wire [15:0] _6738;
    wire _6731;
    wire _6732;
    wire [15:0] _6740;
    wire [15:0] _6742;
    wire [15:0] _380;
    reg [15:0] _4360;
    wire _6749;
    wire _6746;
    wire _6747;
    wire _6750;
    wire [15:0] _6751;
    wire _6744;
    wire _6745;
    wire [15:0] _6753;
    wire [15:0] _6755;
    wire [15:0] _381;
    reg [15:0] _4357;
    wire _6762;
    wire _6759;
    wire _6760;
    wire _6763;
    wire [15:0] _6764;
    wire _6757;
    wire _6758;
    wire [15:0] _6766;
    wire [15:0] _6768;
    wire [15:0] _382;
    reg [15:0] _4354;
    wire _6775;
    wire _6772;
    wire _6773;
    wire _6776;
    wire [15:0] _6777;
    wire _6770;
    wire _6771;
    wire [15:0] _6779;
    wire [15:0] _6781;
    wire [15:0] _383;
    reg [15:0] _4351;
    wire _6788;
    wire _6785;
    wire _6786;
    wire _6789;
    wire [15:0] _6790;
    wire _6783;
    wire _6784;
    wire [15:0] _6792;
    wire [15:0] _6794;
    wire [15:0] _384;
    reg [15:0] _4348;
    wire _6801;
    wire _6798;
    wire _6799;
    wire _6802;
    wire [15:0] _6803;
    wire _6796;
    wire _6797;
    wire [15:0] _6805;
    wire [15:0] _6807;
    wire [15:0] _385;
    reg [15:0] _4345;
    wire _6814;
    wire _6811;
    wire _6812;
    wire _6815;
    wire [15:0] _6816;
    wire _6809;
    wire _6810;
    wire [15:0] _6818;
    wire [15:0] _6820;
    wire [15:0] _386;
    reg [15:0] _4342;
    wire _6827;
    wire _6824;
    wire _6825;
    wire _6828;
    wire [15:0] _6829;
    wire _6822;
    wire _6823;
    wire [15:0] _6831;
    wire [15:0] _6833;
    wire [15:0] _387;
    reg [15:0] _4339;
    wire _6840;
    wire _6837;
    wire _6838;
    wire _6841;
    wire [15:0] _6842;
    wire _6835;
    wire _6836;
    wire [15:0] _6844;
    wire [15:0] _6846;
    wire [15:0] _388;
    reg [15:0] _4336;
    wire _6853;
    wire _6850;
    wire _6851;
    wire _6854;
    wire [15:0] _6855;
    wire _6848;
    wire _6849;
    wire [15:0] _6857;
    wire [15:0] _6859;
    wire [15:0] _389;
    reg [15:0] _4333;
    wire _6866;
    wire _6863;
    wire _6864;
    wire _6867;
    wire [15:0] _6868;
    wire _6861;
    wire _6862;
    wire [15:0] _6870;
    wire [15:0] _6872;
    wire [15:0] _390;
    reg [15:0] _4330;
    wire _6879;
    wire _6876;
    wire _6877;
    wire _6880;
    wire [15:0] _6881;
    wire _6874;
    wire _6875;
    wire [15:0] _6883;
    wire [15:0] _6885;
    wire [15:0] _391;
    reg [15:0] _4327;
    wire _6892;
    wire _6889;
    wire _6890;
    wire _6893;
    wire [15:0] _6894;
    wire _6887;
    wire _6888;
    wire [15:0] _6896;
    wire [15:0] _6898;
    wire [15:0] _392;
    reg [15:0] _4324;
    wire _6905;
    wire _6902;
    wire _6903;
    wire _6906;
    wire [15:0] _6907;
    wire _6900;
    wire _6901;
    wire [15:0] _6909;
    wire [15:0] _6911;
    wire [15:0] _393;
    reg [15:0] _4321;
    wire _6918;
    wire _6915;
    wire _6916;
    wire _6919;
    wire [15:0] _6920;
    wire _6913;
    wire _6914;
    wire [15:0] _6922;
    wire [15:0] _6924;
    wire [15:0] _394;
    reg [15:0] _4318;
    wire _6931;
    wire _6928;
    wire _6929;
    wire _6932;
    wire [15:0] _6933;
    wire _6926;
    wire _6927;
    wire [15:0] _6935;
    wire [15:0] _6937;
    wire [15:0] _395;
    reg [15:0] _4315;
    wire _6944;
    wire _6941;
    wire _6942;
    wire _6945;
    wire [15:0] _6946;
    wire _6939;
    wire _6940;
    wire [15:0] _6948;
    wire [15:0] _6950;
    wire [15:0] _396;
    reg [15:0] _4312;
    wire _6957;
    wire _6954;
    wire _6955;
    wire _6958;
    wire [15:0] _6959;
    wire _6952;
    wire _6953;
    wire [15:0] _6961;
    wire [15:0] _6963;
    wire [15:0] _397;
    reg [15:0] _4309;
    wire _6970;
    wire _6967;
    wire _6968;
    wire _6971;
    wire [15:0] _6972;
    wire _6965;
    wire _6966;
    wire [15:0] _6974;
    wire [15:0] _6976;
    wire [15:0] _398;
    reg [15:0] _4306;
    wire _6983;
    wire _6980;
    wire _6981;
    wire _6984;
    wire [15:0] _6985;
    wire _6978;
    wire _6979;
    wire [15:0] _6987;
    wire [15:0] _6989;
    wire [15:0] _399;
    reg [15:0] _4303;
    wire _6996;
    wire _6993;
    wire _6994;
    wire _6997;
    wire [15:0] _6998;
    wire _6991;
    wire _6992;
    wire [15:0] _7000;
    wire [15:0] _7002;
    wire [15:0] _400;
    reg [15:0] _4300;
    wire _7009;
    wire _7006;
    wire _7007;
    wire _7010;
    wire [15:0] _7011;
    wire _7004;
    wire _7005;
    wire [15:0] _7013;
    wire [15:0] _7015;
    wire [15:0] _401;
    reg [15:0] _4297;
    wire _7022;
    wire _7019;
    wire _7020;
    wire _7023;
    wire [15:0] _7024;
    wire _7017;
    wire _7018;
    wire [15:0] _7026;
    wire [15:0] _7028;
    wire [15:0] _402;
    reg [15:0] _4294;
    wire _7035;
    wire _7032;
    wire _7033;
    wire _7036;
    wire [15:0] _7037;
    wire _7030;
    wire _7031;
    wire [15:0] _7039;
    wire [15:0] _7041;
    wire [15:0] _403;
    reg [15:0] _4291;
    wire _7048;
    wire _7045;
    wire _7046;
    wire _7049;
    wire [15:0] _7050;
    wire _7043;
    wire _7044;
    wire [15:0] _7052;
    wire [15:0] _7054;
    wire [15:0] _404;
    reg [15:0] _4288;
    wire _7061;
    wire _7058;
    wire _7059;
    wire _7062;
    wire [15:0] _7063;
    wire _7056;
    wire _7057;
    wire [15:0] _7065;
    wire [15:0] _7067;
    wire [15:0] _405;
    reg [15:0] _4285;
    wire _7074;
    wire _7071;
    wire _7072;
    wire _7075;
    wire [15:0] _7076;
    wire _7069;
    wire _7070;
    wire [15:0] _7078;
    wire [15:0] _7080;
    wire [15:0] _406;
    reg [15:0] _4282;
    wire _7087;
    wire _7084;
    wire _7085;
    wire _7088;
    wire [15:0] _7089;
    wire _7082;
    wire _7083;
    wire [15:0] _7091;
    wire [15:0] _7093;
    wire [15:0] _407;
    reg [15:0] _4279;
    wire _7100;
    wire _7097;
    wire _7098;
    wire _7101;
    wire [15:0] _7102;
    wire _7095;
    wire _7096;
    wire [15:0] _7104;
    wire [15:0] _7106;
    wire [15:0] _408;
    reg [15:0] _4276;
    wire _7113;
    wire _7110;
    wire _7111;
    wire _7114;
    wire [15:0] _7115;
    wire _7108;
    wire _7109;
    wire [15:0] _7117;
    wire [15:0] _7119;
    wire [15:0] _409;
    reg [15:0] _4273;
    wire _7126;
    wire _7123;
    wire _7124;
    wire _7127;
    wire [15:0] _7128;
    wire _7121;
    wire _7122;
    wire [15:0] _7130;
    wire [15:0] _7132;
    wire [15:0] _410;
    reg [15:0] _4270;
    wire _7139;
    wire _7136;
    wire _7137;
    wire _7140;
    wire [15:0] _7141;
    wire _7134;
    wire _7135;
    wire [15:0] _7143;
    wire [15:0] _7145;
    wire [15:0] _411;
    reg [15:0] _4267;
    wire _7152;
    wire _7149;
    wire _7150;
    wire _7153;
    wire [15:0] _7154;
    wire _7147;
    wire _7148;
    wire [15:0] _7156;
    wire [15:0] _7158;
    wire [15:0] _412;
    reg [15:0] _4264;
    wire _7165;
    wire _7162;
    wire _7163;
    wire _7166;
    wire [15:0] _7167;
    wire _7160;
    wire _7161;
    wire [15:0] _7169;
    wire [15:0] _7171;
    wire [15:0] _413;
    reg [15:0] _4261;
    wire _7178;
    wire _7175;
    wire _7176;
    wire _7179;
    wire [15:0] _7180;
    wire _7173;
    wire _7174;
    wire [15:0] _7182;
    wire [15:0] _7184;
    wire [15:0] _414;
    reg [15:0] _4258;
    wire _7191;
    wire _7188;
    wire _7189;
    wire _7192;
    wire [15:0] _7193;
    wire _7186;
    wire _7187;
    wire [15:0] _7195;
    wire [15:0] _7197;
    wire [15:0] _415;
    reg [15:0] _4255;
    wire _7204;
    wire _7201;
    wire _7202;
    wire _7205;
    wire [15:0] _7206;
    wire _7199;
    wire _7200;
    wire [15:0] _7208;
    wire [15:0] _7210;
    wire [15:0] _416;
    reg [15:0] _4252;
    wire _7217;
    wire _7214;
    wire _7215;
    wire _7218;
    wire [15:0] _7219;
    wire _7212;
    wire _7213;
    wire [15:0] _7221;
    wire [15:0] _7223;
    wire [15:0] _417;
    reg [15:0] _4249;
    wire _7230;
    wire _7227;
    wire _7228;
    wire _7231;
    wire [15:0] _7232;
    wire _7225;
    wire _7226;
    wire [15:0] _7234;
    wire [15:0] _7236;
    wire [15:0] _418;
    reg [15:0] _4246;
    wire _7243;
    wire _7240;
    wire _7241;
    wire _7244;
    wire [15:0] _7245;
    wire _7238;
    wire _7239;
    wire [15:0] _7247;
    wire [15:0] _7249;
    wire [15:0] _419;
    reg [15:0] _4243;
    wire _7256;
    wire _7253;
    wire _7254;
    wire _7257;
    wire [15:0] _7258;
    wire _7251;
    wire _7252;
    wire [15:0] _7260;
    wire [15:0] _7262;
    wire [15:0] _420;
    reg [15:0] _4240;
    wire _7269;
    wire _7266;
    wire _7267;
    wire _7270;
    wire [15:0] _7271;
    wire _7264;
    wire _7265;
    wire [15:0] _7273;
    wire [15:0] _7275;
    wire [15:0] _421;
    reg [15:0] _4237;
    wire _7282;
    wire _7279;
    wire _7280;
    wire _7283;
    wire [15:0] _7284;
    wire _7277;
    wire _7278;
    wire [15:0] _7286;
    wire [15:0] _7288;
    wire [15:0] _422;
    reg [15:0] _4234;
    wire _7295;
    wire _7292;
    wire _7293;
    wire _7296;
    wire [15:0] _7297;
    wire _7290;
    wire _7291;
    wire [15:0] _7299;
    wire [15:0] _7301;
    wire [15:0] _423;
    reg [15:0] _4231;
    wire _7308;
    wire _7305;
    wire _7306;
    wire _7309;
    wire [15:0] _7310;
    wire _7303;
    wire _7304;
    wire [15:0] _7312;
    wire [15:0] _7314;
    wire [15:0] _424;
    reg [15:0] _4228;
    wire _7321;
    wire _7318;
    wire _7319;
    wire _7322;
    wire [15:0] _7323;
    wire _7316;
    wire _7317;
    wire [15:0] _7325;
    wire [15:0] _7327;
    wire [15:0] _425;
    reg [15:0] _4225;
    wire _7334;
    wire _7331;
    wire _7332;
    wire _7335;
    wire [15:0] _7336;
    wire _7329;
    wire _7330;
    wire [15:0] _7338;
    wire [15:0] _7340;
    wire [15:0] _426;
    reg [15:0] _4222;
    wire _7347;
    wire _7344;
    wire _7345;
    wire _7348;
    wire [15:0] _7349;
    wire _7342;
    wire _7343;
    wire [15:0] _7351;
    wire [15:0] _7353;
    wire [15:0] _427;
    reg [15:0] _4219;
    wire _7360;
    wire _7357;
    wire _7358;
    wire _7361;
    wire [15:0] _7362;
    wire _7355;
    wire _7356;
    wire [15:0] _7364;
    wire [15:0] _7366;
    wire [15:0] _428;
    reg [15:0] _4216;
    wire _7373;
    wire _7370;
    wire _7371;
    wire _7374;
    wire [15:0] _7375;
    wire _7368;
    wire _7369;
    wire [15:0] _7377;
    wire [15:0] _7379;
    wire [15:0] _429;
    reg [15:0] _4213;
    wire _7386;
    wire _7383;
    wire _7384;
    wire _7387;
    wire [15:0] _7388;
    wire _7381;
    wire _7382;
    wire [15:0] _7390;
    wire [15:0] _7392;
    wire [15:0] _430;
    reg [15:0] _4210;
    wire _7399;
    wire _7396;
    wire _7397;
    wire _7400;
    wire [15:0] _7401;
    wire _7394;
    wire _7395;
    wire [15:0] _7403;
    wire [15:0] _7405;
    wire [15:0] _431;
    reg [15:0] _4207;
    wire _7412;
    wire _7409;
    wire _7410;
    wire _7413;
    wire [15:0] _7414;
    wire _7407;
    wire _7408;
    wire [15:0] _7416;
    wire [15:0] _7418;
    wire [15:0] _432;
    reg [15:0] _4204;
    wire _7425;
    wire _7422;
    wire _7423;
    wire _7426;
    wire [15:0] _7427;
    wire _7420;
    wire _7421;
    wire [15:0] _7429;
    wire [15:0] _7431;
    wire [15:0] _433;
    reg [15:0] _4201;
    wire _7438;
    wire _7435;
    wire _7436;
    wire _7439;
    wire [15:0] _7440;
    wire _7433;
    wire _7434;
    wire [15:0] _7442;
    wire [15:0] _7444;
    wire [15:0] _434;
    reg [15:0] _4198;
    wire _7451;
    wire _7448;
    wire _7449;
    wire _7452;
    wire [15:0] _7453;
    wire _7446;
    wire _7447;
    wire [15:0] _7455;
    wire [15:0] _7457;
    wire [15:0] _435;
    reg [15:0] _4195;
    wire _7464;
    wire _7461;
    wire _7462;
    wire _7465;
    wire [15:0] _7466;
    wire _7459;
    wire _7460;
    wire [15:0] _7468;
    wire [15:0] _7470;
    wire [15:0] _436;
    reg [15:0] _4192;
    wire _7477;
    wire _7474;
    wire _7475;
    wire _7478;
    wire [15:0] _7479;
    wire _7472;
    wire _7473;
    wire [15:0] _7481;
    wire [15:0] _7483;
    wire [15:0] _437;
    reg [15:0] _4189;
    wire _7490;
    wire _7487;
    wire _7488;
    wire _7491;
    wire [15:0] _7492;
    wire _7485;
    wire _7486;
    wire [15:0] _7494;
    wire [15:0] _7496;
    wire [15:0] _438;
    reg [15:0] _4186;
    wire _7503;
    wire _7500;
    wire _7501;
    wire _7504;
    wire [15:0] _7505;
    wire _7498;
    wire _7499;
    wire [15:0] _7507;
    wire [15:0] _7509;
    wire [15:0] _439;
    reg [15:0] _4183;
    wire _7516;
    wire _7513;
    wire _7514;
    wire _7517;
    wire [15:0] _7518;
    wire _7511;
    wire _7512;
    wire [15:0] _7520;
    wire [15:0] _7522;
    wire [15:0] _440;
    reg [15:0] _4180;
    wire _7529;
    wire _7526;
    wire _7527;
    wire _7530;
    wire [15:0] _7531;
    wire _7524;
    wire _7525;
    wire [15:0] _7533;
    wire [15:0] _7535;
    wire [15:0] _441;
    reg [15:0] _4177;
    wire _7542;
    wire _7539;
    wire _7540;
    wire _7543;
    wire [15:0] _7544;
    wire _7537;
    wire _7538;
    wire [15:0] _7546;
    wire [15:0] _7548;
    wire [15:0] _442;
    reg [15:0] _4174;
    wire _7555;
    wire _7552;
    wire _7553;
    wire _7556;
    wire [15:0] _7557;
    wire _7550;
    wire _7551;
    wire [15:0] _7559;
    wire [15:0] _7561;
    wire [15:0] _443;
    reg [15:0] _4171;
    wire _7568;
    wire _7565;
    wire _7566;
    wire _7569;
    wire [15:0] _7570;
    wire _7563;
    wire _7564;
    wire [15:0] _7572;
    wire [15:0] _7574;
    wire [15:0] _444;
    reg [15:0] _4168;
    wire _7581;
    wire _7578;
    wire _7579;
    wire _7582;
    wire [15:0] _7583;
    wire _7576;
    wire _7577;
    wire [15:0] _7585;
    wire [15:0] _7587;
    wire [15:0] _445;
    reg [15:0] _4165;
    wire _7594;
    wire _7591;
    wire _7592;
    wire _7595;
    wire [15:0] _7596;
    wire _7589;
    wire _7590;
    wire [15:0] _7598;
    wire [15:0] _7600;
    wire [15:0] _446;
    reg [15:0] _4162;
    wire _7607;
    wire _7604;
    wire _7605;
    wire _7608;
    wire [15:0] _7609;
    wire _7602;
    wire _7603;
    wire [15:0] _7611;
    wire [15:0] _7613;
    wire [15:0] _447;
    reg [15:0] _4159;
    wire _7620;
    wire _7617;
    wire _7618;
    wire _7621;
    wire [15:0] _7622;
    wire _7615;
    wire _7616;
    wire [15:0] _7624;
    wire [15:0] _7626;
    wire [15:0] _448;
    reg [15:0] _4156;
    wire _7633;
    wire _7630;
    wire _7631;
    wire _7634;
    wire [15:0] _7635;
    wire _7628;
    wire _7629;
    wire [15:0] _7637;
    wire [15:0] _7639;
    wire [15:0] _449;
    reg [15:0] _4153;
    wire _7646;
    wire _7643;
    wire _7644;
    wire _7647;
    wire [15:0] _7648;
    wire _7641;
    wire _7642;
    wire [15:0] _7650;
    wire [15:0] _7652;
    wire [15:0] _450;
    reg [15:0] _4150;
    wire _7659;
    wire _7656;
    wire _7657;
    wire _7660;
    wire [15:0] _7661;
    wire _7654;
    wire _7655;
    wire [15:0] _7663;
    wire [15:0] _7665;
    wire [15:0] _451;
    reg [15:0] _4147;
    wire _7672;
    wire _7669;
    wire _7670;
    wire _7673;
    wire [15:0] _7674;
    wire _7667;
    wire _7668;
    wire [15:0] _7676;
    wire [15:0] _7678;
    wire [15:0] _452;
    reg [15:0] _4144;
    wire _7685;
    wire _7682;
    wire _7683;
    wire _7686;
    wire [15:0] _7687;
    wire _7680;
    wire _7681;
    wire [15:0] _7689;
    wire [15:0] _7691;
    wire [15:0] _453;
    reg [15:0] _4141;
    wire _7698;
    wire _7695;
    wire _7696;
    wire _7699;
    wire [15:0] _7700;
    wire _7693;
    wire _7694;
    wire [15:0] _7702;
    wire [15:0] _7704;
    wire [15:0] _454;
    reg [15:0] _4138;
    wire _7711;
    wire _7708;
    wire _7709;
    wire _7712;
    wire [15:0] _7713;
    wire _7706;
    wire _7707;
    wire [15:0] _7715;
    wire [15:0] _7717;
    wire [15:0] _455;
    reg [15:0] _4135;
    wire _7724;
    wire _7721;
    wire _7722;
    wire _7725;
    wire [15:0] _7726;
    wire _7719;
    wire _7720;
    wire [15:0] _7728;
    wire [15:0] _7730;
    wire [15:0] _456;
    reg [15:0] _4132;
    wire _7737;
    wire _7734;
    wire _7735;
    wire _7738;
    wire [15:0] _7739;
    wire _7732;
    wire _7733;
    wire [15:0] _7741;
    wire [15:0] _7743;
    wire [15:0] _457;
    reg [15:0] _4129;
    wire _7750;
    wire _7747;
    wire _7748;
    wire _7751;
    wire [15:0] _7752;
    wire _7745;
    wire _7746;
    wire [15:0] _7754;
    wire [15:0] _7756;
    wire [15:0] _458;
    reg [15:0] _4126;
    wire _7763;
    wire _7760;
    wire _7761;
    wire _7764;
    wire [15:0] _7765;
    wire _7758;
    wire _7759;
    wire [15:0] _7767;
    wire [15:0] _7769;
    wire [15:0] _459;
    reg [15:0] _4123;
    wire _7776;
    wire _7773;
    wire _7774;
    wire _7777;
    wire [15:0] _7778;
    wire _7771;
    wire _7772;
    wire [15:0] _7780;
    wire [15:0] _7782;
    wire [15:0] _460;
    reg [15:0] _4120;
    wire _7789;
    wire _7786;
    wire _7787;
    wire _7790;
    wire [15:0] _7791;
    wire _7784;
    wire _7785;
    wire [15:0] _7793;
    wire [15:0] _7795;
    wire [15:0] _461;
    reg [15:0] _4117;
    wire _7802;
    wire _7799;
    wire _7800;
    wire _7803;
    wire [15:0] _7804;
    wire _7797;
    wire _7798;
    wire [15:0] _7806;
    wire [15:0] _7808;
    wire [15:0] _462;
    reg [15:0] _4114;
    wire _7815;
    wire _7812;
    wire _7813;
    wire _7816;
    wire [15:0] _7817;
    wire _7810;
    wire _7811;
    wire [15:0] _7819;
    wire [15:0] _7821;
    wire [15:0] _463;
    reg [15:0] _4111;
    wire _7828;
    wire _7825;
    wire _7826;
    wire _7829;
    wire [15:0] _7830;
    wire _7823;
    wire _7824;
    wire [15:0] _7832;
    wire [15:0] _7834;
    wire [15:0] _464;
    reg [15:0] _4108;
    wire _7841;
    wire _7838;
    wire _7839;
    wire _7842;
    wire [15:0] _7843;
    wire _7836;
    wire _7837;
    wire [15:0] _7845;
    wire [15:0] _7847;
    wire [15:0] _465;
    reg [15:0] _4105;
    wire _7854;
    wire _7851;
    wire _7852;
    wire _7855;
    wire [15:0] _7856;
    wire _7849;
    wire _7850;
    wire [15:0] _7858;
    wire [15:0] _7860;
    wire [15:0] _466;
    reg [15:0] _4102;
    wire _7867;
    wire _7864;
    wire _7865;
    wire _7868;
    wire [15:0] _7869;
    wire _7862;
    wire _7863;
    wire [15:0] _7871;
    wire [15:0] _7873;
    wire [15:0] _467;
    reg [15:0] _4099;
    wire _7880;
    wire _7877;
    wire _7878;
    wire _7881;
    wire [15:0] _7882;
    wire _7875;
    wire _7876;
    wire [15:0] _7884;
    wire [15:0] _7886;
    wire [15:0] _468;
    reg [15:0] _4096;
    wire _7893;
    wire _7890;
    wire _7891;
    wire _7894;
    wire [15:0] _7895;
    wire _7888;
    wire _7889;
    wire [15:0] _7897;
    wire [15:0] _7899;
    wire [15:0] _469;
    reg [15:0] _4093;
    wire _7906;
    wire _7903;
    wire _7904;
    wire _7907;
    wire [15:0] _7908;
    wire _7901;
    wire _7902;
    wire [15:0] _7910;
    wire [15:0] _7912;
    wire [15:0] _470;
    reg [15:0] _4090;
    wire _7919;
    wire _7916;
    wire _7917;
    wire _7920;
    wire [15:0] _7921;
    wire _7914;
    wire _7915;
    wire [15:0] _7923;
    wire [15:0] _7925;
    wire [15:0] _471;
    reg [15:0] _4087;
    wire _7932;
    wire _7929;
    wire _7930;
    wire _7933;
    wire [15:0] _7934;
    wire _7927;
    wire _7928;
    wire [15:0] _7936;
    wire [15:0] _7938;
    wire [15:0] _472;
    reg [15:0] _4084;
    wire _7945;
    wire _7942;
    wire _7943;
    wire _7946;
    wire [15:0] _7947;
    wire _7940;
    wire _7941;
    wire [15:0] _7949;
    wire [15:0] _7951;
    wire [15:0] _473;
    reg [15:0] _4081;
    wire _7958;
    wire _7955;
    wire _7956;
    wire _7959;
    wire [15:0] _7960;
    wire _7953;
    wire _7954;
    wire [15:0] _7962;
    wire [15:0] _7964;
    wire [15:0] _474;
    reg [15:0] _4078;
    wire _7971;
    wire _7968;
    wire _7969;
    wire _7972;
    wire [15:0] _7973;
    wire _7966;
    wire _7967;
    wire [15:0] _7975;
    wire [15:0] _7977;
    wire [15:0] _475;
    reg [15:0] _4075;
    wire _7984;
    wire _7981;
    wire _7982;
    wire _7985;
    wire [15:0] _7986;
    wire _7979;
    wire _7980;
    wire [15:0] _7988;
    wire [15:0] _7990;
    wire [15:0] _476;
    reg [15:0] _4072;
    wire _7997;
    wire _7994;
    wire _7995;
    wire _7998;
    wire [15:0] _7999;
    wire _7992;
    wire _7993;
    wire [15:0] _8001;
    wire [15:0] _8003;
    wire [15:0] _477;
    reg [15:0] _4069;
    wire _8010;
    wire _8007;
    wire _8008;
    wire _8011;
    wire [15:0] _8012;
    wire _8005;
    wire _8006;
    wire [15:0] _8014;
    wire [15:0] _8016;
    wire [15:0] _478;
    reg [15:0] _4066;
    wire _8023;
    wire _8020;
    wire _8021;
    wire _8024;
    wire [15:0] _8025;
    wire _8018;
    wire _8019;
    wire [15:0] _8027;
    wire [15:0] _8029;
    wire [15:0] _479;
    reg [15:0] _4063;
    wire _8036;
    wire _8033;
    wire _8034;
    wire _8037;
    wire [15:0] _8038;
    wire _8031;
    wire _8032;
    wire [15:0] _8040;
    wire [15:0] _8042;
    wire [15:0] _480;
    reg [15:0] _4060;
    wire _8049;
    wire _8046;
    wire _8047;
    wire _8050;
    wire [15:0] _8051;
    wire _8044;
    wire _8045;
    wire [15:0] _8053;
    wire [15:0] _8055;
    wire [15:0] _481;
    reg [15:0] _4057;
    wire _8062;
    wire _8059;
    wire _8060;
    wire _8063;
    wire [15:0] _8064;
    wire _8057;
    wire _8058;
    wire [15:0] _8066;
    wire [15:0] _8068;
    wire [15:0] _482;
    reg [15:0] _4054;
    wire _8075;
    wire _8072;
    wire _8073;
    wire _8076;
    wire [15:0] _8077;
    wire _8070;
    wire _8071;
    wire [15:0] _8079;
    wire [15:0] _8081;
    wire [15:0] _483;
    reg [15:0] _4051;
    wire _8088;
    wire _8085;
    wire _8086;
    wire _8089;
    wire [15:0] _8090;
    wire _8083;
    wire _8084;
    wire [15:0] _8092;
    wire [15:0] _8094;
    wire [15:0] _484;
    reg [15:0] _4048;
    wire _8101;
    wire _8098;
    wire _8099;
    wire _8102;
    wire [15:0] _8103;
    wire _8096;
    wire _8097;
    wire [15:0] _8105;
    wire [15:0] _8107;
    wire [15:0] _485;
    reg [15:0] _4045;
    wire _8114;
    wire _8111;
    wire _8112;
    wire _8115;
    wire [15:0] _8116;
    wire _8109;
    wire _8110;
    wire [15:0] _8118;
    wire [15:0] _8120;
    wire [15:0] _486;
    reg [15:0] _4042;
    wire _8127;
    wire _8124;
    wire _8125;
    wire _8128;
    wire [15:0] _8129;
    wire _8122;
    wire _8123;
    wire [15:0] _8131;
    wire [15:0] _8133;
    wire [15:0] _487;
    reg [15:0] _4039;
    wire _8140;
    wire _8137;
    wire _8138;
    wire _8141;
    wire [15:0] _8142;
    wire _8135;
    wire _8136;
    wire [15:0] _8144;
    wire [15:0] _8146;
    wire [15:0] _488;
    reg [15:0] _4036;
    wire _8153;
    wire _8150;
    wire _8151;
    wire _8154;
    wire [15:0] _8155;
    wire _8148;
    wire _8149;
    wire [15:0] _8157;
    wire [15:0] _8159;
    wire [15:0] _489;
    reg [15:0] _4033;
    wire _8166;
    wire _8163;
    wire _8164;
    wire _8167;
    wire [15:0] _8168;
    wire _8161;
    wire _8162;
    wire [15:0] _8170;
    wire [15:0] _8172;
    wire [15:0] _490;
    reg [15:0] _4030;
    wire _8179;
    wire _8176;
    wire _8177;
    wire _8180;
    wire [15:0] _8181;
    wire _8174;
    wire _8175;
    wire [15:0] _8183;
    wire [15:0] _8185;
    wire [15:0] _491;
    reg [15:0] _4027;
    wire _8192;
    wire _8189;
    wire _8190;
    wire _8193;
    wire [15:0] _8194;
    wire _8187;
    wire _8188;
    wire [15:0] _8196;
    wire [15:0] _8198;
    wire [15:0] _492;
    reg [15:0] _4024;
    wire _8205;
    wire _8202;
    wire _8203;
    wire _8206;
    wire [15:0] _8207;
    wire _8200;
    wire _8201;
    wire [15:0] _8209;
    wire [15:0] _8211;
    wire [15:0] _493;
    reg [15:0] _4021;
    wire _8218;
    wire _8215;
    wire _8216;
    wire _8219;
    wire [15:0] _8220;
    wire _8213;
    wire _8214;
    wire [15:0] _8222;
    wire [15:0] _8224;
    wire [15:0] _494;
    reg [15:0] _4018;
    wire _8231;
    wire _8228;
    wire _8229;
    wire _8232;
    wire [15:0] _8233;
    wire _8226;
    wire _8227;
    wire [15:0] _8235;
    wire [15:0] _8237;
    wire [15:0] _495;
    reg [15:0] _4015;
    wire _8244;
    wire _8241;
    wire _8242;
    wire _8245;
    wire [15:0] _8246;
    wire _8239;
    wire _8240;
    wire [15:0] _8248;
    wire [15:0] _8250;
    wire [15:0] _496;
    reg [15:0] _4012;
    wire _8257;
    wire _8254;
    wire _8255;
    wire _8258;
    wire [15:0] _8259;
    wire _8252;
    wire _8253;
    wire [15:0] _8261;
    wire [15:0] _8263;
    wire [15:0] _497;
    reg [15:0] _4009;
    wire _8270;
    wire _8267;
    wire _8268;
    wire _8271;
    wire [15:0] _8272;
    wire _8265;
    wire _8266;
    wire [15:0] _8274;
    wire [15:0] _8276;
    wire [15:0] _498;
    reg [15:0] _4006;
    wire _8283;
    wire _8280;
    wire _8281;
    wire _8284;
    wire [15:0] _8285;
    wire _8278;
    wire _8279;
    wire [15:0] _8287;
    wire [15:0] _8289;
    wire [15:0] _499;
    reg [15:0] _4003;
    wire _8296;
    wire _8293;
    wire _8294;
    wire _8297;
    wire [15:0] _8298;
    wire _8291;
    wire _8292;
    wire [15:0] _8300;
    wire [15:0] _8302;
    wire [15:0] _500;
    reg [15:0] _4000;
    wire _8309;
    wire _8306;
    wire _8307;
    wire _8310;
    wire [15:0] _8311;
    wire _8304;
    wire _8305;
    wire [15:0] _8313;
    wire [15:0] _8315;
    wire [15:0] _501;
    reg [15:0] _3997;
    wire _8322;
    wire _8319;
    wire _8320;
    wire _8323;
    wire [15:0] _8324;
    wire _8317;
    wire _8318;
    wire [15:0] _8326;
    wire [15:0] _8328;
    wire [15:0] _502;
    reg [15:0] _3994;
    wire _8335;
    wire _8332;
    wire _8333;
    wire _8336;
    wire [15:0] _8337;
    wire _8330;
    wire _8331;
    wire [15:0] _8339;
    wire [15:0] _8341;
    wire [15:0] _503;
    reg [15:0] _3991;
    wire _8348;
    wire _8345;
    wire _8346;
    wire _8349;
    wire [15:0] _8350;
    wire _8343;
    wire _8344;
    wire [15:0] _8352;
    wire [15:0] _8354;
    wire [15:0] _504;
    reg [15:0] _3988;
    wire _8361;
    wire _8358;
    wire _8359;
    wire _8362;
    wire [15:0] _8363;
    wire _8356;
    wire _8357;
    wire [15:0] _8365;
    wire [15:0] _8367;
    wire [15:0] _505;
    reg [15:0] _3985;
    wire _8374;
    wire _8371;
    wire _8372;
    wire _8375;
    wire [15:0] _8376;
    wire _8369;
    wire _8370;
    wire [15:0] _8378;
    wire [15:0] _8380;
    wire [15:0] _506;
    reg [15:0] _3982;
    wire _8387;
    wire _8384;
    wire _8385;
    wire _8388;
    wire [15:0] _8389;
    wire _8382;
    wire _8383;
    wire [15:0] _8391;
    wire [15:0] _8393;
    wire [15:0] _507;
    reg [15:0] _3979;
    wire _8400;
    wire _8397;
    wire _8398;
    wire _8401;
    wire [15:0] _8402;
    wire _8395;
    wire _8396;
    wire [15:0] _8404;
    wire [15:0] _8406;
    wire [15:0] _508;
    reg [15:0] _3976;
    wire _8413;
    wire _8410;
    wire _8411;
    wire _8414;
    wire [15:0] _8415;
    wire _8408;
    wire _8409;
    wire [15:0] _8417;
    wire [15:0] _8419;
    wire [15:0] _509;
    reg [15:0] _3973;
    wire _8426;
    wire _8423;
    wire _8424;
    wire _8427;
    wire [15:0] _8428;
    wire _8421;
    wire _8422;
    wire [15:0] _8430;
    wire [15:0] _8432;
    wire [15:0] _510;
    reg [15:0] _3970;
    wire _8439;
    wire _8436;
    wire _8437;
    wire _8440;
    wire [15:0] _8441;
    wire _8434;
    wire _8435;
    wire [15:0] _8443;
    wire [15:0] _8445;
    wire [15:0] _511;
    reg [15:0] _3967;
    wire _8452;
    wire _8449;
    wire _8450;
    wire _8453;
    wire [15:0] _8454;
    wire _8447;
    wire _8448;
    wire [15:0] _8456;
    wire [15:0] _8458;
    wire [15:0] _512;
    reg [15:0] _3964;
    wire _8465;
    wire _8462;
    wire _8463;
    wire _8466;
    wire [15:0] _8467;
    wire _8460;
    wire _8461;
    wire [15:0] _8469;
    wire [15:0] _8471;
    wire [15:0] _513;
    reg [15:0] _3961;
    wire _8478;
    wire _8475;
    wire _8476;
    wire _8479;
    wire [15:0] _8480;
    wire _8473;
    wire _8474;
    wire [15:0] _8482;
    wire [15:0] _8484;
    wire [15:0] _514;
    reg [15:0] _3958;
    wire _8491;
    wire _8488;
    wire _8489;
    wire _8492;
    wire [15:0] _8493;
    wire _8486;
    wire _8487;
    wire [15:0] _8495;
    wire [15:0] _8497;
    wire [15:0] _515;
    reg [15:0] _3955;
    wire _8504;
    wire _8501;
    wire _8502;
    wire _8505;
    wire [15:0] _8506;
    wire _8499;
    wire _8500;
    wire [15:0] _8508;
    wire [15:0] _8510;
    wire [15:0] _516;
    reg [15:0] _3952;
    wire _8517;
    wire _8514;
    wire _8515;
    wire _8518;
    wire [15:0] _8519;
    wire _8512;
    wire _8513;
    wire [15:0] _8521;
    wire [15:0] _8523;
    wire [15:0] _517;
    reg [15:0] _3949;
    wire _8530;
    wire _8527;
    wire _8528;
    wire _8531;
    wire [15:0] _8532;
    wire _8525;
    wire _8526;
    wire [15:0] _8534;
    wire [15:0] _8536;
    wire [15:0] _518;
    reg [15:0] _3946;
    wire _8543;
    wire _8540;
    wire _8541;
    wire _8544;
    wire [15:0] _8545;
    wire _8538;
    wire _8539;
    wire [15:0] _8547;
    wire [15:0] _8549;
    wire [15:0] _519;
    reg [15:0] _3943;
    wire _8556;
    wire _8553;
    wire _8554;
    wire _8557;
    wire [15:0] _8558;
    wire _8551;
    wire _8552;
    wire [15:0] _8560;
    wire [15:0] _8562;
    wire [15:0] _520;
    reg [15:0] _3940;
    wire _8569;
    wire _8566;
    wire _8567;
    wire _8570;
    wire [15:0] _8571;
    wire _8564;
    wire _8565;
    wire [15:0] _8573;
    wire [15:0] _8575;
    wire [15:0] _521;
    reg [15:0] _3937;
    wire _8582;
    wire _8579;
    wire _8580;
    wire _8583;
    wire [15:0] _8584;
    wire _8577;
    wire _8578;
    wire [15:0] _8586;
    wire [15:0] _8588;
    wire [15:0] _522;
    reg [15:0] _3934;
    wire _8595;
    wire _8592;
    wire _8593;
    wire _8596;
    wire [15:0] _8597;
    wire _8590;
    wire _8591;
    wire [15:0] _8599;
    wire [15:0] _8601;
    wire [15:0] _523;
    reg [15:0] _3931;
    wire _8608;
    wire _8605;
    wire _8606;
    wire _8609;
    wire [15:0] _8610;
    wire _8603;
    wire _8604;
    wire [15:0] _8612;
    wire [15:0] _8614;
    wire [15:0] _524;
    reg [15:0] _3928;
    reg [15:0] _4692;
    wire [15:0] _4693;
    wire _8622;
    wire _8618;
    wire _8619;
    wire _8623;
    wire [7:0] _8624;
    wire _8616;
    wire _8617;
    wire [7:0] _8626;
    wire [7:0] _8628;
    wire [7:0] _525;
    reg [7:0] _3903;
    wire _8635;
    wire _8632;
    wire _8633;
    wire _8636;
    wire [7:0] _8637;
    wire _8630;
    wire _8631;
    wire [7:0] _8639;
    wire [7:0] _8641;
    wire [7:0] _526;
    reg [7:0] _3900;
    wire _8648;
    wire _8645;
    wire _8646;
    wire _8649;
    wire [7:0] _8650;
    wire _8643;
    wire _8644;
    wire [7:0] _8652;
    wire [7:0] _8654;
    wire [7:0] _527;
    reg [7:0] _3897;
    wire _8661;
    wire _8658;
    wire _8659;
    wire _8662;
    wire [7:0] _8663;
    wire _8656;
    wire _8657;
    wire [7:0] _8665;
    wire [7:0] _8667;
    wire [7:0] _528;
    reg [7:0] _3894;
    wire _8674;
    wire _8671;
    wire _8672;
    wire _8675;
    wire [7:0] _8676;
    wire _8669;
    wire _8670;
    wire [7:0] _8678;
    wire [7:0] _8680;
    wire [7:0] _529;
    reg [7:0] _3891;
    wire _8687;
    wire _8684;
    wire _8685;
    wire _8688;
    wire [7:0] _8689;
    wire _8682;
    wire _8683;
    wire [7:0] _8691;
    wire [7:0] _8693;
    wire [7:0] _530;
    reg [7:0] _3888;
    wire _8700;
    wire _8697;
    wire _8698;
    wire _8701;
    wire [7:0] _8702;
    wire _8695;
    wire _8696;
    wire [7:0] _8704;
    wire [7:0] _8706;
    wire [7:0] _531;
    reg [7:0] _3885;
    wire _8713;
    wire _8710;
    wire _8711;
    wire _8714;
    wire [7:0] _8715;
    wire _8708;
    wire _8709;
    wire [7:0] _8717;
    wire [7:0] _8719;
    wire [7:0] _532;
    reg [7:0] _3882;
    wire _8726;
    wire _8723;
    wire _8724;
    wire _8727;
    wire [7:0] _8728;
    wire _8721;
    wire _8722;
    wire [7:0] _8730;
    wire [7:0] _8732;
    wire [7:0] _533;
    reg [7:0] _3879;
    wire _8739;
    wire _8736;
    wire _8737;
    wire _8740;
    wire [7:0] _8741;
    wire _8734;
    wire _8735;
    wire [7:0] _8743;
    wire [7:0] _8745;
    wire [7:0] _534;
    reg [7:0] _3876;
    wire _8752;
    wire _8749;
    wire _8750;
    wire _8753;
    wire [7:0] _8754;
    wire _8747;
    wire _8748;
    wire [7:0] _8756;
    wire [7:0] _8758;
    wire [7:0] _535;
    reg [7:0] _3873;
    wire _8765;
    wire _8762;
    wire _8763;
    wire _8766;
    wire [7:0] _8767;
    wire _8760;
    wire _8761;
    wire [7:0] _8769;
    wire [7:0] _8771;
    wire [7:0] _536;
    reg [7:0] _3870;
    wire _8778;
    wire _8775;
    wire _8776;
    wire _8779;
    wire [7:0] _8780;
    wire _8773;
    wire _8774;
    wire [7:0] _8782;
    wire [7:0] _8784;
    wire [7:0] _537;
    reg [7:0] _3867;
    wire _8791;
    wire _8788;
    wire _8789;
    wire _8792;
    wire [7:0] _8793;
    wire _8786;
    wire _8787;
    wire [7:0] _8795;
    wire [7:0] _8797;
    wire [7:0] _538;
    reg [7:0] _3864;
    wire _8804;
    wire _8801;
    wire _8802;
    wire _8805;
    wire [7:0] _8806;
    wire _8799;
    wire _8800;
    wire [7:0] _8808;
    wire [7:0] _8810;
    wire [7:0] _539;
    reg [7:0] _3861;
    wire _8817;
    wire _8814;
    wire _8815;
    wire _8818;
    wire [7:0] _8819;
    wire _8812;
    wire _8813;
    wire [7:0] _8821;
    wire [7:0] _8823;
    wire [7:0] _540;
    reg [7:0] _3858;
    wire _8830;
    wire _8827;
    wire _8828;
    wire _8831;
    wire [7:0] _8832;
    wire _8825;
    wire _8826;
    wire [7:0] _8834;
    wire [7:0] _8836;
    wire [7:0] _541;
    reg [7:0] _3855;
    wire _8843;
    wire _8840;
    wire _8841;
    wire _8844;
    wire [7:0] _8845;
    wire _8838;
    wire _8839;
    wire [7:0] _8847;
    wire [7:0] _8849;
    wire [7:0] _542;
    reg [7:0] _3852;
    wire _8856;
    wire _8853;
    wire _8854;
    wire _8857;
    wire [7:0] _8858;
    wire _8851;
    wire _8852;
    wire [7:0] _8860;
    wire [7:0] _8862;
    wire [7:0] _543;
    reg [7:0] _3849;
    wire _8869;
    wire _8866;
    wire _8867;
    wire _8870;
    wire [7:0] _8871;
    wire _8864;
    wire _8865;
    wire [7:0] _8873;
    wire [7:0] _8875;
    wire [7:0] _544;
    reg [7:0] _3846;
    wire _8882;
    wire _8879;
    wire _8880;
    wire _8883;
    wire [7:0] _8884;
    wire _8877;
    wire _8878;
    wire [7:0] _8886;
    wire [7:0] _8888;
    wire [7:0] _545;
    reg [7:0] _3843;
    wire _8895;
    wire _8892;
    wire _8893;
    wire _8896;
    wire [7:0] _8897;
    wire _8890;
    wire _8891;
    wire [7:0] _8899;
    wire [7:0] _8901;
    wire [7:0] _546;
    reg [7:0] _3840;
    wire _8908;
    wire _8905;
    wire _8906;
    wire _8909;
    wire [7:0] _8910;
    wire _8903;
    wire _8904;
    wire [7:0] _8912;
    wire [7:0] _8914;
    wire [7:0] _547;
    reg [7:0] _3837;
    wire _8921;
    wire _8918;
    wire _8919;
    wire _8922;
    wire [7:0] _8923;
    wire _8916;
    wire _8917;
    wire [7:0] _8925;
    wire [7:0] _8927;
    wire [7:0] _548;
    reg [7:0] _3834;
    wire _8934;
    wire _8931;
    wire _8932;
    wire _8935;
    wire [7:0] _8936;
    wire _8929;
    wire _8930;
    wire [7:0] _8938;
    wire [7:0] _8940;
    wire [7:0] _549;
    reg [7:0] _3831;
    wire _8947;
    wire _8944;
    wire _8945;
    wire _8948;
    wire [7:0] _8949;
    wire _8942;
    wire _8943;
    wire [7:0] _8951;
    wire [7:0] _8953;
    wire [7:0] _550;
    reg [7:0] _3828;
    wire _8960;
    wire _8957;
    wire _8958;
    wire _8961;
    wire [7:0] _8962;
    wire _8955;
    wire _8956;
    wire [7:0] _8964;
    wire [7:0] _8966;
    wire [7:0] _551;
    reg [7:0] _3825;
    wire _8973;
    wire _8970;
    wire _8971;
    wire _8974;
    wire [7:0] _8975;
    wire _8968;
    wire _8969;
    wire [7:0] _8977;
    wire [7:0] _8979;
    wire [7:0] _552;
    reg [7:0] _3822;
    wire _8986;
    wire _8983;
    wire _8984;
    wire _8987;
    wire [7:0] _8988;
    wire _8981;
    wire _8982;
    wire [7:0] _8990;
    wire [7:0] _8992;
    wire [7:0] _553;
    reg [7:0] _3819;
    wire _8999;
    wire _8996;
    wire _8997;
    wire _9000;
    wire [7:0] _9001;
    wire _8994;
    wire _8995;
    wire [7:0] _9003;
    wire [7:0] _9005;
    wire [7:0] _554;
    reg [7:0] _3816;
    wire _9012;
    wire _9009;
    wire _9010;
    wire _9013;
    wire [7:0] _9014;
    wire _9007;
    wire _9008;
    wire [7:0] _9016;
    wire [7:0] _9018;
    wire [7:0] _555;
    reg [7:0] _3813;
    wire _9025;
    wire _9022;
    wire _9023;
    wire _9026;
    wire [7:0] _9027;
    wire _9020;
    wire _9021;
    wire [7:0] _9029;
    wire [7:0] _9031;
    wire [7:0] _556;
    reg [7:0] _3810;
    wire _9038;
    wire _9035;
    wire _9036;
    wire _9039;
    wire [7:0] _9040;
    wire _9033;
    wire _9034;
    wire [7:0] _9042;
    wire [7:0] _9044;
    wire [7:0] _557;
    reg [7:0] _3807;
    wire _9051;
    wire _9048;
    wire _9049;
    wire _9052;
    wire [7:0] _9053;
    wire _9046;
    wire _9047;
    wire [7:0] _9055;
    wire [7:0] _9057;
    wire [7:0] _558;
    reg [7:0] _3804;
    wire _9064;
    wire _9061;
    wire _9062;
    wire _9065;
    wire [7:0] _9066;
    wire _9059;
    wire _9060;
    wire [7:0] _9068;
    wire [7:0] _9070;
    wire [7:0] _559;
    reg [7:0] _3801;
    wire _9077;
    wire _9074;
    wire _9075;
    wire _9078;
    wire [7:0] _9079;
    wire _9072;
    wire _9073;
    wire [7:0] _9081;
    wire [7:0] _9083;
    wire [7:0] _560;
    reg [7:0] _3798;
    wire _9090;
    wire _9087;
    wire _9088;
    wire _9091;
    wire [7:0] _9092;
    wire _9085;
    wire _9086;
    wire [7:0] _9094;
    wire [7:0] _9096;
    wire [7:0] _561;
    reg [7:0] _3795;
    wire _9103;
    wire _9100;
    wire _9101;
    wire _9104;
    wire [7:0] _9105;
    wire _9098;
    wire _9099;
    wire [7:0] _9107;
    wire [7:0] _9109;
    wire [7:0] _562;
    reg [7:0] _3792;
    wire _9116;
    wire _9113;
    wire _9114;
    wire _9117;
    wire [7:0] _9118;
    wire _9111;
    wire _9112;
    wire [7:0] _9120;
    wire [7:0] _9122;
    wire [7:0] _563;
    reg [7:0] _3789;
    wire _9129;
    wire _9126;
    wire _9127;
    wire _9130;
    wire [7:0] _9131;
    wire _9124;
    wire _9125;
    wire [7:0] _9133;
    wire [7:0] _9135;
    wire [7:0] _564;
    reg [7:0] _3786;
    wire _9142;
    wire _9139;
    wire _9140;
    wire _9143;
    wire [7:0] _9144;
    wire _9137;
    wire _9138;
    wire [7:0] _9146;
    wire [7:0] _9148;
    wire [7:0] _565;
    reg [7:0] _3783;
    wire _9155;
    wire _9152;
    wire _9153;
    wire _9156;
    wire [7:0] _9157;
    wire _9150;
    wire _9151;
    wire [7:0] _9159;
    wire [7:0] _9161;
    wire [7:0] _566;
    reg [7:0] _3780;
    wire _9168;
    wire _9165;
    wire _9166;
    wire _9169;
    wire [7:0] _9170;
    wire _9163;
    wire _9164;
    wire [7:0] _9172;
    wire [7:0] _9174;
    wire [7:0] _567;
    reg [7:0] _3777;
    wire _9181;
    wire _9178;
    wire _9179;
    wire _9182;
    wire [7:0] _9183;
    wire _9176;
    wire _9177;
    wire [7:0] _9185;
    wire [7:0] _9187;
    wire [7:0] _568;
    reg [7:0] _3774;
    wire _9194;
    wire _9191;
    wire _9192;
    wire _9195;
    wire [7:0] _9196;
    wire _9189;
    wire _9190;
    wire [7:0] _9198;
    wire [7:0] _9200;
    wire [7:0] _569;
    reg [7:0] _3771;
    wire _9207;
    wire _9204;
    wire _9205;
    wire _9208;
    wire [7:0] _9209;
    wire _9202;
    wire _9203;
    wire [7:0] _9211;
    wire [7:0] _9213;
    wire [7:0] _570;
    reg [7:0] _3768;
    wire _9220;
    wire _9217;
    wire _9218;
    wire _9221;
    wire [7:0] _9222;
    wire _9215;
    wire _9216;
    wire [7:0] _9224;
    wire [7:0] _9226;
    wire [7:0] _571;
    reg [7:0] _3765;
    wire _9233;
    wire _9230;
    wire _9231;
    wire _9234;
    wire [7:0] _9235;
    wire _9228;
    wire _9229;
    wire [7:0] _9237;
    wire [7:0] _9239;
    wire [7:0] _572;
    reg [7:0] _3762;
    wire _9246;
    wire _9243;
    wire _9244;
    wire _9247;
    wire [7:0] _9248;
    wire _9241;
    wire _9242;
    wire [7:0] _9250;
    wire [7:0] _9252;
    wire [7:0] _573;
    reg [7:0] _3759;
    wire _9259;
    wire _9256;
    wire _9257;
    wire _9260;
    wire [7:0] _9261;
    wire _9254;
    wire _9255;
    wire [7:0] _9263;
    wire [7:0] _9265;
    wire [7:0] _574;
    reg [7:0] _3756;
    wire _9272;
    wire _9269;
    wire _9270;
    wire _9273;
    wire [7:0] _9274;
    wire _9267;
    wire _9268;
    wire [7:0] _9276;
    wire [7:0] _9278;
    wire [7:0] _575;
    reg [7:0] _3753;
    wire _9285;
    wire _9282;
    wire _9283;
    wire _9286;
    wire [7:0] _9287;
    wire _9280;
    wire _9281;
    wire [7:0] _9289;
    wire [7:0] _9291;
    wire [7:0] _576;
    reg [7:0] _3750;
    wire _9298;
    wire _9295;
    wire _9296;
    wire _9299;
    wire [7:0] _9300;
    wire _9293;
    wire _9294;
    wire [7:0] _9302;
    wire [7:0] _9304;
    wire [7:0] _577;
    reg [7:0] _3747;
    wire _9311;
    wire _9308;
    wire _9309;
    wire _9312;
    wire [7:0] _9313;
    wire _9306;
    wire _9307;
    wire [7:0] _9315;
    wire [7:0] _9317;
    wire [7:0] _578;
    reg [7:0] _3744;
    wire _9324;
    wire _9321;
    wire _9322;
    wire _9325;
    wire [7:0] _9326;
    wire _9319;
    wire _9320;
    wire [7:0] _9328;
    wire [7:0] _9330;
    wire [7:0] _579;
    reg [7:0] _3741;
    wire _9337;
    wire _9334;
    wire _9335;
    wire _9338;
    wire [7:0] _9339;
    wire _9332;
    wire _9333;
    wire [7:0] _9341;
    wire [7:0] _9343;
    wire [7:0] _580;
    reg [7:0] _3738;
    wire _9350;
    wire _9347;
    wire _9348;
    wire _9351;
    wire [7:0] _9352;
    wire _9345;
    wire _9346;
    wire [7:0] _9354;
    wire [7:0] _9356;
    wire [7:0] _581;
    reg [7:0] _3735;
    wire _9363;
    wire _9360;
    wire _9361;
    wire _9364;
    wire [7:0] _9365;
    wire _9358;
    wire _9359;
    wire [7:0] _9367;
    wire [7:0] _9369;
    wire [7:0] _582;
    reg [7:0] _3732;
    wire _9376;
    wire _9373;
    wire _9374;
    wire _9377;
    wire [7:0] _9378;
    wire _9371;
    wire _9372;
    wire [7:0] _9380;
    wire [7:0] _9382;
    wire [7:0] _583;
    reg [7:0] _3729;
    wire _9389;
    wire _9386;
    wire _9387;
    wire _9390;
    wire [7:0] _9391;
    wire _9384;
    wire _9385;
    wire [7:0] _9393;
    wire [7:0] _9395;
    wire [7:0] _584;
    reg [7:0] _3726;
    wire _9402;
    wire _9399;
    wire _9400;
    wire _9403;
    wire [7:0] _9404;
    wire _9397;
    wire _9398;
    wire [7:0] _9406;
    wire [7:0] _9408;
    wire [7:0] _585;
    reg [7:0] _3723;
    wire _9415;
    wire _9412;
    wire _9413;
    wire _9416;
    wire [7:0] _9417;
    wire _9410;
    wire _9411;
    wire [7:0] _9419;
    wire [7:0] _9421;
    wire [7:0] _586;
    reg [7:0] _3720;
    wire _9428;
    wire _9425;
    wire _9426;
    wire _9429;
    wire [7:0] _9430;
    wire _9423;
    wire _9424;
    wire [7:0] _9432;
    wire [7:0] _9434;
    wire [7:0] _587;
    reg [7:0] _3717;
    wire _9441;
    wire _9438;
    wire _9439;
    wire _9442;
    wire [7:0] _9443;
    wire _9436;
    wire _9437;
    wire [7:0] _9445;
    wire [7:0] _9447;
    wire [7:0] _588;
    reg [7:0] _3714;
    wire _9454;
    wire _9451;
    wire _9452;
    wire _9455;
    wire [7:0] _9456;
    wire _9449;
    wire _9450;
    wire [7:0] _9458;
    wire [7:0] _9460;
    wire [7:0] _589;
    reg [7:0] _3711;
    wire _9467;
    wire _9464;
    wire _9465;
    wire _9468;
    wire [7:0] _9469;
    wire _9462;
    wire _9463;
    wire [7:0] _9471;
    wire [7:0] _9473;
    wire [7:0] _590;
    reg [7:0] _3708;
    wire _9480;
    wire _9477;
    wire _9478;
    wire _9481;
    wire [7:0] _9482;
    wire _9475;
    wire _9476;
    wire [7:0] _9484;
    wire [7:0] _9486;
    wire [7:0] _591;
    reg [7:0] _3705;
    wire _9493;
    wire _9490;
    wire _9491;
    wire _9494;
    wire [7:0] _9495;
    wire _9488;
    wire _9489;
    wire [7:0] _9497;
    wire [7:0] _9499;
    wire [7:0] _592;
    reg [7:0] _3702;
    wire _9506;
    wire _9503;
    wire _9504;
    wire _9507;
    wire [7:0] _9508;
    wire _9501;
    wire _9502;
    wire [7:0] _9510;
    wire [7:0] _9512;
    wire [7:0] _593;
    reg [7:0] _3699;
    wire _9519;
    wire _9516;
    wire _9517;
    wire _9520;
    wire [7:0] _9521;
    wire _9514;
    wire _9515;
    wire [7:0] _9523;
    wire [7:0] _9525;
    wire [7:0] _594;
    reg [7:0] _3696;
    wire _9532;
    wire _9529;
    wire _9530;
    wire _9533;
    wire [7:0] _9534;
    wire _9527;
    wire _9528;
    wire [7:0] _9536;
    wire [7:0] _9538;
    wire [7:0] _595;
    reg [7:0] _3693;
    wire _9545;
    wire _9542;
    wire _9543;
    wire _9546;
    wire [7:0] _9547;
    wire _9540;
    wire _9541;
    wire [7:0] _9549;
    wire [7:0] _9551;
    wire [7:0] _596;
    reg [7:0] _3690;
    wire _9558;
    wire _9555;
    wire _9556;
    wire _9559;
    wire [7:0] _9560;
    wire _9553;
    wire _9554;
    wire [7:0] _9562;
    wire [7:0] _9564;
    wire [7:0] _597;
    reg [7:0] _3687;
    wire _9571;
    wire _9568;
    wire _9569;
    wire _9572;
    wire [7:0] _9573;
    wire _9566;
    wire _9567;
    wire [7:0] _9575;
    wire [7:0] _9577;
    wire [7:0] _598;
    reg [7:0] _3684;
    wire _9584;
    wire _9581;
    wire _9582;
    wire _9585;
    wire [7:0] _9586;
    wire _9579;
    wire _9580;
    wire [7:0] _9588;
    wire [7:0] _9590;
    wire [7:0] _599;
    reg [7:0] _3681;
    wire _9597;
    wire _9594;
    wire _9595;
    wire _9598;
    wire [7:0] _9599;
    wire _9592;
    wire _9593;
    wire [7:0] _9601;
    wire [7:0] _9603;
    wire [7:0] _600;
    reg [7:0] _3678;
    wire _9610;
    wire _9607;
    wire _9608;
    wire _9611;
    wire [7:0] _9612;
    wire _9605;
    wire _9606;
    wire [7:0] _9614;
    wire [7:0] _9616;
    wire [7:0] _601;
    reg [7:0] _3675;
    wire _9623;
    wire _9620;
    wire _9621;
    wire _9624;
    wire [7:0] _9625;
    wire _9618;
    wire _9619;
    wire [7:0] _9627;
    wire [7:0] _9629;
    wire [7:0] _602;
    reg [7:0] _3672;
    wire _9636;
    wire _9633;
    wire _9634;
    wire _9637;
    wire [7:0] _9638;
    wire _9631;
    wire _9632;
    wire [7:0] _9640;
    wire [7:0] _9642;
    wire [7:0] _603;
    reg [7:0] _3669;
    wire _9649;
    wire _9646;
    wire _9647;
    wire _9650;
    wire [7:0] _9651;
    wire _9644;
    wire _9645;
    wire [7:0] _9653;
    wire [7:0] _9655;
    wire [7:0] _604;
    reg [7:0] _3666;
    wire _9662;
    wire _9659;
    wire _9660;
    wire _9663;
    wire [7:0] _9664;
    wire _9657;
    wire _9658;
    wire [7:0] _9666;
    wire [7:0] _9668;
    wire [7:0] _605;
    reg [7:0] _3663;
    wire _9675;
    wire _9672;
    wire _9673;
    wire _9676;
    wire [7:0] _9677;
    wire _9670;
    wire _9671;
    wire [7:0] _9679;
    wire [7:0] _9681;
    wire [7:0] _606;
    reg [7:0] _3660;
    wire _9688;
    wire _9685;
    wire _9686;
    wire _9689;
    wire [7:0] _9690;
    wire _9683;
    wire _9684;
    wire [7:0] _9692;
    wire [7:0] _9694;
    wire [7:0] _607;
    reg [7:0] _3657;
    wire _9701;
    wire _9698;
    wire _9699;
    wire _9702;
    wire [7:0] _9703;
    wire _9696;
    wire _9697;
    wire [7:0] _9705;
    wire [7:0] _9707;
    wire [7:0] _608;
    reg [7:0] _3654;
    wire _9714;
    wire _9711;
    wire _9712;
    wire _9715;
    wire [7:0] _9716;
    wire _9709;
    wire _9710;
    wire [7:0] _9718;
    wire [7:0] _9720;
    wire [7:0] _609;
    reg [7:0] _3651;
    wire _9727;
    wire _9724;
    wire _9725;
    wire _9728;
    wire [7:0] _9729;
    wire _9722;
    wire _9723;
    wire [7:0] _9731;
    wire [7:0] _9733;
    wire [7:0] _610;
    reg [7:0] _3648;
    wire _9740;
    wire _9737;
    wire _9738;
    wire _9741;
    wire [7:0] _9742;
    wire _9735;
    wire _9736;
    wire [7:0] _9744;
    wire [7:0] _9746;
    wire [7:0] _611;
    reg [7:0] _3645;
    wire _9753;
    wire _9750;
    wire _9751;
    wire _9754;
    wire [7:0] _9755;
    wire _9748;
    wire _9749;
    wire [7:0] _9757;
    wire [7:0] _9759;
    wire [7:0] _612;
    reg [7:0] _3642;
    wire _9766;
    wire _9763;
    wire _9764;
    wire _9767;
    wire [7:0] _9768;
    wire _9761;
    wire _9762;
    wire [7:0] _9770;
    wire [7:0] _9772;
    wire [7:0] _613;
    reg [7:0] _3639;
    wire _9779;
    wire _9776;
    wire _9777;
    wire _9780;
    wire [7:0] _9781;
    wire _9774;
    wire _9775;
    wire [7:0] _9783;
    wire [7:0] _9785;
    wire [7:0] _614;
    reg [7:0] _3636;
    wire _9792;
    wire _9789;
    wire _9790;
    wire _9793;
    wire [7:0] _9794;
    wire _9787;
    wire _9788;
    wire [7:0] _9796;
    wire [7:0] _9798;
    wire [7:0] _615;
    reg [7:0] _3633;
    wire _9805;
    wire _9802;
    wire _9803;
    wire _9806;
    wire [7:0] _9807;
    wire _9800;
    wire _9801;
    wire [7:0] _9809;
    wire [7:0] _9811;
    wire [7:0] _616;
    reg [7:0] _3630;
    wire _9818;
    wire _9815;
    wire _9816;
    wire _9819;
    wire [7:0] _9820;
    wire _9813;
    wire _9814;
    wire [7:0] _9822;
    wire [7:0] _9824;
    wire [7:0] _617;
    reg [7:0] _3627;
    wire _9831;
    wire _9828;
    wire _9829;
    wire _9832;
    wire [7:0] _9833;
    wire _9826;
    wire _9827;
    wire [7:0] _9835;
    wire [7:0] _9837;
    wire [7:0] _618;
    reg [7:0] _3624;
    wire _9844;
    wire _9841;
    wire _9842;
    wire _9845;
    wire [7:0] _9846;
    wire _9839;
    wire _9840;
    wire [7:0] _9848;
    wire [7:0] _9850;
    wire [7:0] _619;
    reg [7:0] _3621;
    wire _9857;
    wire _9854;
    wire _9855;
    wire _9858;
    wire [7:0] _9859;
    wire _9852;
    wire _9853;
    wire [7:0] _9861;
    wire [7:0] _9863;
    wire [7:0] _620;
    reg [7:0] _3618;
    wire _9870;
    wire _9867;
    wire _9868;
    wire _9871;
    wire [7:0] _9872;
    wire _9865;
    wire _9866;
    wire [7:0] _9874;
    wire [7:0] _9876;
    wire [7:0] _621;
    reg [7:0] _3615;
    wire _9883;
    wire _9880;
    wire _9881;
    wire _9884;
    wire [7:0] _9885;
    wire _9878;
    wire _9879;
    wire [7:0] _9887;
    wire [7:0] _9889;
    wire [7:0] _622;
    reg [7:0] _3612;
    wire _9896;
    wire _9893;
    wire _9894;
    wire _9897;
    wire [7:0] _9898;
    wire _9891;
    wire _9892;
    wire [7:0] _9900;
    wire [7:0] _9902;
    wire [7:0] _623;
    reg [7:0] _3609;
    wire _9909;
    wire _9906;
    wire _9907;
    wire _9910;
    wire [7:0] _9911;
    wire _9904;
    wire _9905;
    wire [7:0] _9913;
    wire [7:0] _9915;
    wire [7:0] _624;
    reg [7:0] _3606;
    wire _9922;
    wire _9919;
    wire _9920;
    wire _9923;
    wire [7:0] _9924;
    wire _9917;
    wire _9918;
    wire [7:0] _9926;
    wire [7:0] _9928;
    wire [7:0] _625;
    reg [7:0] _3603;
    wire _9935;
    wire _9932;
    wire _9933;
    wire _9936;
    wire [7:0] _9937;
    wire _9930;
    wire _9931;
    wire [7:0] _9939;
    wire [7:0] _9941;
    wire [7:0] _626;
    reg [7:0] _3600;
    wire _9948;
    wire _9945;
    wire _9946;
    wire _9949;
    wire [7:0] _9950;
    wire _9943;
    wire _9944;
    wire [7:0] _9952;
    wire [7:0] _9954;
    wire [7:0] _627;
    reg [7:0] _3597;
    wire _9961;
    wire _9958;
    wire _9959;
    wire _9962;
    wire [7:0] _9963;
    wire _9956;
    wire _9957;
    wire [7:0] _9965;
    wire [7:0] _9967;
    wire [7:0] _628;
    reg [7:0] _3594;
    wire _9974;
    wire _9971;
    wire _9972;
    wire _9975;
    wire [7:0] _9976;
    wire _9969;
    wire _9970;
    wire [7:0] _9978;
    wire [7:0] _9980;
    wire [7:0] _629;
    reg [7:0] _3591;
    wire _9987;
    wire _9984;
    wire _9985;
    wire _9988;
    wire [7:0] _9989;
    wire _9982;
    wire _9983;
    wire [7:0] _9991;
    wire [7:0] _9993;
    wire [7:0] _630;
    reg [7:0] _3588;
    wire _10000;
    wire _9997;
    wire _9998;
    wire _10001;
    wire [7:0] _10002;
    wire _9995;
    wire _9996;
    wire [7:0] _10004;
    wire [7:0] _10006;
    wire [7:0] _631;
    reg [7:0] _3585;
    wire _10013;
    wire _10010;
    wire _10011;
    wire _10014;
    wire [7:0] _10015;
    wire _10008;
    wire _10009;
    wire [7:0] _10017;
    wire [7:0] _10019;
    wire [7:0] _632;
    reg [7:0] _3582;
    wire _10026;
    wire _10023;
    wire _10024;
    wire _10027;
    wire [7:0] _10028;
    wire _10021;
    wire _10022;
    wire [7:0] _10030;
    wire [7:0] _10032;
    wire [7:0] _633;
    reg [7:0] _3579;
    wire _10039;
    wire _10036;
    wire _10037;
    wire _10040;
    wire [7:0] _10041;
    wire _10034;
    wire _10035;
    wire [7:0] _10043;
    wire [7:0] _10045;
    wire [7:0] _634;
    reg [7:0] _3576;
    wire _10052;
    wire _10049;
    wire _10050;
    wire _10053;
    wire [7:0] _10054;
    wire _10047;
    wire _10048;
    wire [7:0] _10056;
    wire [7:0] _10058;
    wire [7:0] _635;
    reg [7:0] _3573;
    wire _10065;
    wire _10062;
    wire _10063;
    wire _10066;
    wire [7:0] _10067;
    wire _10060;
    wire _10061;
    wire [7:0] _10069;
    wire [7:0] _10071;
    wire [7:0] _636;
    reg [7:0] _3570;
    wire _10078;
    wire _10075;
    wire _10076;
    wire _10079;
    wire [7:0] _10080;
    wire _10073;
    wire _10074;
    wire [7:0] _10082;
    wire [7:0] _10084;
    wire [7:0] _637;
    reg [7:0] _3567;
    wire _10091;
    wire _10088;
    wire _10089;
    wire _10092;
    wire [7:0] _10093;
    wire _10086;
    wire _10087;
    wire [7:0] _10095;
    wire [7:0] _10097;
    wire [7:0] _638;
    reg [7:0] _3564;
    wire _10104;
    wire _10101;
    wire _10102;
    wire _10105;
    wire [7:0] _10106;
    wire _10099;
    wire _10100;
    wire [7:0] _10108;
    wire [7:0] _10110;
    wire [7:0] _639;
    reg [7:0] _3561;
    wire _10117;
    wire _10114;
    wire _10115;
    wire _10118;
    wire [7:0] _10119;
    wire _10112;
    wire _10113;
    wire [7:0] _10121;
    wire [7:0] _10123;
    wire [7:0] _640;
    reg [7:0] _3558;
    wire _10130;
    wire _10127;
    wire _10128;
    wire _10131;
    wire [7:0] _10132;
    wire _10125;
    wire _10126;
    wire [7:0] _10134;
    wire [7:0] _10136;
    wire [7:0] _641;
    reg [7:0] _3555;
    wire _10143;
    wire _10140;
    wire _10141;
    wire _10144;
    wire [7:0] _10145;
    wire _10138;
    wire _10139;
    wire [7:0] _10147;
    wire [7:0] _10149;
    wire [7:0] _642;
    reg [7:0] _3552;
    wire _10156;
    wire _10153;
    wire _10154;
    wire _10157;
    wire [7:0] _10158;
    wire _10151;
    wire _10152;
    wire [7:0] _10160;
    wire [7:0] _10162;
    wire [7:0] _643;
    reg [7:0] _3549;
    wire _10169;
    wire _10166;
    wire _10167;
    wire _10170;
    wire [7:0] _10171;
    wire _10164;
    wire _10165;
    wire [7:0] _10173;
    wire [7:0] _10175;
    wire [7:0] _644;
    reg [7:0] _3546;
    wire _10182;
    wire _10179;
    wire _10180;
    wire _10183;
    wire [7:0] _10184;
    wire _10177;
    wire _10178;
    wire [7:0] _10186;
    wire [7:0] _10188;
    wire [7:0] _645;
    reg [7:0] _3543;
    wire _10195;
    wire _10192;
    wire _10193;
    wire _10196;
    wire [7:0] _10197;
    wire _10190;
    wire _10191;
    wire [7:0] _10199;
    wire [7:0] _10201;
    wire [7:0] _646;
    reg [7:0] _3540;
    wire _10208;
    wire _10205;
    wire _10206;
    wire _10209;
    wire [7:0] _10210;
    wire _10203;
    wire _10204;
    wire [7:0] _10212;
    wire [7:0] _10214;
    wire [7:0] _647;
    reg [7:0] _3537;
    wire _10221;
    wire _10218;
    wire _10219;
    wire _10222;
    wire [7:0] _10223;
    wire _10216;
    wire _10217;
    wire [7:0] _10225;
    wire [7:0] _10227;
    wire [7:0] _648;
    reg [7:0] _3534;
    wire _10234;
    wire _10231;
    wire _10232;
    wire _10235;
    wire [7:0] _10236;
    wire _10229;
    wire _10230;
    wire [7:0] _10238;
    wire [7:0] _10240;
    wire [7:0] _649;
    reg [7:0] _3531;
    wire _10247;
    wire _10244;
    wire _10245;
    wire _10248;
    wire [7:0] _10249;
    wire _10242;
    wire _10243;
    wire [7:0] _10251;
    wire [7:0] _10253;
    wire [7:0] _650;
    reg [7:0] _3528;
    wire _10260;
    wire _10257;
    wire _10258;
    wire _10261;
    wire [7:0] _10262;
    wire _10255;
    wire _10256;
    wire [7:0] _10264;
    wire [7:0] _10266;
    wire [7:0] _651;
    reg [7:0] _3525;
    wire _10273;
    wire _10270;
    wire _10271;
    wire _10274;
    wire [7:0] _10275;
    wire _10268;
    wire _10269;
    wire [7:0] _10277;
    wire [7:0] _10279;
    wire [7:0] _652;
    reg [7:0] _3522;
    wire _10286;
    wire _10283;
    wire _10284;
    wire _10287;
    wire [7:0] _10288;
    wire _10281;
    wire _10282;
    wire [7:0] _10290;
    wire [7:0] _10292;
    wire [7:0] _653;
    reg [7:0] _3519;
    wire _10299;
    wire _10296;
    wire _10297;
    wire _10300;
    wire [7:0] _10301;
    wire _10294;
    wire _10295;
    wire [7:0] _10303;
    wire [7:0] _10305;
    wire [7:0] _654;
    reg [7:0] _3516;
    wire _10312;
    wire _10309;
    wire _10310;
    wire _10313;
    wire [7:0] _10314;
    wire _10307;
    wire _10308;
    wire [7:0] _10316;
    wire [7:0] _10318;
    wire [7:0] _655;
    reg [7:0] _3513;
    wire _10325;
    wire _10322;
    wire _10323;
    wire _10326;
    wire [7:0] _10327;
    wire _10320;
    wire _10321;
    wire [7:0] _10329;
    wire [7:0] _10331;
    wire [7:0] _656;
    reg [7:0] _3510;
    wire _10338;
    wire _10335;
    wire _10336;
    wire _10339;
    wire [7:0] _10340;
    wire _10333;
    wire _10334;
    wire [7:0] _10342;
    wire [7:0] _10344;
    wire [7:0] _657;
    reg [7:0] _3507;
    wire _10351;
    wire _10348;
    wire _10349;
    wire _10352;
    wire [7:0] _10353;
    wire _10346;
    wire _10347;
    wire [7:0] _10355;
    wire [7:0] _10357;
    wire [7:0] _658;
    reg [7:0] _3504;
    wire _10364;
    wire _10361;
    wire _10362;
    wire _10365;
    wire [7:0] _10366;
    wire _10359;
    wire _10360;
    wire [7:0] _10368;
    wire [7:0] _10370;
    wire [7:0] _659;
    reg [7:0] _3501;
    wire _10377;
    wire _10374;
    wire _10375;
    wire _10378;
    wire [7:0] _10379;
    wire _10372;
    wire _10373;
    wire [7:0] _10381;
    wire [7:0] _10383;
    wire [7:0] _660;
    reg [7:0] _3498;
    wire _10390;
    wire _10387;
    wire _10388;
    wire _10391;
    wire [7:0] _10392;
    wire _10385;
    wire _10386;
    wire [7:0] _10394;
    wire [7:0] _10396;
    wire [7:0] _661;
    reg [7:0] _3495;
    wire _10403;
    wire _10400;
    wire _10401;
    wire _10404;
    wire [7:0] _10405;
    wire _10398;
    wire _10399;
    wire [7:0] _10407;
    wire [7:0] _10409;
    wire [7:0] _662;
    reg [7:0] _3492;
    wire _10416;
    wire _10413;
    wire _10414;
    wire _10417;
    wire [7:0] _10418;
    wire _10411;
    wire _10412;
    wire [7:0] _10420;
    wire [7:0] _10422;
    wire [7:0] _663;
    reg [7:0] _3489;
    wire _10429;
    wire _10426;
    wire _10427;
    wire _10430;
    wire [7:0] _10431;
    wire _10424;
    wire _10425;
    wire [7:0] _10433;
    wire [7:0] _10435;
    wire [7:0] _664;
    reg [7:0] _3486;
    wire _10442;
    wire _10439;
    wire _10440;
    wire _10443;
    wire [7:0] _10444;
    wire _10437;
    wire _10438;
    wire [7:0] _10446;
    wire [7:0] _10448;
    wire [7:0] _665;
    reg [7:0] _3483;
    wire _10455;
    wire _10452;
    wire _10453;
    wire _10456;
    wire [7:0] _10457;
    wire _10450;
    wire _10451;
    wire [7:0] _10459;
    wire [7:0] _10461;
    wire [7:0] _666;
    reg [7:0] _3480;
    wire _10468;
    wire _10465;
    wire _10466;
    wire _10469;
    wire [7:0] _10470;
    wire _10463;
    wire _10464;
    wire [7:0] _10472;
    wire [7:0] _10474;
    wire [7:0] _667;
    reg [7:0] _3477;
    wire _10481;
    wire _10478;
    wire _10479;
    wire _10482;
    wire [7:0] _10483;
    wire _10476;
    wire _10477;
    wire [7:0] _10485;
    wire [7:0] _10487;
    wire [7:0] _668;
    reg [7:0] _3474;
    wire _10494;
    wire _10491;
    wire _10492;
    wire _10495;
    wire [7:0] _10496;
    wire _10489;
    wire _10490;
    wire [7:0] _10498;
    wire [7:0] _10500;
    wire [7:0] _669;
    reg [7:0] _3471;
    wire _10507;
    wire _10504;
    wire _10505;
    wire _10508;
    wire [7:0] _10509;
    wire _10502;
    wire _10503;
    wire [7:0] _10511;
    wire [7:0] _10513;
    wire [7:0] _670;
    reg [7:0] _3468;
    wire _10520;
    wire _10517;
    wire _10518;
    wire _10521;
    wire [7:0] _10522;
    wire _10515;
    wire _10516;
    wire [7:0] _10524;
    wire [7:0] _10526;
    wire [7:0] _671;
    reg [7:0] _3465;
    wire _10533;
    wire _10530;
    wire _10531;
    wire _10534;
    wire [7:0] _10535;
    wire _10528;
    wire _10529;
    wire [7:0] _10537;
    wire [7:0] _10539;
    wire [7:0] _672;
    reg [7:0] _3462;
    wire _10546;
    wire _10543;
    wire _10544;
    wire _10547;
    wire [7:0] _10548;
    wire _10541;
    wire _10542;
    wire [7:0] _10550;
    wire [7:0] _10552;
    wire [7:0] _673;
    reg [7:0] _3459;
    wire _10559;
    wire _10556;
    wire _10557;
    wire _10560;
    wire [7:0] _10561;
    wire _10554;
    wire _10555;
    wire [7:0] _10563;
    wire [7:0] _10565;
    wire [7:0] _674;
    reg [7:0] _3456;
    wire _10572;
    wire _10569;
    wire _10570;
    wire _10573;
    wire [7:0] _10574;
    wire _10567;
    wire _10568;
    wire [7:0] _10576;
    wire [7:0] _10578;
    wire [7:0] _675;
    reg [7:0] _3453;
    wire _10585;
    wire _10582;
    wire _10583;
    wire _10586;
    wire [7:0] _10587;
    wire _10580;
    wire _10581;
    wire [7:0] _10589;
    wire [7:0] _10591;
    wire [7:0] _676;
    reg [7:0] _3450;
    wire _10598;
    wire _10595;
    wire _10596;
    wire _10599;
    wire [7:0] _10600;
    wire _10593;
    wire _10594;
    wire [7:0] _10602;
    wire [7:0] _10604;
    wire [7:0] _677;
    reg [7:0] _3447;
    wire _10611;
    wire _10608;
    wire _10609;
    wire _10612;
    wire [7:0] _10613;
    wire _10606;
    wire _10607;
    wire [7:0] _10615;
    wire [7:0] _10617;
    wire [7:0] _678;
    reg [7:0] _3444;
    wire _10624;
    wire _10621;
    wire _10622;
    wire _10625;
    wire [7:0] _10626;
    wire _10619;
    wire _10620;
    wire [7:0] _10628;
    wire [7:0] _10630;
    wire [7:0] _679;
    reg [7:0] _3441;
    wire _10637;
    wire _10634;
    wire _10635;
    wire _10638;
    wire [7:0] _10639;
    wire _10632;
    wire _10633;
    wire [7:0] _10641;
    wire [7:0] _10643;
    wire [7:0] _680;
    reg [7:0] _3438;
    wire _10650;
    wire _10647;
    wire _10648;
    wire _10651;
    wire [7:0] _10652;
    wire _10645;
    wire _10646;
    wire [7:0] _10654;
    wire [7:0] _10656;
    wire [7:0] _681;
    reg [7:0] _3435;
    wire _10663;
    wire _10660;
    wire _10661;
    wire _10664;
    wire [7:0] _10665;
    wire _10658;
    wire _10659;
    wire [7:0] _10667;
    wire [7:0] _10669;
    wire [7:0] _682;
    reg [7:0] _3432;
    wire _10676;
    wire _10673;
    wire _10674;
    wire _10677;
    wire [7:0] _10678;
    wire _10671;
    wire _10672;
    wire [7:0] _10680;
    wire [7:0] _10682;
    wire [7:0] _683;
    reg [7:0] _3429;
    wire _10689;
    wire _10686;
    wire _10687;
    wire _10690;
    wire [7:0] _10691;
    wire _10684;
    wire _10685;
    wire [7:0] _10693;
    wire [7:0] _10695;
    wire [7:0] _684;
    reg [7:0] _3426;
    wire _10702;
    wire _10699;
    wire _10700;
    wire _10703;
    wire [7:0] _10704;
    wire _10697;
    wire _10698;
    wire [7:0] _10706;
    wire [7:0] _10708;
    wire [7:0] _685;
    reg [7:0] _3423;
    wire _10715;
    wire _10712;
    wire _10713;
    wire _10716;
    wire [7:0] _10717;
    wire _10710;
    wire _10711;
    wire [7:0] _10719;
    wire [7:0] _10721;
    wire [7:0] _686;
    reg [7:0] _3420;
    wire _10728;
    wire _10725;
    wire _10726;
    wire _10729;
    wire [7:0] _10730;
    wire _10723;
    wire _10724;
    wire [7:0] _10732;
    wire [7:0] _10734;
    wire [7:0] _687;
    reg [7:0] _3417;
    wire _10741;
    wire _10738;
    wire _10739;
    wire _10742;
    wire [7:0] _10743;
    wire _10736;
    wire _10737;
    wire [7:0] _10745;
    wire [7:0] _10747;
    wire [7:0] _688;
    reg [7:0] _3414;
    wire _10754;
    wire _10751;
    wire _10752;
    wire _10755;
    wire [7:0] _10756;
    wire _10749;
    wire _10750;
    wire [7:0] _10758;
    wire [7:0] _10760;
    wire [7:0] _689;
    reg [7:0] _3411;
    wire _10767;
    wire _10764;
    wire _10765;
    wire _10768;
    wire [7:0] _10769;
    wire _10762;
    wire _10763;
    wire [7:0] _10771;
    wire [7:0] _10773;
    wire [7:0] _690;
    reg [7:0] _3408;
    wire _10780;
    wire _10777;
    wire _10778;
    wire _10781;
    wire [7:0] _10782;
    wire _10775;
    wire _10776;
    wire [7:0] _10784;
    wire [7:0] _10786;
    wire [7:0] _691;
    reg [7:0] _3405;
    wire _10793;
    wire _10790;
    wire _10791;
    wire _10794;
    wire [7:0] _10795;
    wire _10788;
    wire _10789;
    wire [7:0] _10797;
    wire [7:0] _10799;
    wire [7:0] _692;
    reg [7:0] _3402;
    wire _10806;
    wire _10803;
    wire _10804;
    wire _10807;
    wire [7:0] _10808;
    wire _10801;
    wire _10802;
    wire [7:0] _10810;
    wire [7:0] _10812;
    wire [7:0] _693;
    reg [7:0] _3399;
    wire _10819;
    wire _10816;
    wire _10817;
    wire _10820;
    wire [7:0] _10821;
    wire _10814;
    wire _10815;
    wire [7:0] _10823;
    wire [7:0] _10825;
    wire [7:0] _694;
    reg [7:0] _3396;
    wire _10832;
    wire _10829;
    wire _10830;
    wire _10833;
    wire [7:0] _10834;
    wire _10827;
    wire _10828;
    wire [7:0] _10836;
    wire [7:0] _10838;
    wire [7:0] _695;
    reg [7:0] _3393;
    wire _10845;
    wire _10842;
    wire _10843;
    wire _10846;
    wire [7:0] _10847;
    wire _10840;
    wire _10841;
    wire [7:0] _10849;
    wire [7:0] _10851;
    wire [7:0] _696;
    reg [7:0] _3390;
    wire _10858;
    wire _10855;
    wire _10856;
    wire _10859;
    wire [7:0] _10860;
    wire _10853;
    wire _10854;
    wire [7:0] _10862;
    wire [7:0] _10864;
    wire [7:0] _697;
    reg [7:0] _3387;
    wire _10871;
    wire _10868;
    wire _10869;
    wire _10872;
    wire [7:0] _10873;
    wire _10866;
    wire _10867;
    wire [7:0] _10875;
    wire [7:0] _10877;
    wire [7:0] _698;
    reg [7:0] _3384;
    wire _10884;
    wire _10881;
    wire _10882;
    wire _10885;
    wire [7:0] _10886;
    wire _10879;
    wire _10880;
    wire [7:0] _10888;
    wire [7:0] _10890;
    wire [7:0] _699;
    reg [7:0] _3381;
    wire _10897;
    wire _10894;
    wire _10895;
    wire _10898;
    wire [7:0] _10899;
    wire _10892;
    wire _10893;
    wire [7:0] _10901;
    wire [7:0] _10903;
    wire [7:0] _700;
    reg [7:0] _3378;
    wire _10910;
    wire _10907;
    wire _10908;
    wire _10911;
    wire [7:0] _10912;
    wire _10905;
    wire _10906;
    wire [7:0] _10914;
    wire [7:0] _10916;
    wire [7:0] _701;
    reg [7:0] _3375;
    wire _10923;
    wire _10920;
    wire _10921;
    wire _10924;
    wire [7:0] _10925;
    wire _10918;
    wire _10919;
    wire [7:0] _10927;
    wire [7:0] _10929;
    wire [7:0] _702;
    reg [7:0] _3372;
    wire _10936;
    wire _10933;
    wire _10934;
    wire _10937;
    wire [7:0] _10938;
    wire _10931;
    wire _10932;
    wire [7:0] _10940;
    wire [7:0] _10942;
    wire [7:0] _703;
    reg [7:0] _3369;
    wire _10949;
    wire _10946;
    wire _10947;
    wire _10950;
    wire [7:0] _10951;
    wire _10944;
    wire _10945;
    wire [7:0] _10953;
    wire [7:0] _10955;
    wire [7:0] _704;
    reg [7:0] _3366;
    wire _10962;
    wire _10959;
    wire _10960;
    wire _10963;
    wire [7:0] _10964;
    wire _10957;
    wire _10958;
    wire [7:0] _10966;
    wire [7:0] _10968;
    wire [7:0] _705;
    reg [7:0] _3363;
    wire _10975;
    wire _10972;
    wire _10973;
    wire _10976;
    wire [7:0] _10977;
    wire _10970;
    wire _10971;
    wire [7:0] _10979;
    wire [7:0] _10981;
    wire [7:0] _706;
    reg [7:0] _3360;
    wire _10988;
    wire _10985;
    wire _10986;
    wire _10989;
    wire [7:0] _10990;
    wire _10983;
    wire _10984;
    wire [7:0] _10992;
    wire [7:0] _10994;
    wire [7:0] _707;
    reg [7:0] _3357;
    wire _11001;
    wire _10998;
    wire _10999;
    wire _11002;
    wire [7:0] _11003;
    wire _10996;
    wire _10997;
    wire [7:0] _11005;
    wire [7:0] _11007;
    wire [7:0] _708;
    reg [7:0] _3354;
    wire _11014;
    wire _11011;
    wire _11012;
    wire _11015;
    wire [7:0] _11016;
    wire _11009;
    wire _11010;
    wire [7:0] _11018;
    wire [7:0] _11020;
    wire [7:0] _709;
    reg [7:0] _3351;
    wire _11027;
    wire _11024;
    wire _11025;
    wire _11028;
    wire [7:0] _11029;
    wire _11022;
    wire _11023;
    wire [7:0] _11031;
    wire [7:0] _11033;
    wire [7:0] _710;
    reg [7:0] _3348;
    wire _11040;
    wire _11037;
    wire _11038;
    wire _11041;
    wire [7:0] _11042;
    wire _11035;
    wire _11036;
    wire [7:0] _11044;
    wire [7:0] _11046;
    wire [7:0] _711;
    reg [7:0] _3345;
    wire _11053;
    wire _11050;
    wire _11051;
    wire _11054;
    wire [7:0] _11055;
    wire _11048;
    wire _11049;
    wire [7:0] _11057;
    wire [7:0] _11059;
    wire [7:0] _712;
    reg [7:0] _3342;
    wire _11066;
    wire _11063;
    wire _11064;
    wire _11067;
    wire [7:0] _11068;
    wire _11061;
    wire _11062;
    wire [7:0] _11070;
    wire [7:0] _11072;
    wire [7:0] _713;
    reg [7:0] _3339;
    wire _11079;
    wire _11076;
    wire _11077;
    wire _11080;
    wire [7:0] _11081;
    wire _11074;
    wire _11075;
    wire [7:0] _11083;
    wire [7:0] _11085;
    wire [7:0] _714;
    reg [7:0] _3336;
    wire _11092;
    wire _11089;
    wire _11090;
    wire _11093;
    wire [7:0] _11094;
    wire _11087;
    wire _11088;
    wire [7:0] _11096;
    wire [7:0] _11098;
    wire [7:0] _715;
    reg [7:0] _3333;
    wire _11105;
    wire _11102;
    wire _11103;
    wire _11106;
    wire [7:0] _11107;
    wire _11100;
    wire _11101;
    wire [7:0] _11109;
    wire [7:0] _11111;
    wire [7:0] _716;
    reg [7:0] _3330;
    wire _11118;
    wire _11115;
    wire _11116;
    wire _11119;
    wire [7:0] _11120;
    wire _11113;
    wire _11114;
    wire [7:0] _11122;
    wire [7:0] _11124;
    wire [7:0] _717;
    reg [7:0] _3327;
    wire _11131;
    wire _11128;
    wire _11129;
    wire _11132;
    wire [7:0] _11133;
    wire _11126;
    wire _11127;
    wire [7:0] _11135;
    wire [7:0] _11137;
    wire [7:0] _718;
    reg [7:0] _3324;
    wire _11144;
    wire _11141;
    wire _11142;
    wire _11145;
    wire [7:0] _11146;
    wire _11139;
    wire _11140;
    wire [7:0] _11148;
    wire [7:0] _11150;
    wire [7:0] _719;
    reg [7:0] _3321;
    wire _11157;
    wire _11154;
    wire _11155;
    wire _11158;
    wire [7:0] _11159;
    wire _11152;
    wire _11153;
    wire [7:0] _11161;
    wire [7:0] _11163;
    wire [7:0] _720;
    reg [7:0] _3318;
    wire _11170;
    wire _11167;
    wire _11168;
    wire _11171;
    wire [7:0] _11172;
    wire _11165;
    wire _11166;
    wire [7:0] _11174;
    wire [7:0] _11176;
    wire [7:0] _721;
    reg [7:0] _3315;
    wire _11183;
    wire _11180;
    wire _11181;
    wire _11184;
    wire [7:0] _11185;
    wire _11178;
    wire _11179;
    wire [7:0] _11187;
    wire [7:0] _11189;
    wire [7:0] _722;
    reg [7:0] _3312;
    wire _11196;
    wire _11193;
    wire _11194;
    wire _11197;
    wire [7:0] _11198;
    wire _11191;
    wire _11192;
    wire [7:0] _11200;
    wire [7:0] _11202;
    wire [7:0] _723;
    reg [7:0] _3309;
    wire _11209;
    wire _11206;
    wire _11207;
    wire _11210;
    wire [7:0] _11211;
    wire _11204;
    wire _11205;
    wire [7:0] _11213;
    wire [7:0] _11215;
    wire [7:0] _724;
    reg [7:0] _3306;
    wire _11222;
    wire _11219;
    wire _11220;
    wire _11223;
    wire [7:0] _11224;
    wire _11217;
    wire _11218;
    wire [7:0] _11226;
    wire [7:0] _11228;
    wire [7:0] _725;
    reg [7:0] _3303;
    wire _11235;
    wire _11232;
    wire _11233;
    wire _11236;
    wire [7:0] _11237;
    wire _11230;
    wire _11231;
    wire [7:0] _11239;
    wire [7:0] _11241;
    wire [7:0] _726;
    reg [7:0] _3300;
    wire _11248;
    wire _11245;
    wire _11246;
    wire _11249;
    wire [7:0] _11250;
    wire _11243;
    wire _11244;
    wire [7:0] _11252;
    wire [7:0] _11254;
    wire [7:0] _727;
    reg [7:0] _3297;
    wire _11261;
    wire _11258;
    wire _11259;
    wire _11262;
    wire [7:0] _11263;
    wire _11256;
    wire _11257;
    wire [7:0] _11265;
    wire [7:0] _11267;
    wire [7:0] _728;
    reg [7:0] _3294;
    wire _11274;
    wire _11271;
    wire _11272;
    wire _11275;
    wire [7:0] _11276;
    wire _11269;
    wire _11270;
    wire [7:0] _11278;
    wire [7:0] _11280;
    wire [7:0] _729;
    reg [7:0] _3291;
    wire _11287;
    wire _11284;
    wire _11285;
    wire _11288;
    wire [7:0] _11289;
    wire _11282;
    wire _11283;
    wire [7:0] _11291;
    wire [7:0] _11293;
    wire [7:0] _730;
    reg [7:0] _3288;
    wire _11300;
    wire _11297;
    wire _11298;
    wire _11301;
    wire [7:0] _11302;
    wire _11295;
    wire _11296;
    wire [7:0] _11304;
    wire [7:0] _11306;
    wire [7:0] _731;
    reg [7:0] _3285;
    wire _11313;
    wire _11310;
    wire _11311;
    wire _11314;
    wire [7:0] _11315;
    wire _11308;
    wire _11309;
    wire [7:0] _11317;
    wire [7:0] _11319;
    wire [7:0] _732;
    reg [7:0] _3282;
    wire _11326;
    wire _11323;
    wire _11324;
    wire _11327;
    wire [7:0] _11328;
    wire _11321;
    wire _11322;
    wire [7:0] _11330;
    wire [7:0] _11332;
    wire [7:0] _733;
    reg [7:0] _3279;
    wire _11339;
    wire _11336;
    wire _11337;
    wire _11340;
    wire [7:0] _11341;
    wire _11334;
    wire _11335;
    wire [7:0] _11343;
    wire [7:0] _11345;
    wire [7:0] _734;
    reg [7:0] _3276;
    wire _11352;
    wire _11349;
    wire _11350;
    wire _11353;
    wire [7:0] _11354;
    wire _11347;
    wire _11348;
    wire [7:0] _11356;
    wire [7:0] _11358;
    wire [7:0] _735;
    reg [7:0] _3273;
    wire _11365;
    wire _11362;
    wire _11363;
    wire _11366;
    wire [7:0] _11367;
    wire _11360;
    wire _11361;
    wire [7:0] _11369;
    wire [7:0] _11371;
    wire [7:0] _736;
    reg [7:0] _3270;
    wire _11378;
    wire _11375;
    wire _11376;
    wire _11379;
    wire [7:0] _11380;
    wire _11373;
    wire _11374;
    wire [7:0] _11382;
    wire [7:0] _11384;
    wire [7:0] _737;
    reg [7:0] _3267;
    wire _11391;
    wire _11388;
    wire _11389;
    wire _11392;
    wire [7:0] _11393;
    wire _11386;
    wire _11387;
    wire [7:0] _11395;
    wire [7:0] _11397;
    wire [7:0] _738;
    reg [7:0] _3264;
    wire _11404;
    wire _11401;
    wire _11402;
    wire _11405;
    wire [7:0] _11406;
    wire _11399;
    wire _11400;
    wire [7:0] _11408;
    wire [7:0] _11410;
    wire [7:0] _739;
    reg [7:0] _3261;
    wire _11417;
    wire _11414;
    wire _11415;
    wire _11418;
    wire [7:0] _11419;
    wire _11412;
    wire _11413;
    wire [7:0] _11421;
    wire [7:0] _11423;
    wire [7:0] _740;
    reg [7:0] _3258;
    wire _11430;
    wire _11427;
    wire _11428;
    wire _11431;
    wire [7:0] _11432;
    wire _11425;
    wire _11426;
    wire [7:0] _11434;
    wire [7:0] _11436;
    wire [7:0] _741;
    reg [7:0] _3255;
    wire _11443;
    wire _11440;
    wire _11441;
    wire _11444;
    wire [7:0] _11445;
    wire _11438;
    wire _11439;
    wire [7:0] _11447;
    wire [7:0] _11449;
    wire [7:0] _742;
    reg [7:0] _3252;
    wire _11456;
    wire _11453;
    wire _11454;
    wire _11457;
    wire [7:0] _11458;
    wire _11451;
    wire _11452;
    wire [7:0] _11460;
    wire [7:0] _11462;
    wire [7:0] _743;
    reg [7:0] _3249;
    wire _11469;
    wire _11466;
    wire _11467;
    wire _11470;
    wire [7:0] _11471;
    wire _11464;
    wire _11465;
    wire [7:0] _11473;
    wire [7:0] _11475;
    wire [7:0] _744;
    reg [7:0] _3246;
    wire _11482;
    wire _11479;
    wire _11480;
    wire _11483;
    wire [7:0] _11484;
    wire _11477;
    wire _11478;
    wire [7:0] _11486;
    wire [7:0] _11488;
    wire [7:0] _745;
    reg [7:0] _3243;
    wire _11495;
    wire _11492;
    wire _11493;
    wire _11496;
    wire [7:0] _11497;
    wire _11490;
    wire _11491;
    wire [7:0] _11499;
    wire [7:0] _11501;
    wire [7:0] _746;
    reg [7:0] _3240;
    wire _11508;
    wire _11505;
    wire _11506;
    wire _11509;
    wire [7:0] _11510;
    wire _11503;
    wire _11504;
    wire [7:0] _11512;
    wire [7:0] _11514;
    wire [7:0] _747;
    reg [7:0] _3237;
    wire _11521;
    wire _11518;
    wire _11519;
    wire _11522;
    wire [7:0] _11523;
    wire _11516;
    wire _11517;
    wire [7:0] _11525;
    wire [7:0] _11527;
    wire [7:0] _748;
    reg [7:0] _3234;
    wire _11534;
    wire _11531;
    wire _11532;
    wire _11535;
    wire [7:0] _11536;
    wire _11529;
    wire _11530;
    wire [7:0] _11538;
    wire [7:0] _11540;
    wire [7:0] _749;
    reg [7:0] _3231;
    wire _11547;
    wire _11544;
    wire _11545;
    wire _11548;
    wire [7:0] _11549;
    wire _11542;
    wire _11543;
    wire [7:0] _11551;
    wire [7:0] _11553;
    wire [7:0] _750;
    reg [7:0] _3228;
    wire _11560;
    wire _11557;
    wire _11558;
    wire _11561;
    wire [7:0] _11562;
    wire _11555;
    wire _11556;
    wire [7:0] _11564;
    wire [7:0] _11566;
    wire [7:0] _751;
    reg [7:0] _3225;
    wire _11573;
    wire _11570;
    wire _11571;
    wire _11574;
    wire [7:0] _11575;
    wire _11568;
    wire _11569;
    wire [7:0] _11577;
    wire [7:0] _11579;
    wire [7:0] _752;
    reg [7:0] _3222;
    wire _11586;
    wire _11583;
    wire _11584;
    wire _11587;
    wire [7:0] _11588;
    wire _11581;
    wire _11582;
    wire [7:0] _11590;
    wire [7:0] _11592;
    wire [7:0] _753;
    reg [7:0] _3219;
    wire _11599;
    wire _11596;
    wire _11597;
    wire _11600;
    wire [7:0] _11601;
    wire _11594;
    wire _11595;
    wire [7:0] _11603;
    wire [7:0] _11605;
    wire [7:0] _754;
    reg [7:0] _3216;
    wire _11612;
    wire _11609;
    wire _11610;
    wire _11613;
    wire [7:0] _11614;
    wire _11607;
    wire _11608;
    wire [7:0] _11616;
    wire [7:0] _11618;
    wire [7:0] _755;
    reg [7:0] _3213;
    wire _11625;
    wire _11622;
    wire _11623;
    wire _11626;
    wire [7:0] _11627;
    wire _11620;
    wire _11621;
    wire [7:0] _11629;
    wire [7:0] _11631;
    wire [7:0] _756;
    reg [7:0] _3210;
    wire _11638;
    wire _11635;
    wire _11636;
    wire _11639;
    wire [7:0] _11640;
    wire _11633;
    wire _11634;
    wire [7:0] _11642;
    wire [7:0] _11644;
    wire [7:0] _757;
    reg [7:0] _3207;
    wire _11651;
    wire _11648;
    wire _11649;
    wire _11652;
    wire [7:0] _11653;
    wire _11646;
    wire _11647;
    wire [7:0] _11655;
    wire [7:0] _11657;
    wire [7:0] _758;
    reg [7:0] _3204;
    wire _11664;
    wire _11661;
    wire _11662;
    wire _11665;
    wire [7:0] _11666;
    wire _11659;
    wire _11660;
    wire [7:0] _11668;
    wire [7:0] _11670;
    wire [7:0] _759;
    reg [7:0] _3201;
    wire _11677;
    wire _11674;
    wire _11675;
    wire _11678;
    wire [7:0] _11679;
    wire _11672;
    wire _11673;
    wire [7:0] _11681;
    wire [7:0] _11683;
    wire [7:0] _760;
    reg [7:0] _3198;
    wire _11690;
    wire _11687;
    wire _11688;
    wire _11691;
    wire [7:0] _11692;
    wire _11685;
    wire _11686;
    wire [7:0] _11694;
    wire [7:0] _11696;
    wire [7:0] _761;
    reg [7:0] _3195;
    wire _11703;
    wire _11700;
    wire _11701;
    wire _11704;
    wire [7:0] _11705;
    wire _11698;
    wire _11699;
    wire [7:0] _11707;
    wire [7:0] _11709;
    wire [7:0] _762;
    reg [7:0] _3192;
    wire _11716;
    wire _11713;
    wire _11714;
    wire _11717;
    wire [7:0] _11718;
    wire _11711;
    wire _11712;
    wire [7:0] _11720;
    wire [7:0] _11722;
    wire [7:0] _763;
    reg [7:0] _3189;
    wire _11729;
    wire _11726;
    wire _11727;
    wire _11730;
    wire [7:0] _11731;
    wire _11724;
    wire _11725;
    wire [7:0] _11733;
    wire [7:0] _11735;
    wire [7:0] _764;
    reg [7:0] _3186;
    wire _11742;
    wire _11739;
    wire _11740;
    wire _11743;
    wire [7:0] _11744;
    wire _11737;
    wire _11738;
    wire [7:0] _11746;
    wire [7:0] _11748;
    wire [7:0] _765;
    reg [7:0] _3183;
    wire _11755;
    wire _11752;
    wire _11753;
    wire _11756;
    wire [7:0] _11757;
    wire _11750;
    wire _11751;
    wire [7:0] _11759;
    wire [7:0] _11761;
    wire [7:0] _766;
    reg [7:0] _3180;
    wire _11768;
    wire _11765;
    wire _11766;
    wire _11769;
    wire [7:0] _11770;
    wire _11763;
    wire _11764;
    wire [7:0] _11772;
    wire [7:0] _11774;
    wire [7:0] _767;
    reg [7:0] _3177;
    wire _11781;
    wire _11778;
    wire _11779;
    wire _11782;
    wire [7:0] _11783;
    wire _11776;
    wire _11777;
    wire [7:0] _11785;
    wire [7:0] _11787;
    wire [7:0] _768;
    reg [7:0] _3174;
    wire _11794;
    wire _11791;
    wire _11792;
    wire _11795;
    wire [7:0] _11796;
    wire _11789;
    wire _11790;
    wire [7:0] _11798;
    wire [7:0] _11800;
    wire [7:0] _769;
    reg [7:0] _3171;
    wire _11807;
    wire _11804;
    wire _11805;
    wire _11808;
    wire [7:0] _11809;
    wire _11802;
    wire _11803;
    wire [7:0] _11811;
    wire [7:0] _11813;
    wire [7:0] _770;
    reg [7:0] _3168;
    wire _11820;
    wire _11817;
    wire _11818;
    wire _11821;
    wire [7:0] _11822;
    wire _11815;
    wire _11816;
    wire [7:0] _11824;
    wire [7:0] _11826;
    wire [7:0] _771;
    reg [7:0] _3165;
    wire _11833;
    wire _11830;
    wire _11831;
    wire _11834;
    wire [7:0] _11835;
    wire _11828;
    wire _11829;
    wire [7:0] _11837;
    wire [7:0] _11839;
    wire [7:0] _772;
    reg [7:0] _3162;
    wire _11846;
    wire _11843;
    wire _11844;
    wire _11847;
    wire [7:0] _11848;
    wire _11841;
    wire _11842;
    wire [7:0] _11850;
    wire [7:0] _11852;
    wire [7:0] _773;
    reg [7:0] _3159;
    wire _11859;
    wire _11856;
    wire _11857;
    wire _11860;
    wire [7:0] _11861;
    wire _11854;
    wire _11855;
    wire [7:0] _11863;
    wire [7:0] _11865;
    wire [7:0] _774;
    reg [7:0] _3156;
    wire _11872;
    wire _11869;
    wire _11870;
    wire _11873;
    wire [7:0] _11874;
    wire _11867;
    wire _11868;
    wire [7:0] _11876;
    wire [7:0] _11878;
    wire [7:0] _775;
    reg [7:0] _3153;
    wire _11885;
    wire _11882;
    wire _11883;
    wire _11886;
    wire [7:0] _11887;
    wire _11880;
    wire _11881;
    wire [7:0] _11889;
    wire [7:0] _11891;
    wire [7:0] _776;
    reg [7:0] _3150;
    wire _11898;
    wire _11895;
    wire _11896;
    wire _11899;
    wire [7:0] _11900;
    wire _11893;
    wire _11894;
    wire [7:0] _11902;
    wire [7:0] _11904;
    wire [7:0] _777;
    reg [7:0] _3147;
    wire _11911;
    wire _11908;
    wire _11909;
    wire _11912;
    wire [7:0] _11913;
    wire _11906;
    wire _11907;
    wire [7:0] _11915;
    wire [7:0] _11917;
    wire [7:0] _778;
    reg [7:0] _3144;
    wire _11924;
    wire _11921;
    wire _11922;
    wire _11925;
    wire [7:0] _11926;
    wire _11919;
    wire _11920;
    wire [7:0] _11928;
    wire [7:0] _11930;
    wire [7:0] _779;
    reg [7:0] _3141;
    wire [7:0] _781;
    reg [7:0] _3912;
    reg [7:0] _3913;
    reg [7:0] _3914;
    reg [7:0] _3915;
    reg [7:0] _3916;
    reg [7:0] _3917;
    reg [7:0] _3918;
    reg [7:0] _3919;
    wire [7:0] _5304;
    wire _11937;
    wire _11934;
    wire _11935;
    wire _11938;
    wire [15:0] _11939;
    wire _11932;
    wire _11933;
    wire [15:0] _11941;
    wire [15:0] _11943;
    wire [15:0] _782;
    reg [15:0] _3925;
    reg [15:0] _4691;
    wire _5302;
    wire _5303;
    wire [7:0] _8620;
    wire _11950;
    wire _11947;
    wire _11948;
    wire _11951;
    wire [7:0] _11952;
    wire _11945;
    wire _11946;
    wire [7:0] _11954;
    wire [7:0] _11956;
    wire [7:0] _783;
    reg [7:0] _3138;
    wire [7:0] _785;
    reg [7:0] _3904;
    reg [7:0] _3905;
    reg [7:0] _3906;
    reg [7:0] _3907;
    reg [7:0] _3908;
    reg [7:0] _3909;
    reg [7:0] _3910;
    reg [7:0] _3911;
    wire _3920;
    wire _3921;
    wire _3922;
    wire _4698;
    wire _11989;
    wire [2:0] _11993;
    wire _11988;
    wire [2:0] _11994;
    wire _11986;
    wire _11987;
    wire [2:0] _11995;
    wire _11984;
    wire _11985;
    wire [2:0] _11996;
    wire [7:0] _11978;
    wire [7:0] _11972;
    wire _11968;
    wire _11969;
    wire _11970;
    wire [7:0] _11974;
    wire [7:0] _787;
    wire vdd;
    wire _789;
    wire _791;
    wire [7:0] _11962;
    wire [7:0] _11958;
    wire _793;
    wire _795;
    wire [2:0] _3131;
    wire _3132;
    wire _3133;
    wire _797;
    wire _3129;
    wire _3130;
    wire _3134;
    wire _3135;
    wire [2:0] _3127;
    wire _3128;
    wire _4715;
    wire _4716;
    wire [7:0] _11960;
    wire [7:0] _11963;
    wire [7:0] _798;
    reg [7:0] _4729;
    wire _5269;
    wire [2:0] _4713;
    wire _4714;
    wire _5270;
    wire [7:0] _11976;
    wire _11966;
    wire _11967;
    wire [7:0] _11979;
    wire [7:0] _799;
    reg [7:0] _5296;
    wire _11964;
    wire [2:0] _5291;
    wire _5292;
    wire _5293;
    wire _11965;
    wire [2:0] _5289;
    wire _5290;
    wire _11983;
    wire [2:0] _11997;
    wire _801;
    wire _803;
    wire _814;
    wire _11980;
    wire _11981;
    wire _11982;
    wire [2:0] _11998;
    wire _805;
    wire [2:0] _11999;
    wire [2:0] _806;
    reg [2:0] _811;
    wire _813;
    assign _4700 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    always @* begin
        case (_781)
        0:
            _4708 <= _3123;
        1:
            _4708 <= _3109;
        2:
            _4708 <= _3100;
        3:
            _4708 <= _3091;
        4:
            _4708 <= _3082;
        5:
            _4708 <= _3073;
        6:
            _4708 <= _3064;
        7:
            _4708 <= _3055;
        8:
            _4708 <= _3046;
        9:
            _4708 <= _3037;
        10:
            _4708 <= _3028;
        11:
            _4708 <= _3019;
        12:
            _4708 <= _3010;
        13:
            _4708 <= _3001;
        14:
            _4708 <= _2992;
        15:
            _4708 <= _2983;
        16:
            _4708 <= _2974;
        17:
            _4708 <= _2965;
        18:
            _4708 <= _2956;
        19:
            _4708 <= _2947;
        20:
            _4708 <= _2938;
        21:
            _4708 <= _2929;
        22:
            _4708 <= _2920;
        23:
            _4708 <= _2911;
        24:
            _4708 <= _2902;
        25:
            _4708 <= _2893;
        26:
            _4708 <= _2884;
        27:
            _4708 <= _2875;
        28:
            _4708 <= _2866;
        29:
            _4708 <= _2857;
        30:
            _4708 <= _2848;
        31:
            _4708 <= _2839;
        32:
            _4708 <= _2830;
        33:
            _4708 <= _2821;
        34:
            _4708 <= _2812;
        35:
            _4708 <= _2803;
        36:
            _4708 <= _2794;
        37:
            _4708 <= _2785;
        38:
            _4708 <= _2776;
        39:
            _4708 <= _2767;
        40:
            _4708 <= _2758;
        41:
            _4708 <= _2749;
        42:
            _4708 <= _2740;
        43:
            _4708 <= _2731;
        44:
            _4708 <= _2722;
        45:
            _4708 <= _2713;
        46:
            _4708 <= _2704;
        47:
            _4708 <= _2695;
        48:
            _4708 <= _2686;
        49:
            _4708 <= _2677;
        50:
            _4708 <= _2668;
        51:
            _4708 <= _2659;
        52:
            _4708 <= _2650;
        53:
            _4708 <= _2641;
        54:
            _4708 <= _2632;
        55:
            _4708 <= _2623;
        56:
            _4708 <= _2614;
        57:
            _4708 <= _2605;
        58:
            _4708 <= _2596;
        59:
            _4708 <= _2587;
        60:
            _4708 <= _2578;
        61:
            _4708 <= _2569;
        62:
            _4708 <= _2560;
        63:
            _4708 <= _2551;
        64:
            _4708 <= _2542;
        65:
            _4708 <= _2533;
        66:
            _4708 <= _2524;
        67:
            _4708 <= _2515;
        68:
            _4708 <= _2506;
        69:
            _4708 <= _2497;
        70:
            _4708 <= _2488;
        71:
            _4708 <= _2479;
        72:
            _4708 <= _2470;
        73:
            _4708 <= _2461;
        74:
            _4708 <= _2452;
        75:
            _4708 <= _2443;
        76:
            _4708 <= _2434;
        77:
            _4708 <= _2425;
        78:
            _4708 <= _2416;
        79:
            _4708 <= _2407;
        80:
            _4708 <= _2398;
        81:
            _4708 <= _2389;
        82:
            _4708 <= _2380;
        83:
            _4708 <= _2371;
        84:
            _4708 <= _2362;
        85:
            _4708 <= _2353;
        86:
            _4708 <= _2344;
        87:
            _4708 <= _2335;
        88:
            _4708 <= _2326;
        89:
            _4708 <= _2317;
        90:
            _4708 <= _2308;
        91:
            _4708 <= _2299;
        92:
            _4708 <= _2290;
        93:
            _4708 <= _2281;
        94:
            _4708 <= _2272;
        95:
            _4708 <= _2263;
        96:
            _4708 <= _2254;
        97:
            _4708 <= _2245;
        98:
            _4708 <= _2236;
        99:
            _4708 <= _2227;
        100:
            _4708 <= _2218;
        101:
            _4708 <= _2209;
        102:
            _4708 <= _2200;
        103:
            _4708 <= _2191;
        104:
            _4708 <= _2182;
        105:
            _4708 <= _2173;
        106:
            _4708 <= _2164;
        107:
            _4708 <= _2155;
        108:
            _4708 <= _2146;
        109:
            _4708 <= _2137;
        110:
            _4708 <= _2128;
        111:
            _4708 <= _2119;
        112:
            _4708 <= _2110;
        113:
            _4708 <= _2101;
        114:
            _4708 <= _2092;
        115:
            _4708 <= _2083;
        116:
            _4708 <= _2074;
        117:
            _4708 <= _2065;
        118:
            _4708 <= _2056;
        119:
            _4708 <= _2047;
        120:
            _4708 <= _2038;
        121:
            _4708 <= _2029;
        122:
            _4708 <= _2020;
        123:
            _4708 <= _2011;
        124:
            _4708 <= _2002;
        125:
            _4708 <= _1993;
        126:
            _4708 <= _1984;
        127:
            _4708 <= _1975;
        128:
            _4708 <= _1966;
        129:
            _4708 <= _1957;
        130:
            _4708 <= _1948;
        131:
            _4708 <= _1939;
        132:
            _4708 <= _1930;
        133:
            _4708 <= _1921;
        134:
            _4708 <= _1912;
        135:
            _4708 <= _1903;
        136:
            _4708 <= _1894;
        137:
            _4708 <= _1885;
        138:
            _4708 <= _1876;
        139:
            _4708 <= _1867;
        140:
            _4708 <= _1858;
        141:
            _4708 <= _1849;
        142:
            _4708 <= _1840;
        143:
            _4708 <= _1831;
        144:
            _4708 <= _1822;
        145:
            _4708 <= _1813;
        146:
            _4708 <= _1804;
        147:
            _4708 <= _1795;
        148:
            _4708 <= _1786;
        149:
            _4708 <= _1777;
        150:
            _4708 <= _1768;
        151:
            _4708 <= _1759;
        152:
            _4708 <= _1750;
        153:
            _4708 <= _1741;
        154:
            _4708 <= _1732;
        155:
            _4708 <= _1723;
        156:
            _4708 <= _1714;
        157:
            _4708 <= _1705;
        158:
            _4708 <= _1696;
        159:
            _4708 <= _1687;
        160:
            _4708 <= _1678;
        161:
            _4708 <= _1669;
        162:
            _4708 <= _1660;
        163:
            _4708 <= _1651;
        164:
            _4708 <= _1642;
        165:
            _4708 <= _1633;
        166:
            _4708 <= _1624;
        167:
            _4708 <= _1615;
        168:
            _4708 <= _1606;
        169:
            _4708 <= _1597;
        170:
            _4708 <= _1588;
        171:
            _4708 <= _1579;
        172:
            _4708 <= _1570;
        173:
            _4708 <= _1561;
        174:
            _4708 <= _1552;
        175:
            _4708 <= _1543;
        176:
            _4708 <= _1534;
        177:
            _4708 <= _1525;
        178:
            _4708 <= _1516;
        179:
            _4708 <= _1507;
        180:
            _4708 <= _1498;
        181:
            _4708 <= _1489;
        182:
            _4708 <= _1480;
        183:
            _4708 <= _1471;
        184:
            _4708 <= _1462;
        185:
            _4708 <= _1453;
        186:
            _4708 <= _1444;
        187:
            _4708 <= _1435;
        188:
            _4708 <= _1426;
        189:
            _4708 <= _1417;
        190:
            _4708 <= _1408;
        191:
            _4708 <= _1399;
        192:
            _4708 <= _1390;
        193:
            _4708 <= _1381;
        194:
            _4708 <= _1372;
        195:
            _4708 <= _1363;
        196:
            _4708 <= _1354;
        197:
            _4708 <= _1345;
        198:
            _4708 <= _1336;
        199:
            _4708 <= _1327;
        200:
            _4708 <= _1318;
        201:
            _4708 <= _1309;
        202:
            _4708 <= _1300;
        203:
            _4708 <= _1291;
        204:
            _4708 <= _1282;
        205:
            _4708 <= _1273;
        206:
            _4708 <= _1264;
        207:
            _4708 <= _1255;
        208:
            _4708 <= _1246;
        209:
            _4708 <= _1237;
        210:
            _4708 <= _1228;
        211:
            _4708 <= _1219;
        212:
            _4708 <= _1210;
        213:
            _4708 <= _1201;
        214:
            _4708 <= _1192;
        215:
            _4708 <= _1183;
        216:
            _4708 <= _1174;
        217:
            _4708 <= _1165;
        218:
            _4708 <= _1156;
        219:
            _4708 <= _1147;
        220:
            _4708 <= _1138;
        221:
            _4708 <= _1129;
        222:
            _4708 <= _1120;
        223:
            _4708 <= _1111;
        224:
            _4708 <= _1102;
        225:
            _4708 <= _1093;
        226:
            _4708 <= _1084;
        227:
            _4708 <= _1075;
        228:
            _4708 <= _1066;
        229:
            _4708 <= _1057;
        230:
            _4708 <= _1048;
        231:
            _4708 <= _1039;
        232:
            _4708 <= _1030;
        233:
            _4708 <= _1021;
        234:
            _4708 <= _1012;
        235:
            _4708 <= _1003;
        236:
            _4708 <= _994;
        237:
            _4708 <= _985;
        238:
            _4708 <= _976;
        239:
            _4708 <= _967;
        240:
            _4708 <= _958;
        241:
            _4708 <= _949;
        242:
            _4708 <= _940;
        243:
            _4708 <= _931;
        244:
            _4708 <= _922;
        245:
            _4708 <= _913;
        246:
            _4708 <= _904;
        247:
            _4708 <= _895;
        248:
            _4708 <= _886;
        249:
            _4708 <= _877;
        250:
            _4708 <= _868;
        251:
            _4708 <= _859;
        252:
            _4708 <= _850;
        253:
            _4708 <= _841;
        254:
            _4708 <= _832;
        default:
            _4708 <= _823;
        endcase
    end
    assign _4707 = 32'b00000000000000000000000000000000;
    assign _4709 = { _4707,
                     _4708 };
    assign _818 = 8'b11111111;
    assign _819 = _817 == _818;
    assign _820 = _814 & _819;
    assign _824 = _820 ? _258 : _823;
    assign _826 = _805 ? _4707 : _824;
    assign _2 = _826;
    always @(posedge _791) begin
        if (_789)
            _823 <= _4707;
        else
            _823 <= _2;
    end
    assign _827 = 8'b11111110;
    assign _828 = _817 == _827;
    assign _829 = _814 & _828;
    assign _833 = _829 ? _258 : _832;
    assign _835 = _805 ? _4707 : _833;
    assign _3 = _835;
    always @(posedge _791) begin
        if (_789)
            _832 <= _4707;
        else
            _832 <= _3;
    end
    assign _836 = 8'b11111101;
    assign _837 = _817 == _836;
    assign _838 = _814 & _837;
    assign _842 = _838 ? _258 : _841;
    assign _844 = _805 ? _4707 : _842;
    assign _4 = _844;
    always @(posedge _791) begin
        if (_789)
            _841 <= _4707;
        else
            _841 <= _4;
    end
    assign _845 = 8'b11111100;
    assign _846 = _817 == _845;
    assign _847 = _814 & _846;
    assign _851 = _847 ? _258 : _850;
    assign _853 = _805 ? _4707 : _851;
    assign _5 = _853;
    always @(posedge _791) begin
        if (_789)
            _850 <= _4707;
        else
            _850 <= _5;
    end
    assign _854 = 8'b11111011;
    assign _855 = _817 == _854;
    assign _856 = _814 & _855;
    assign _860 = _856 ? _258 : _859;
    assign _862 = _805 ? _4707 : _860;
    assign _6 = _862;
    always @(posedge _791) begin
        if (_789)
            _859 <= _4707;
        else
            _859 <= _6;
    end
    assign _863 = 8'b11111010;
    assign _864 = _817 == _863;
    assign _865 = _814 & _864;
    assign _869 = _865 ? _258 : _868;
    assign _871 = _805 ? _4707 : _869;
    assign _7 = _871;
    always @(posedge _791) begin
        if (_789)
            _868 <= _4707;
        else
            _868 <= _7;
    end
    assign _872 = 8'b11111001;
    assign _873 = _817 == _872;
    assign _874 = _814 & _873;
    assign _878 = _874 ? _258 : _877;
    assign _880 = _805 ? _4707 : _878;
    assign _8 = _880;
    always @(posedge _791) begin
        if (_789)
            _877 <= _4707;
        else
            _877 <= _8;
    end
    assign _881 = 8'b11111000;
    assign _882 = _817 == _881;
    assign _883 = _814 & _882;
    assign _887 = _883 ? _258 : _886;
    assign _889 = _805 ? _4707 : _887;
    assign _9 = _889;
    always @(posedge _791) begin
        if (_789)
            _886 <= _4707;
        else
            _886 <= _9;
    end
    assign _890 = 8'b11110111;
    assign _891 = _817 == _890;
    assign _892 = _814 & _891;
    assign _896 = _892 ? _258 : _895;
    assign _898 = _805 ? _4707 : _896;
    assign _10 = _898;
    always @(posedge _791) begin
        if (_789)
            _895 <= _4707;
        else
            _895 <= _10;
    end
    assign _899 = 8'b11110110;
    assign _900 = _817 == _899;
    assign _901 = _814 & _900;
    assign _905 = _901 ? _258 : _904;
    assign _907 = _805 ? _4707 : _905;
    assign _11 = _907;
    always @(posedge _791) begin
        if (_789)
            _904 <= _4707;
        else
            _904 <= _11;
    end
    assign _908 = 8'b11110101;
    assign _909 = _817 == _908;
    assign _910 = _814 & _909;
    assign _914 = _910 ? _258 : _913;
    assign _916 = _805 ? _4707 : _914;
    assign _12 = _916;
    always @(posedge _791) begin
        if (_789)
            _913 <= _4707;
        else
            _913 <= _12;
    end
    assign _917 = 8'b11110100;
    assign _918 = _817 == _917;
    assign _919 = _814 & _918;
    assign _923 = _919 ? _258 : _922;
    assign _925 = _805 ? _4707 : _923;
    assign _13 = _925;
    always @(posedge _791) begin
        if (_789)
            _922 <= _4707;
        else
            _922 <= _13;
    end
    assign _926 = 8'b11110011;
    assign _927 = _817 == _926;
    assign _928 = _814 & _927;
    assign _932 = _928 ? _258 : _931;
    assign _934 = _805 ? _4707 : _932;
    assign _14 = _934;
    always @(posedge _791) begin
        if (_789)
            _931 <= _4707;
        else
            _931 <= _14;
    end
    assign _935 = 8'b11110010;
    assign _936 = _817 == _935;
    assign _937 = _814 & _936;
    assign _941 = _937 ? _258 : _940;
    assign _943 = _805 ? _4707 : _941;
    assign _15 = _943;
    always @(posedge _791) begin
        if (_789)
            _940 <= _4707;
        else
            _940 <= _15;
    end
    assign _944 = 8'b11110001;
    assign _945 = _817 == _944;
    assign _946 = _814 & _945;
    assign _950 = _946 ? _258 : _949;
    assign _952 = _805 ? _4707 : _950;
    assign _16 = _952;
    always @(posedge _791) begin
        if (_789)
            _949 <= _4707;
        else
            _949 <= _16;
    end
    assign _953 = 8'b11110000;
    assign _954 = _817 == _953;
    assign _955 = _814 & _954;
    assign _959 = _955 ? _258 : _958;
    assign _961 = _805 ? _4707 : _959;
    assign _17 = _961;
    always @(posedge _791) begin
        if (_789)
            _958 <= _4707;
        else
            _958 <= _17;
    end
    assign _962 = 8'b11101111;
    assign _963 = _817 == _962;
    assign _964 = _814 & _963;
    assign _968 = _964 ? _258 : _967;
    assign _970 = _805 ? _4707 : _968;
    assign _18 = _970;
    always @(posedge _791) begin
        if (_789)
            _967 <= _4707;
        else
            _967 <= _18;
    end
    assign _971 = 8'b11101110;
    assign _972 = _817 == _971;
    assign _973 = _814 & _972;
    assign _977 = _973 ? _258 : _976;
    assign _979 = _805 ? _4707 : _977;
    assign _19 = _979;
    always @(posedge _791) begin
        if (_789)
            _976 <= _4707;
        else
            _976 <= _19;
    end
    assign _980 = 8'b11101101;
    assign _981 = _817 == _980;
    assign _982 = _814 & _981;
    assign _986 = _982 ? _258 : _985;
    assign _988 = _805 ? _4707 : _986;
    assign _20 = _988;
    always @(posedge _791) begin
        if (_789)
            _985 <= _4707;
        else
            _985 <= _20;
    end
    assign _989 = 8'b11101100;
    assign _990 = _817 == _989;
    assign _991 = _814 & _990;
    assign _995 = _991 ? _258 : _994;
    assign _997 = _805 ? _4707 : _995;
    assign _21 = _997;
    always @(posedge _791) begin
        if (_789)
            _994 <= _4707;
        else
            _994 <= _21;
    end
    assign _998 = 8'b11101011;
    assign _999 = _817 == _998;
    assign _1000 = _814 & _999;
    assign _1004 = _1000 ? _258 : _1003;
    assign _1006 = _805 ? _4707 : _1004;
    assign _22 = _1006;
    always @(posedge _791) begin
        if (_789)
            _1003 <= _4707;
        else
            _1003 <= _22;
    end
    assign _1007 = 8'b11101010;
    assign _1008 = _817 == _1007;
    assign _1009 = _814 & _1008;
    assign _1013 = _1009 ? _258 : _1012;
    assign _1015 = _805 ? _4707 : _1013;
    assign _23 = _1015;
    always @(posedge _791) begin
        if (_789)
            _1012 <= _4707;
        else
            _1012 <= _23;
    end
    assign _1016 = 8'b11101001;
    assign _1017 = _817 == _1016;
    assign _1018 = _814 & _1017;
    assign _1022 = _1018 ? _258 : _1021;
    assign _1024 = _805 ? _4707 : _1022;
    assign _24 = _1024;
    always @(posedge _791) begin
        if (_789)
            _1021 <= _4707;
        else
            _1021 <= _24;
    end
    assign _1025 = 8'b11101000;
    assign _1026 = _817 == _1025;
    assign _1027 = _814 & _1026;
    assign _1031 = _1027 ? _258 : _1030;
    assign _1033 = _805 ? _4707 : _1031;
    assign _25 = _1033;
    always @(posedge _791) begin
        if (_789)
            _1030 <= _4707;
        else
            _1030 <= _25;
    end
    assign _1034 = 8'b11100111;
    assign _1035 = _817 == _1034;
    assign _1036 = _814 & _1035;
    assign _1040 = _1036 ? _258 : _1039;
    assign _1042 = _805 ? _4707 : _1040;
    assign _26 = _1042;
    always @(posedge _791) begin
        if (_789)
            _1039 <= _4707;
        else
            _1039 <= _26;
    end
    assign _1043 = 8'b11100110;
    assign _1044 = _817 == _1043;
    assign _1045 = _814 & _1044;
    assign _1049 = _1045 ? _258 : _1048;
    assign _1051 = _805 ? _4707 : _1049;
    assign _27 = _1051;
    always @(posedge _791) begin
        if (_789)
            _1048 <= _4707;
        else
            _1048 <= _27;
    end
    assign _1052 = 8'b11100101;
    assign _1053 = _817 == _1052;
    assign _1054 = _814 & _1053;
    assign _1058 = _1054 ? _258 : _1057;
    assign _1060 = _805 ? _4707 : _1058;
    assign _28 = _1060;
    always @(posedge _791) begin
        if (_789)
            _1057 <= _4707;
        else
            _1057 <= _28;
    end
    assign _1061 = 8'b11100100;
    assign _1062 = _817 == _1061;
    assign _1063 = _814 & _1062;
    assign _1067 = _1063 ? _258 : _1066;
    assign _1069 = _805 ? _4707 : _1067;
    assign _29 = _1069;
    always @(posedge _791) begin
        if (_789)
            _1066 <= _4707;
        else
            _1066 <= _29;
    end
    assign _1070 = 8'b11100011;
    assign _1071 = _817 == _1070;
    assign _1072 = _814 & _1071;
    assign _1076 = _1072 ? _258 : _1075;
    assign _1078 = _805 ? _4707 : _1076;
    assign _30 = _1078;
    always @(posedge _791) begin
        if (_789)
            _1075 <= _4707;
        else
            _1075 <= _30;
    end
    assign _1079 = 8'b11100010;
    assign _1080 = _817 == _1079;
    assign _1081 = _814 & _1080;
    assign _1085 = _1081 ? _258 : _1084;
    assign _1087 = _805 ? _4707 : _1085;
    assign _31 = _1087;
    always @(posedge _791) begin
        if (_789)
            _1084 <= _4707;
        else
            _1084 <= _31;
    end
    assign _1088 = 8'b11100001;
    assign _1089 = _817 == _1088;
    assign _1090 = _814 & _1089;
    assign _1094 = _1090 ? _258 : _1093;
    assign _1096 = _805 ? _4707 : _1094;
    assign _32 = _1096;
    always @(posedge _791) begin
        if (_789)
            _1093 <= _4707;
        else
            _1093 <= _32;
    end
    assign _1097 = 8'b11100000;
    assign _1098 = _817 == _1097;
    assign _1099 = _814 & _1098;
    assign _1103 = _1099 ? _258 : _1102;
    assign _1105 = _805 ? _4707 : _1103;
    assign _33 = _1105;
    always @(posedge _791) begin
        if (_789)
            _1102 <= _4707;
        else
            _1102 <= _33;
    end
    assign _1106 = 8'b11011111;
    assign _1107 = _817 == _1106;
    assign _1108 = _814 & _1107;
    assign _1112 = _1108 ? _258 : _1111;
    assign _1114 = _805 ? _4707 : _1112;
    assign _34 = _1114;
    always @(posedge _791) begin
        if (_789)
            _1111 <= _4707;
        else
            _1111 <= _34;
    end
    assign _1115 = 8'b11011110;
    assign _1116 = _817 == _1115;
    assign _1117 = _814 & _1116;
    assign _1121 = _1117 ? _258 : _1120;
    assign _1123 = _805 ? _4707 : _1121;
    assign _35 = _1123;
    always @(posedge _791) begin
        if (_789)
            _1120 <= _4707;
        else
            _1120 <= _35;
    end
    assign _1124 = 8'b11011101;
    assign _1125 = _817 == _1124;
    assign _1126 = _814 & _1125;
    assign _1130 = _1126 ? _258 : _1129;
    assign _1132 = _805 ? _4707 : _1130;
    assign _36 = _1132;
    always @(posedge _791) begin
        if (_789)
            _1129 <= _4707;
        else
            _1129 <= _36;
    end
    assign _1133 = 8'b11011100;
    assign _1134 = _817 == _1133;
    assign _1135 = _814 & _1134;
    assign _1139 = _1135 ? _258 : _1138;
    assign _1141 = _805 ? _4707 : _1139;
    assign _37 = _1141;
    always @(posedge _791) begin
        if (_789)
            _1138 <= _4707;
        else
            _1138 <= _37;
    end
    assign _1142 = 8'b11011011;
    assign _1143 = _817 == _1142;
    assign _1144 = _814 & _1143;
    assign _1148 = _1144 ? _258 : _1147;
    assign _1150 = _805 ? _4707 : _1148;
    assign _38 = _1150;
    always @(posedge _791) begin
        if (_789)
            _1147 <= _4707;
        else
            _1147 <= _38;
    end
    assign _1151 = 8'b11011010;
    assign _1152 = _817 == _1151;
    assign _1153 = _814 & _1152;
    assign _1157 = _1153 ? _258 : _1156;
    assign _1159 = _805 ? _4707 : _1157;
    assign _39 = _1159;
    always @(posedge _791) begin
        if (_789)
            _1156 <= _4707;
        else
            _1156 <= _39;
    end
    assign _1160 = 8'b11011001;
    assign _1161 = _817 == _1160;
    assign _1162 = _814 & _1161;
    assign _1166 = _1162 ? _258 : _1165;
    assign _1168 = _805 ? _4707 : _1166;
    assign _40 = _1168;
    always @(posedge _791) begin
        if (_789)
            _1165 <= _4707;
        else
            _1165 <= _40;
    end
    assign _1169 = 8'b11011000;
    assign _1170 = _817 == _1169;
    assign _1171 = _814 & _1170;
    assign _1175 = _1171 ? _258 : _1174;
    assign _1177 = _805 ? _4707 : _1175;
    assign _41 = _1177;
    always @(posedge _791) begin
        if (_789)
            _1174 <= _4707;
        else
            _1174 <= _41;
    end
    assign _1178 = 8'b11010111;
    assign _1179 = _817 == _1178;
    assign _1180 = _814 & _1179;
    assign _1184 = _1180 ? _258 : _1183;
    assign _1186 = _805 ? _4707 : _1184;
    assign _42 = _1186;
    always @(posedge _791) begin
        if (_789)
            _1183 <= _4707;
        else
            _1183 <= _42;
    end
    assign _1187 = 8'b11010110;
    assign _1188 = _817 == _1187;
    assign _1189 = _814 & _1188;
    assign _1193 = _1189 ? _258 : _1192;
    assign _1195 = _805 ? _4707 : _1193;
    assign _43 = _1195;
    always @(posedge _791) begin
        if (_789)
            _1192 <= _4707;
        else
            _1192 <= _43;
    end
    assign _1196 = 8'b11010101;
    assign _1197 = _817 == _1196;
    assign _1198 = _814 & _1197;
    assign _1202 = _1198 ? _258 : _1201;
    assign _1204 = _805 ? _4707 : _1202;
    assign _44 = _1204;
    always @(posedge _791) begin
        if (_789)
            _1201 <= _4707;
        else
            _1201 <= _44;
    end
    assign _1205 = 8'b11010100;
    assign _1206 = _817 == _1205;
    assign _1207 = _814 & _1206;
    assign _1211 = _1207 ? _258 : _1210;
    assign _1213 = _805 ? _4707 : _1211;
    assign _45 = _1213;
    always @(posedge _791) begin
        if (_789)
            _1210 <= _4707;
        else
            _1210 <= _45;
    end
    assign _1214 = 8'b11010011;
    assign _1215 = _817 == _1214;
    assign _1216 = _814 & _1215;
    assign _1220 = _1216 ? _258 : _1219;
    assign _1222 = _805 ? _4707 : _1220;
    assign _46 = _1222;
    always @(posedge _791) begin
        if (_789)
            _1219 <= _4707;
        else
            _1219 <= _46;
    end
    assign _1223 = 8'b11010010;
    assign _1224 = _817 == _1223;
    assign _1225 = _814 & _1224;
    assign _1229 = _1225 ? _258 : _1228;
    assign _1231 = _805 ? _4707 : _1229;
    assign _47 = _1231;
    always @(posedge _791) begin
        if (_789)
            _1228 <= _4707;
        else
            _1228 <= _47;
    end
    assign _1232 = 8'b11010001;
    assign _1233 = _817 == _1232;
    assign _1234 = _814 & _1233;
    assign _1238 = _1234 ? _258 : _1237;
    assign _1240 = _805 ? _4707 : _1238;
    assign _48 = _1240;
    always @(posedge _791) begin
        if (_789)
            _1237 <= _4707;
        else
            _1237 <= _48;
    end
    assign _1241 = 8'b11010000;
    assign _1242 = _817 == _1241;
    assign _1243 = _814 & _1242;
    assign _1247 = _1243 ? _258 : _1246;
    assign _1249 = _805 ? _4707 : _1247;
    assign _49 = _1249;
    always @(posedge _791) begin
        if (_789)
            _1246 <= _4707;
        else
            _1246 <= _49;
    end
    assign _1250 = 8'b11001111;
    assign _1251 = _817 == _1250;
    assign _1252 = _814 & _1251;
    assign _1256 = _1252 ? _258 : _1255;
    assign _1258 = _805 ? _4707 : _1256;
    assign _50 = _1258;
    always @(posedge _791) begin
        if (_789)
            _1255 <= _4707;
        else
            _1255 <= _50;
    end
    assign _1259 = 8'b11001110;
    assign _1260 = _817 == _1259;
    assign _1261 = _814 & _1260;
    assign _1265 = _1261 ? _258 : _1264;
    assign _1267 = _805 ? _4707 : _1265;
    assign _51 = _1267;
    always @(posedge _791) begin
        if (_789)
            _1264 <= _4707;
        else
            _1264 <= _51;
    end
    assign _1268 = 8'b11001101;
    assign _1269 = _817 == _1268;
    assign _1270 = _814 & _1269;
    assign _1274 = _1270 ? _258 : _1273;
    assign _1276 = _805 ? _4707 : _1274;
    assign _52 = _1276;
    always @(posedge _791) begin
        if (_789)
            _1273 <= _4707;
        else
            _1273 <= _52;
    end
    assign _1277 = 8'b11001100;
    assign _1278 = _817 == _1277;
    assign _1279 = _814 & _1278;
    assign _1283 = _1279 ? _258 : _1282;
    assign _1285 = _805 ? _4707 : _1283;
    assign _53 = _1285;
    always @(posedge _791) begin
        if (_789)
            _1282 <= _4707;
        else
            _1282 <= _53;
    end
    assign _1286 = 8'b11001011;
    assign _1287 = _817 == _1286;
    assign _1288 = _814 & _1287;
    assign _1292 = _1288 ? _258 : _1291;
    assign _1294 = _805 ? _4707 : _1292;
    assign _54 = _1294;
    always @(posedge _791) begin
        if (_789)
            _1291 <= _4707;
        else
            _1291 <= _54;
    end
    assign _1295 = 8'b11001010;
    assign _1296 = _817 == _1295;
    assign _1297 = _814 & _1296;
    assign _1301 = _1297 ? _258 : _1300;
    assign _1303 = _805 ? _4707 : _1301;
    assign _55 = _1303;
    always @(posedge _791) begin
        if (_789)
            _1300 <= _4707;
        else
            _1300 <= _55;
    end
    assign _1304 = 8'b11001001;
    assign _1305 = _817 == _1304;
    assign _1306 = _814 & _1305;
    assign _1310 = _1306 ? _258 : _1309;
    assign _1312 = _805 ? _4707 : _1310;
    assign _56 = _1312;
    always @(posedge _791) begin
        if (_789)
            _1309 <= _4707;
        else
            _1309 <= _56;
    end
    assign _1313 = 8'b11001000;
    assign _1314 = _817 == _1313;
    assign _1315 = _814 & _1314;
    assign _1319 = _1315 ? _258 : _1318;
    assign _1321 = _805 ? _4707 : _1319;
    assign _57 = _1321;
    always @(posedge _791) begin
        if (_789)
            _1318 <= _4707;
        else
            _1318 <= _57;
    end
    assign _1322 = 8'b11000111;
    assign _1323 = _817 == _1322;
    assign _1324 = _814 & _1323;
    assign _1328 = _1324 ? _258 : _1327;
    assign _1330 = _805 ? _4707 : _1328;
    assign _58 = _1330;
    always @(posedge _791) begin
        if (_789)
            _1327 <= _4707;
        else
            _1327 <= _58;
    end
    assign _1331 = 8'b11000110;
    assign _1332 = _817 == _1331;
    assign _1333 = _814 & _1332;
    assign _1337 = _1333 ? _258 : _1336;
    assign _1339 = _805 ? _4707 : _1337;
    assign _59 = _1339;
    always @(posedge _791) begin
        if (_789)
            _1336 <= _4707;
        else
            _1336 <= _59;
    end
    assign _1340 = 8'b11000101;
    assign _1341 = _817 == _1340;
    assign _1342 = _814 & _1341;
    assign _1346 = _1342 ? _258 : _1345;
    assign _1348 = _805 ? _4707 : _1346;
    assign _60 = _1348;
    always @(posedge _791) begin
        if (_789)
            _1345 <= _4707;
        else
            _1345 <= _60;
    end
    assign _1349 = 8'b11000100;
    assign _1350 = _817 == _1349;
    assign _1351 = _814 & _1350;
    assign _1355 = _1351 ? _258 : _1354;
    assign _1357 = _805 ? _4707 : _1355;
    assign _61 = _1357;
    always @(posedge _791) begin
        if (_789)
            _1354 <= _4707;
        else
            _1354 <= _61;
    end
    assign _1358 = 8'b11000011;
    assign _1359 = _817 == _1358;
    assign _1360 = _814 & _1359;
    assign _1364 = _1360 ? _258 : _1363;
    assign _1366 = _805 ? _4707 : _1364;
    assign _62 = _1366;
    always @(posedge _791) begin
        if (_789)
            _1363 <= _4707;
        else
            _1363 <= _62;
    end
    assign _1367 = 8'b11000010;
    assign _1368 = _817 == _1367;
    assign _1369 = _814 & _1368;
    assign _1373 = _1369 ? _258 : _1372;
    assign _1375 = _805 ? _4707 : _1373;
    assign _63 = _1375;
    always @(posedge _791) begin
        if (_789)
            _1372 <= _4707;
        else
            _1372 <= _63;
    end
    assign _1376 = 8'b11000001;
    assign _1377 = _817 == _1376;
    assign _1378 = _814 & _1377;
    assign _1382 = _1378 ? _258 : _1381;
    assign _1384 = _805 ? _4707 : _1382;
    assign _64 = _1384;
    always @(posedge _791) begin
        if (_789)
            _1381 <= _4707;
        else
            _1381 <= _64;
    end
    assign _1385 = 8'b11000000;
    assign _1386 = _817 == _1385;
    assign _1387 = _814 & _1386;
    assign _1391 = _1387 ? _258 : _1390;
    assign _1393 = _805 ? _4707 : _1391;
    assign _65 = _1393;
    always @(posedge _791) begin
        if (_789)
            _1390 <= _4707;
        else
            _1390 <= _65;
    end
    assign _1394 = 8'b10111111;
    assign _1395 = _817 == _1394;
    assign _1396 = _814 & _1395;
    assign _1400 = _1396 ? _258 : _1399;
    assign _1402 = _805 ? _4707 : _1400;
    assign _66 = _1402;
    always @(posedge _791) begin
        if (_789)
            _1399 <= _4707;
        else
            _1399 <= _66;
    end
    assign _1403 = 8'b10111110;
    assign _1404 = _817 == _1403;
    assign _1405 = _814 & _1404;
    assign _1409 = _1405 ? _258 : _1408;
    assign _1411 = _805 ? _4707 : _1409;
    assign _67 = _1411;
    always @(posedge _791) begin
        if (_789)
            _1408 <= _4707;
        else
            _1408 <= _67;
    end
    assign _1412 = 8'b10111101;
    assign _1413 = _817 == _1412;
    assign _1414 = _814 & _1413;
    assign _1418 = _1414 ? _258 : _1417;
    assign _1420 = _805 ? _4707 : _1418;
    assign _68 = _1420;
    always @(posedge _791) begin
        if (_789)
            _1417 <= _4707;
        else
            _1417 <= _68;
    end
    assign _1421 = 8'b10111100;
    assign _1422 = _817 == _1421;
    assign _1423 = _814 & _1422;
    assign _1427 = _1423 ? _258 : _1426;
    assign _1429 = _805 ? _4707 : _1427;
    assign _69 = _1429;
    always @(posedge _791) begin
        if (_789)
            _1426 <= _4707;
        else
            _1426 <= _69;
    end
    assign _1430 = 8'b10111011;
    assign _1431 = _817 == _1430;
    assign _1432 = _814 & _1431;
    assign _1436 = _1432 ? _258 : _1435;
    assign _1438 = _805 ? _4707 : _1436;
    assign _70 = _1438;
    always @(posedge _791) begin
        if (_789)
            _1435 <= _4707;
        else
            _1435 <= _70;
    end
    assign _1439 = 8'b10111010;
    assign _1440 = _817 == _1439;
    assign _1441 = _814 & _1440;
    assign _1445 = _1441 ? _258 : _1444;
    assign _1447 = _805 ? _4707 : _1445;
    assign _71 = _1447;
    always @(posedge _791) begin
        if (_789)
            _1444 <= _4707;
        else
            _1444 <= _71;
    end
    assign _1448 = 8'b10111001;
    assign _1449 = _817 == _1448;
    assign _1450 = _814 & _1449;
    assign _1454 = _1450 ? _258 : _1453;
    assign _1456 = _805 ? _4707 : _1454;
    assign _72 = _1456;
    always @(posedge _791) begin
        if (_789)
            _1453 <= _4707;
        else
            _1453 <= _72;
    end
    assign _1457 = 8'b10111000;
    assign _1458 = _817 == _1457;
    assign _1459 = _814 & _1458;
    assign _1463 = _1459 ? _258 : _1462;
    assign _1465 = _805 ? _4707 : _1463;
    assign _73 = _1465;
    always @(posedge _791) begin
        if (_789)
            _1462 <= _4707;
        else
            _1462 <= _73;
    end
    assign _1466 = 8'b10110111;
    assign _1467 = _817 == _1466;
    assign _1468 = _814 & _1467;
    assign _1472 = _1468 ? _258 : _1471;
    assign _1474 = _805 ? _4707 : _1472;
    assign _74 = _1474;
    always @(posedge _791) begin
        if (_789)
            _1471 <= _4707;
        else
            _1471 <= _74;
    end
    assign _1475 = 8'b10110110;
    assign _1476 = _817 == _1475;
    assign _1477 = _814 & _1476;
    assign _1481 = _1477 ? _258 : _1480;
    assign _1483 = _805 ? _4707 : _1481;
    assign _75 = _1483;
    always @(posedge _791) begin
        if (_789)
            _1480 <= _4707;
        else
            _1480 <= _75;
    end
    assign _1484 = 8'b10110101;
    assign _1485 = _817 == _1484;
    assign _1486 = _814 & _1485;
    assign _1490 = _1486 ? _258 : _1489;
    assign _1492 = _805 ? _4707 : _1490;
    assign _76 = _1492;
    always @(posedge _791) begin
        if (_789)
            _1489 <= _4707;
        else
            _1489 <= _76;
    end
    assign _1493 = 8'b10110100;
    assign _1494 = _817 == _1493;
    assign _1495 = _814 & _1494;
    assign _1499 = _1495 ? _258 : _1498;
    assign _1501 = _805 ? _4707 : _1499;
    assign _77 = _1501;
    always @(posedge _791) begin
        if (_789)
            _1498 <= _4707;
        else
            _1498 <= _77;
    end
    assign _1502 = 8'b10110011;
    assign _1503 = _817 == _1502;
    assign _1504 = _814 & _1503;
    assign _1508 = _1504 ? _258 : _1507;
    assign _1510 = _805 ? _4707 : _1508;
    assign _78 = _1510;
    always @(posedge _791) begin
        if (_789)
            _1507 <= _4707;
        else
            _1507 <= _78;
    end
    assign _1511 = 8'b10110010;
    assign _1512 = _817 == _1511;
    assign _1513 = _814 & _1512;
    assign _1517 = _1513 ? _258 : _1516;
    assign _1519 = _805 ? _4707 : _1517;
    assign _79 = _1519;
    always @(posedge _791) begin
        if (_789)
            _1516 <= _4707;
        else
            _1516 <= _79;
    end
    assign _1520 = 8'b10110001;
    assign _1521 = _817 == _1520;
    assign _1522 = _814 & _1521;
    assign _1526 = _1522 ? _258 : _1525;
    assign _1528 = _805 ? _4707 : _1526;
    assign _80 = _1528;
    always @(posedge _791) begin
        if (_789)
            _1525 <= _4707;
        else
            _1525 <= _80;
    end
    assign _1529 = 8'b10110000;
    assign _1530 = _817 == _1529;
    assign _1531 = _814 & _1530;
    assign _1535 = _1531 ? _258 : _1534;
    assign _1537 = _805 ? _4707 : _1535;
    assign _81 = _1537;
    always @(posedge _791) begin
        if (_789)
            _1534 <= _4707;
        else
            _1534 <= _81;
    end
    assign _1538 = 8'b10101111;
    assign _1539 = _817 == _1538;
    assign _1540 = _814 & _1539;
    assign _1544 = _1540 ? _258 : _1543;
    assign _1546 = _805 ? _4707 : _1544;
    assign _82 = _1546;
    always @(posedge _791) begin
        if (_789)
            _1543 <= _4707;
        else
            _1543 <= _82;
    end
    assign _1547 = 8'b10101110;
    assign _1548 = _817 == _1547;
    assign _1549 = _814 & _1548;
    assign _1553 = _1549 ? _258 : _1552;
    assign _1555 = _805 ? _4707 : _1553;
    assign _83 = _1555;
    always @(posedge _791) begin
        if (_789)
            _1552 <= _4707;
        else
            _1552 <= _83;
    end
    assign _1556 = 8'b10101101;
    assign _1557 = _817 == _1556;
    assign _1558 = _814 & _1557;
    assign _1562 = _1558 ? _258 : _1561;
    assign _1564 = _805 ? _4707 : _1562;
    assign _84 = _1564;
    always @(posedge _791) begin
        if (_789)
            _1561 <= _4707;
        else
            _1561 <= _84;
    end
    assign _1565 = 8'b10101100;
    assign _1566 = _817 == _1565;
    assign _1567 = _814 & _1566;
    assign _1571 = _1567 ? _258 : _1570;
    assign _1573 = _805 ? _4707 : _1571;
    assign _85 = _1573;
    always @(posedge _791) begin
        if (_789)
            _1570 <= _4707;
        else
            _1570 <= _85;
    end
    assign _1574 = 8'b10101011;
    assign _1575 = _817 == _1574;
    assign _1576 = _814 & _1575;
    assign _1580 = _1576 ? _258 : _1579;
    assign _1582 = _805 ? _4707 : _1580;
    assign _86 = _1582;
    always @(posedge _791) begin
        if (_789)
            _1579 <= _4707;
        else
            _1579 <= _86;
    end
    assign _1583 = 8'b10101010;
    assign _1584 = _817 == _1583;
    assign _1585 = _814 & _1584;
    assign _1589 = _1585 ? _258 : _1588;
    assign _1591 = _805 ? _4707 : _1589;
    assign _87 = _1591;
    always @(posedge _791) begin
        if (_789)
            _1588 <= _4707;
        else
            _1588 <= _87;
    end
    assign _1592 = 8'b10101001;
    assign _1593 = _817 == _1592;
    assign _1594 = _814 & _1593;
    assign _1598 = _1594 ? _258 : _1597;
    assign _1600 = _805 ? _4707 : _1598;
    assign _88 = _1600;
    always @(posedge _791) begin
        if (_789)
            _1597 <= _4707;
        else
            _1597 <= _88;
    end
    assign _1601 = 8'b10101000;
    assign _1602 = _817 == _1601;
    assign _1603 = _814 & _1602;
    assign _1607 = _1603 ? _258 : _1606;
    assign _1609 = _805 ? _4707 : _1607;
    assign _89 = _1609;
    always @(posedge _791) begin
        if (_789)
            _1606 <= _4707;
        else
            _1606 <= _89;
    end
    assign _1610 = 8'b10100111;
    assign _1611 = _817 == _1610;
    assign _1612 = _814 & _1611;
    assign _1616 = _1612 ? _258 : _1615;
    assign _1618 = _805 ? _4707 : _1616;
    assign _90 = _1618;
    always @(posedge _791) begin
        if (_789)
            _1615 <= _4707;
        else
            _1615 <= _90;
    end
    assign _1619 = 8'b10100110;
    assign _1620 = _817 == _1619;
    assign _1621 = _814 & _1620;
    assign _1625 = _1621 ? _258 : _1624;
    assign _1627 = _805 ? _4707 : _1625;
    assign _91 = _1627;
    always @(posedge _791) begin
        if (_789)
            _1624 <= _4707;
        else
            _1624 <= _91;
    end
    assign _1628 = 8'b10100101;
    assign _1629 = _817 == _1628;
    assign _1630 = _814 & _1629;
    assign _1634 = _1630 ? _258 : _1633;
    assign _1636 = _805 ? _4707 : _1634;
    assign _92 = _1636;
    always @(posedge _791) begin
        if (_789)
            _1633 <= _4707;
        else
            _1633 <= _92;
    end
    assign _1637 = 8'b10100100;
    assign _1638 = _817 == _1637;
    assign _1639 = _814 & _1638;
    assign _1643 = _1639 ? _258 : _1642;
    assign _1645 = _805 ? _4707 : _1643;
    assign _93 = _1645;
    always @(posedge _791) begin
        if (_789)
            _1642 <= _4707;
        else
            _1642 <= _93;
    end
    assign _1646 = 8'b10100011;
    assign _1647 = _817 == _1646;
    assign _1648 = _814 & _1647;
    assign _1652 = _1648 ? _258 : _1651;
    assign _1654 = _805 ? _4707 : _1652;
    assign _94 = _1654;
    always @(posedge _791) begin
        if (_789)
            _1651 <= _4707;
        else
            _1651 <= _94;
    end
    assign _1655 = 8'b10100010;
    assign _1656 = _817 == _1655;
    assign _1657 = _814 & _1656;
    assign _1661 = _1657 ? _258 : _1660;
    assign _1663 = _805 ? _4707 : _1661;
    assign _95 = _1663;
    always @(posedge _791) begin
        if (_789)
            _1660 <= _4707;
        else
            _1660 <= _95;
    end
    assign _1664 = 8'b10100001;
    assign _1665 = _817 == _1664;
    assign _1666 = _814 & _1665;
    assign _1670 = _1666 ? _258 : _1669;
    assign _1672 = _805 ? _4707 : _1670;
    assign _96 = _1672;
    always @(posedge _791) begin
        if (_789)
            _1669 <= _4707;
        else
            _1669 <= _96;
    end
    assign _1673 = 8'b10100000;
    assign _1674 = _817 == _1673;
    assign _1675 = _814 & _1674;
    assign _1679 = _1675 ? _258 : _1678;
    assign _1681 = _805 ? _4707 : _1679;
    assign _97 = _1681;
    always @(posedge _791) begin
        if (_789)
            _1678 <= _4707;
        else
            _1678 <= _97;
    end
    assign _1682 = 8'b10011111;
    assign _1683 = _817 == _1682;
    assign _1684 = _814 & _1683;
    assign _1688 = _1684 ? _258 : _1687;
    assign _1690 = _805 ? _4707 : _1688;
    assign _98 = _1690;
    always @(posedge _791) begin
        if (_789)
            _1687 <= _4707;
        else
            _1687 <= _98;
    end
    assign _1691 = 8'b10011110;
    assign _1692 = _817 == _1691;
    assign _1693 = _814 & _1692;
    assign _1697 = _1693 ? _258 : _1696;
    assign _1699 = _805 ? _4707 : _1697;
    assign _99 = _1699;
    always @(posedge _791) begin
        if (_789)
            _1696 <= _4707;
        else
            _1696 <= _99;
    end
    assign _1700 = 8'b10011101;
    assign _1701 = _817 == _1700;
    assign _1702 = _814 & _1701;
    assign _1706 = _1702 ? _258 : _1705;
    assign _1708 = _805 ? _4707 : _1706;
    assign _100 = _1708;
    always @(posedge _791) begin
        if (_789)
            _1705 <= _4707;
        else
            _1705 <= _100;
    end
    assign _1709 = 8'b10011100;
    assign _1710 = _817 == _1709;
    assign _1711 = _814 & _1710;
    assign _1715 = _1711 ? _258 : _1714;
    assign _1717 = _805 ? _4707 : _1715;
    assign _101 = _1717;
    always @(posedge _791) begin
        if (_789)
            _1714 <= _4707;
        else
            _1714 <= _101;
    end
    assign _1718 = 8'b10011011;
    assign _1719 = _817 == _1718;
    assign _1720 = _814 & _1719;
    assign _1724 = _1720 ? _258 : _1723;
    assign _1726 = _805 ? _4707 : _1724;
    assign _102 = _1726;
    always @(posedge _791) begin
        if (_789)
            _1723 <= _4707;
        else
            _1723 <= _102;
    end
    assign _1727 = 8'b10011010;
    assign _1728 = _817 == _1727;
    assign _1729 = _814 & _1728;
    assign _1733 = _1729 ? _258 : _1732;
    assign _1735 = _805 ? _4707 : _1733;
    assign _103 = _1735;
    always @(posedge _791) begin
        if (_789)
            _1732 <= _4707;
        else
            _1732 <= _103;
    end
    assign _1736 = 8'b10011001;
    assign _1737 = _817 == _1736;
    assign _1738 = _814 & _1737;
    assign _1742 = _1738 ? _258 : _1741;
    assign _1744 = _805 ? _4707 : _1742;
    assign _104 = _1744;
    always @(posedge _791) begin
        if (_789)
            _1741 <= _4707;
        else
            _1741 <= _104;
    end
    assign _1745 = 8'b10011000;
    assign _1746 = _817 == _1745;
    assign _1747 = _814 & _1746;
    assign _1751 = _1747 ? _258 : _1750;
    assign _1753 = _805 ? _4707 : _1751;
    assign _105 = _1753;
    always @(posedge _791) begin
        if (_789)
            _1750 <= _4707;
        else
            _1750 <= _105;
    end
    assign _1754 = 8'b10010111;
    assign _1755 = _817 == _1754;
    assign _1756 = _814 & _1755;
    assign _1760 = _1756 ? _258 : _1759;
    assign _1762 = _805 ? _4707 : _1760;
    assign _106 = _1762;
    always @(posedge _791) begin
        if (_789)
            _1759 <= _4707;
        else
            _1759 <= _106;
    end
    assign _1763 = 8'b10010110;
    assign _1764 = _817 == _1763;
    assign _1765 = _814 & _1764;
    assign _1769 = _1765 ? _258 : _1768;
    assign _1771 = _805 ? _4707 : _1769;
    assign _107 = _1771;
    always @(posedge _791) begin
        if (_789)
            _1768 <= _4707;
        else
            _1768 <= _107;
    end
    assign _1772 = 8'b10010101;
    assign _1773 = _817 == _1772;
    assign _1774 = _814 & _1773;
    assign _1778 = _1774 ? _258 : _1777;
    assign _1780 = _805 ? _4707 : _1778;
    assign _108 = _1780;
    always @(posedge _791) begin
        if (_789)
            _1777 <= _4707;
        else
            _1777 <= _108;
    end
    assign _1781 = 8'b10010100;
    assign _1782 = _817 == _1781;
    assign _1783 = _814 & _1782;
    assign _1787 = _1783 ? _258 : _1786;
    assign _1789 = _805 ? _4707 : _1787;
    assign _109 = _1789;
    always @(posedge _791) begin
        if (_789)
            _1786 <= _4707;
        else
            _1786 <= _109;
    end
    assign _1790 = 8'b10010011;
    assign _1791 = _817 == _1790;
    assign _1792 = _814 & _1791;
    assign _1796 = _1792 ? _258 : _1795;
    assign _1798 = _805 ? _4707 : _1796;
    assign _110 = _1798;
    always @(posedge _791) begin
        if (_789)
            _1795 <= _4707;
        else
            _1795 <= _110;
    end
    assign _1799 = 8'b10010010;
    assign _1800 = _817 == _1799;
    assign _1801 = _814 & _1800;
    assign _1805 = _1801 ? _258 : _1804;
    assign _1807 = _805 ? _4707 : _1805;
    assign _111 = _1807;
    always @(posedge _791) begin
        if (_789)
            _1804 <= _4707;
        else
            _1804 <= _111;
    end
    assign _1808 = 8'b10010001;
    assign _1809 = _817 == _1808;
    assign _1810 = _814 & _1809;
    assign _1814 = _1810 ? _258 : _1813;
    assign _1816 = _805 ? _4707 : _1814;
    assign _112 = _1816;
    always @(posedge _791) begin
        if (_789)
            _1813 <= _4707;
        else
            _1813 <= _112;
    end
    assign _1817 = 8'b10010000;
    assign _1818 = _817 == _1817;
    assign _1819 = _814 & _1818;
    assign _1823 = _1819 ? _258 : _1822;
    assign _1825 = _805 ? _4707 : _1823;
    assign _113 = _1825;
    always @(posedge _791) begin
        if (_789)
            _1822 <= _4707;
        else
            _1822 <= _113;
    end
    assign _1826 = 8'b10001111;
    assign _1827 = _817 == _1826;
    assign _1828 = _814 & _1827;
    assign _1832 = _1828 ? _258 : _1831;
    assign _1834 = _805 ? _4707 : _1832;
    assign _114 = _1834;
    always @(posedge _791) begin
        if (_789)
            _1831 <= _4707;
        else
            _1831 <= _114;
    end
    assign _1835 = 8'b10001110;
    assign _1836 = _817 == _1835;
    assign _1837 = _814 & _1836;
    assign _1841 = _1837 ? _258 : _1840;
    assign _1843 = _805 ? _4707 : _1841;
    assign _115 = _1843;
    always @(posedge _791) begin
        if (_789)
            _1840 <= _4707;
        else
            _1840 <= _115;
    end
    assign _1844 = 8'b10001101;
    assign _1845 = _817 == _1844;
    assign _1846 = _814 & _1845;
    assign _1850 = _1846 ? _258 : _1849;
    assign _1852 = _805 ? _4707 : _1850;
    assign _116 = _1852;
    always @(posedge _791) begin
        if (_789)
            _1849 <= _4707;
        else
            _1849 <= _116;
    end
    assign _1853 = 8'b10001100;
    assign _1854 = _817 == _1853;
    assign _1855 = _814 & _1854;
    assign _1859 = _1855 ? _258 : _1858;
    assign _1861 = _805 ? _4707 : _1859;
    assign _117 = _1861;
    always @(posedge _791) begin
        if (_789)
            _1858 <= _4707;
        else
            _1858 <= _117;
    end
    assign _1862 = 8'b10001011;
    assign _1863 = _817 == _1862;
    assign _1864 = _814 & _1863;
    assign _1868 = _1864 ? _258 : _1867;
    assign _1870 = _805 ? _4707 : _1868;
    assign _118 = _1870;
    always @(posedge _791) begin
        if (_789)
            _1867 <= _4707;
        else
            _1867 <= _118;
    end
    assign _1871 = 8'b10001010;
    assign _1872 = _817 == _1871;
    assign _1873 = _814 & _1872;
    assign _1877 = _1873 ? _258 : _1876;
    assign _1879 = _805 ? _4707 : _1877;
    assign _119 = _1879;
    always @(posedge _791) begin
        if (_789)
            _1876 <= _4707;
        else
            _1876 <= _119;
    end
    assign _1880 = 8'b10001001;
    assign _1881 = _817 == _1880;
    assign _1882 = _814 & _1881;
    assign _1886 = _1882 ? _258 : _1885;
    assign _1888 = _805 ? _4707 : _1886;
    assign _120 = _1888;
    always @(posedge _791) begin
        if (_789)
            _1885 <= _4707;
        else
            _1885 <= _120;
    end
    assign _1889 = 8'b10001000;
    assign _1890 = _817 == _1889;
    assign _1891 = _814 & _1890;
    assign _1895 = _1891 ? _258 : _1894;
    assign _1897 = _805 ? _4707 : _1895;
    assign _121 = _1897;
    always @(posedge _791) begin
        if (_789)
            _1894 <= _4707;
        else
            _1894 <= _121;
    end
    assign _1898 = 8'b10000111;
    assign _1899 = _817 == _1898;
    assign _1900 = _814 & _1899;
    assign _1904 = _1900 ? _258 : _1903;
    assign _1906 = _805 ? _4707 : _1904;
    assign _122 = _1906;
    always @(posedge _791) begin
        if (_789)
            _1903 <= _4707;
        else
            _1903 <= _122;
    end
    assign _1907 = 8'b10000110;
    assign _1908 = _817 == _1907;
    assign _1909 = _814 & _1908;
    assign _1913 = _1909 ? _258 : _1912;
    assign _1915 = _805 ? _4707 : _1913;
    assign _123 = _1915;
    always @(posedge _791) begin
        if (_789)
            _1912 <= _4707;
        else
            _1912 <= _123;
    end
    assign _1916 = 8'b10000101;
    assign _1917 = _817 == _1916;
    assign _1918 = _814 & _1917;
    assign _1922 = _1918 ? _258 : _1921;
    assign _1924 = _805 ? _4707 : _1922;
    assign _124 = _1924;
    always @(posedge _791) begin
        if (_789)
            _1921 <= _4707;
        else
            _1921 <= _124;
    end
    assign _1925 = 8'b10000100;
    assign _1926 = _817 == _1925;
    assign _1927 = _814 & _1926;
    assign _1931 = _1927 ? _258 : _1930;
    assign _1933 = _805 ? _4707 : _1931;
    assign _125 = _1933;
    always @(posedge _791) begin
        if (_789)
            _1930 <= _4707;
        else
            _1930 <= _125;
    end
    assign _1934 = 8'b10000011;
    assign _1935 = _817 == _1934;
    assign _1936 = _814 & _1935;
    assign _1940 = _1936 ? _258 : _1939;
    assign _1942 = _805 ? _4707 : _1940;
    assign _126 = _1942;
    always @(posedge _791) begin
        if (_789)
            _1939 <= _4707;
        else
            _1939 <= _126;
    end
    assign _1943 = 8'b10000010;
    assign _1944 = _817 == _1943;
    assign _1945 = _814 & _1944;
    assign _1949 = _1945 ? _258 : _1948;
    assign _1951 = _805 ? _4707 : _1949;
    assign _127 = _1951;
    always @(posedge _791) begin
        if (_789)
            _1948 <= _4707;
        else
            _1948 <= _127;
    end
    assign _1952 = 8'b10000001;
    assign _1953 = _817 == _1952;
    assign _1954 = _814 & _1953;
    assign _1958 = _1954 ? _258 : _1957;
    assign _1960 = _805 ? _4707 : _1958;
    assign _128 = _1960;
    always @(posedge _791) begin
        if (_789)
            _1957 <= _4707;
        else
            _1957 <= _128;
    end
    assign _1961 = 8'b10000000;
    assign _1962 = _817 == _1961;
    assign _1963 = _814 & _1962;
    assign _1967 = _1963 ? _258 : _1966;
    assign _1969 = _805 ? _4707 : _1967;
    assign _129 = _1969;
    always @(posedge _791) begin
        if (_789)
            _1966 <= _4707;
        else
            _1966 <= _129;
    end
    assign _1970 = 8'b01111111;
    assign _1971 = _817 == _1970;
    assign _1972 = _814 & _1971;
    assign _1976 = _1972 ? _258 : _1975;
    assign _1978 = _805 ? _4707 : _1976;
    assign _130 = _1978;
    always @(posedge _791) begin
        if (_789)
            _1975 <= _4707;
        else
            _1975 <= _130;
    end
    assign _1979 = 8'b01111110;
    assign _1980 = _817 == _1979;
    assign _1981 = _814 & _1980;
    assign _1985 = _1981 ? _258 : _1984;
    assign _1987 = _805 ? _4707 : _1985;
    assign _131 = _1987;
    always @(posedge _791) begin
        if (_789)
            _1984 <= _4707;
        else
            _1984 <= _131;
    end
    assign _1988 = 8'b01111101;
    assign _1989 = _817 == _1988;
    assign _1990 = _814 & _1989;
    assign _1994 = _1990 ? _258 : _1993;
    assign _1996 = _805 ? _4707 : _1994;
    assign _132 = _1996;
    always @(posedge _791) begin
        if (_789)
            _1993 <= _4707;
        else
            _1993 <= _132;
    end
    assign _1997 = 8'b01111100;
    assign _1998 = _817 == _1997;
    assign _1999 = _814 & _1998;
    assign _2003 = _1999 ? _258 : _2002;
    assign _2005 = _805 ? _4707 : _2003;
    assign _133 = _2005;
    always @(posedge _791) begin
        if (_789)
            _2002 <= _4707;
        else
            _2002 <= _133;
    end
    assign _2006 = 8'b01111011;
    assign _2007 = _817 == _2006;
    assign _2008 = _814 & _2007;
    assign _2012 = _2008 ? _258 : _2011;
    assign _2014 = _805 ? _4707 : _2012;
    assign _134 = _2014;
    always @(posedge _791) begin
        if (_789)
            _2011 <= _4707;
        else
            _2011 <= _134;
    end
    assign _2015 = 8'b01111010;
    assign _2016 = _817 == _2015;
    assign _2017 = _814 & _2016;
    assign _2021 = _2017 ? _258 : _2020;
    assign _2023 = _805 ? _4707 : _2021;
    assign _135 = _2023;
    always @(posedge _791) begin
        if (_789)
            _2020 <= _4707;
        else
            _2020 <= _135;
    end
    assign _2024 = 8'b01111001;
    assign _2025 = _817 == _2024;
    assign _2026 = _814 & _2025;
    assign _2030 = _2026 ? _258 : _2029;
    assign _2032 = _805 ? _4707 : _2030;
    assign _136 = _2032;
    always @(posedge _791) begin
        if (_789)
            _2029 <= _4707;
        else
            _2029 <= _136;
    end
    assign _2033 = 8'b01111000;
    assign _2034 = _817 == _2033;
    assign _2035 = _814 & _2034;
    assign _2039 = _2035 ? _258 : _2038;
    assign _2041 = _805 ? _4707 : _2039;
    assign _137 = _2041;
    always @(posedge _791) begin
        if (_789)
            _2038 <= _4707;
        else
            _2038 <= _137;
    end
    assign _2042 = 8'b01110111;
    assign _2043 = _817 == _2042;
    assign _2044 = _814 & _2043;
    assign _2048 = _2044 ? _258 : _2047;
    assign _2050 = _805 ? _4707 : _2048;
    assign _138 = _2050;
    always @(posedge _791) begin
        if (_789)
            _2047 <= _4707;
        else
            _2047 <= _138;
    end
    assign _2051 = 8'b01110110;
    assign _2052 = _817 == _2051;
    assign _2053 = _814 & _2052;
    assign _2057 = _2053 ? _258 : _2056;
    assign _2059 = _805 ? _4707 : _2057;
    assign _139 = _2059;
    always @(posedge _791) begin
        if (_789)
            _2056 <= _4707;
        else
            _2056 <= _139;
    end
    assign _2060 = 8'b01110101;
    assign _2061 = _817 == _2060;
    assign _2062 = _814 & _2061;
    assign _2066 = _2062 ? _258 : _2065;
    assign _2068 = _805 ? _4707 : _2066;
    assign _140 = _2068;
    always @(posedge _791) begin
        if (_789)
            _2065 <= _4707;
        else
            _2065 <= _140;
    end
    assign _2069 = 8'b01110100;
    assign _2070 = _817 == _2069;
    assign _2071 = _814 & _2070;
    assign _2075 = _2071 ? _258 : _2074;
    assign _2077 = _805 ? _4707 : _2075;
    assign _141 = _2077;
    always @(posedge _791) begin
        if (_789)
            _2074 <= _4707;
        else
            _2074 <= _141;
    end
    assign _2078 = 8'b01110011;
    assign _2079 = _817 == _2078;
    assign _2080 = _814 & _2079;
    assign _2084 = _2080 ? _258 : _2083;
    assign _2086 = _805 ? _4707 : _2084;
    assign _142 = _2086;
    always @(posedge _791) begin
        if (_789)
            _2083 <= _4707;
        else
            _2083 <= _142;
    end
    assign _2087 = 8'b01110010;
    assign _2088 = _817 == _2087;
    assign _2089 = _814 & _2088;
    assign _2093 = _2089 ? _258 : _2092;
    assign _2095 = _805 ? _4707 : _2093;
    assign _143 = _2095;
    always @(posedge _791) begin
        if (_789)
            _2092 <= _4707;
        else
            _2092 <= _143;
    end
    assign _2096 = 8'b01110001;
    assign _2097 = _817 == _2096;
    assign _2098 = _814 & _2097;
    assign _2102 = _2098 ? _258 : _2101;
    assign _2104 = _805 ? _4707 : _2102;
    assign _144 = _2104;
    always @(posedge _791) begin
        if (_789)
            _2101 <= _4707;
        else
            _2101 <= _144;
    end
    assign _2105 = 8'b01110000;
    assign _2106 = _817 == _2105;
    assign _2107 = _814 & _2106;
    assign _2111 = _2107 ? _258 : _2110;
    assign _2113 = _805 ? _4707 : _2111;
    assign _145 = _2113;
    always @(posedge _791) begin
        if (_789)
            _2110 <= _4707;
        else
            _2110 <= _145;
    end
    assign _2114 = 8'b01101111;
    assign _2115 = _817 == _2114;
    assign _2116 = _814 & _2115;
    assign _2120 = _2116 ? _258 : _2119;
    assign _2122 = _805 ? _4707 : _2120;
    assign _146 = _2122;
    always @(posedge _791) begin
        if (_789)
            _2119 <= _4707;
        else
            _2119 <= _146;
    end
    assign _2123 = 8'b01101110;
    assign _2124 = _817 == _2123;
    assign _2125 = _814 & _2124;
    assign _2129 = _2125 ? _258 : _2128;
    assign _2131 = _805 ? _4707 : _2129;
    assign _147 = _2131;
    always @(posedge _791) begin
        if (_789)
            _2128 <= _4707;
        else
            _2128 <= _147;
    end
    assign _2132 = 8'b01101101;
    assign _2133 = _817 == _2132;
    assign _2134 = _814 & _2133;
    assign _2138 = _2134 ? _258 : _2137;
    assign _2140 = _805 ? _4707 : _2138;
    assign _148 = _2140;
    always @(posedge _791) begin
        if (_789)
            _2137 <= _4707;
        else
            _2137 <= _148;
    end
    assign _2141 = 8'b01101100;
    assign _2142 = _817 == _2141;
    assign _2143 = _814 & _2142;
    assign _2147 = _2143 ? _258 : _2146;
    assign _2149 = _805 ? _4707 : _2147;
    assign _149 = _2149;
    always @(posedge _791) begin
        if (_789)
            _2146 <= _4707;
        else
            _2146 <= _149;
    end
    assign _2150 = 8'b01101011;
    assign _2151 = _817 == _2150;
    assign _2152 = _814 & _2151;
    assign _2156 = _2152 ? _258 : _2155;
    assign _2158 = _805 ? _4707 : _2156;
    assign _150 = _2158;
    always @(posedge _791) begin
        if (_789)
            _2155 <= _4707;
        else
            _2155 <= _150;
    end
    assign _2159 = 8'b01101010;
    assign _2160 = _817 == _2159;
    assign _2161 = _814 & _2160;
    assign _2165 = _2161 ? _258 : _2164;
    assign _2167 = _805 ? _4707 : _2165;
    assign _151 = _2167;
    always @(posedge _791) begin
        if (_789)
            _2164 <= _4707;
        else
            _2164 <= _151;
    end
    assign _2168 = 8'b01101001;
    assign _2169 = _817 == _2168;
    assign _2170 = _814 & _2169;
    assign _2174 = _2170 ? _258 : _2173;
    assign _2176 = _805 ? _4707 : _2174;
    assign _152 = _2176;
    always @(posedge _791) begin
        if (_789)
            _2173 <= _4707;
        else
            _2173 <= _152;
    end
    assign _2177 = 8'b01101000;
    assign _2178 = _817 == _2177;
    assign _2179 = _814 & _2178;
    assign _2183 = _2179 ? _258 : _2182;
    assign _2185 = _805 ? _4707 : _2183;
    assign _153 = _2185;
    always @(posedge _791) begin
        if (_789)
            _2182 <= _4707;
        else
            _2182 <= _153;
    end
    assign _2186 = 8'b01100111;
    assign _2187 = _817 == _2186;
    assign _2188 = _814 & _2187;
    assign _2192 = _2188 ? _258 : _2191;
    assign _2194 = _805 ? _4707 : _2192;
    assign _154 = _2194;
    always @(posedge _791) begin
        if (_789)
            _2191 <= _4707;
        else
            _2191 <= _154;
    end
    assign _2195 = 8'b01100110;
    assign _2196 = _817 == _2195;
    assign _2197 = _814 & _2196;
    assign _2201 = _2197 ? _258 : _2200;
    assign _2203 = _805 ? _4707 : _2201;
    assign _155 = _2203;
    always @(posedge _791) begin
        if (_789)
            _2200 <= _4707;
        else
            _2200 <= _155;
    end
    assign _2204 = 8'b01100101;
    assign _2205 = _817 == _2204;
    assign _2206 = _814 & _2205;
    assign _2210 = _2206 ? _258 : _2209;
    assign _2212 = _805 ? _4707 : _2210;
    assign _156 = _2212;
    always @(posedge _791) begin
        if (_789)
            _2209 <= _4707;
        else
            _2209 <= _156;
    end
    assign _2213 = 8'b01100100;
    assign _2214 = _817 == _2213;
    assign _2215 = _814 & _2214;
    assign _2219 = _2215 ? _258 : _2218;
    assign _2221 = _805 ? _4707 : _2219;
    assign _157 = _2221;
    always @(posedge _791) begin
        if (_789)
            _2218 <= _4707;
        else
            _2218 <= _157;
    end
    assign _2222 = 8'b01100011;
    assign _2223 = _817 == _2222;
    assign _2224 = _814 & _2223;
    assign _2228 = _2224 ? _258 : _2227;
    assign _2230 = _805 ? _4707 : _2228;
    assign _158 = _2230;
    always @(posedge _791) begin
        if (_789)
            _2227 <= _4707;
        else
            _2227 <= _158;
    end
    assign _2231 = 8'b01100010;
    assign _2232 = _817 == _2231;
    assign _2233 = _814 & _2232;
    assign _2237 = _2233 ? _258 : _2236;
    assign _2239 = _805 ? _4707 : _2237;
    assign _159 = _2239;
    always @(posedge _791) begin
        if (_789)
            _2236 <= _4707;
        else
            _2236 <= _159;
    end
    assign _2240 = 8'b01100001;
    assign _2241 = _817 == _2240;
    assign _2242 = _814 & _2241;
    assign _2246 = _2242 ? _258 : _2245;
    assign _2248 = _805 ? _4707 : _2246;
    assign _160 = _2248;
    always @(posedge _791) begin
        if (_789)
            _2245 <= _4707;
        else
            _2245 <= _160;
    end
    assign _2249 = 8'b01100000;
    assign _2250 = _817 == _2249;
    assign _2251 = _814 & _2250;
    assign _2255 = _2251 ? _258 : _2254;
    assign _2257 = _805 ? _4707 : _2255;
    assign _161 = _2257;
    always @(posedge _791) begin
        if (_789)
            _2254 <= _4707;
        else
            _2254 <= _161;
    end
    assign _2258 = 8'b01011111;
    assign _2259 = _817 == _2258;
    assign _2260 = _814 & _2259;
    assign _2264 = _2260 ? _258 : _2263;
    assign _2266 = _805 ? _4707 : _2264;
    assign _162 = _2266;
    always @(posedge _791) begin
        if (_789)
            _2263 <= _4707;
        else
            _2263 <= _162;
    end
    assign _2267 = 8'b01011110;
    assign _2268 = _817 == _2267;
    assign _2269 = _814 & _2268;
    assign _2273 = _2269 ? _258 : _2272;
    assign _2275 = _805 ? _4707 : _2273;
    assign _163 = _2275;
    always @(posedge _791) begin
        if (_789)
            _2272 <= _4707;
        else
            _2272 <= _163;
    end
    assign _2276 = 8'b01011101;
    assign _2277 = _817 == _2276;
    assign _2278 = _814 & _2277;
    assign _2282 = _2278 ? _258 : _2281;
    assign _2284 = _805 ? _4707 : _2282;
    assign _164 = _2284;
    always @(posedge _791) begin
        if (_789)
            _2281 <= _4707;
        else
            _2281 <= _164;
    end
    assign _2285 = 8'b01011100;
    assign _2286 = _817 == _2285;
    assign _2287 = _814 & _2286;
    assign _2291 = _2287 ? _258 : _2290;
    assign _2293 = _805 ? _4707 : _2291;
    assign _165 = _2293;
    always @(posedge _791) begin
        if (_789)
            _2290 <= _4707;
        else
            _2290 <= _165;
    end
    assign _2294 = 8'b01011011;
    assign _2295 = _817 == _2294;
    assign _2296 = _814 & _2295;
    assign _2300 = _2296 ? _258 : _2299;
    assign _2302 = _805 ? _4707 : _2300;
    assign _166 = _2302;
    always @(posedge _791) begin
        if (_789)
            _2299 <= _4707;
        else
            _2299 <= _166;
    end
    assign _2303 = 8'b01011010;
    assign _2304 = _817 == _2303;
    assign _2305 = _814 & _2304;
    assign _2309 = _2305 ? _258 : _2308;
    assign _2311 = _805 ? _4707 : _2309;
    assign _167 = _2311;
    always @(posedge _791) begin
        if (_789)
            _2308 <= _4707;
        else
            _2308 <= _167;
    end
    assign _2312 = 8'b01011001;
    assign _2313 = _817 == _2312;
    assign _2314 = _814 & _2313;
    assign _2318 = _2314 ? _258 : _2317;
    assign _2320 = _805 ? _4707 : _2318;
    assign _168 = _2320;
    always @(posedge _791) begin
        if (_789)
            _2317 <= _4707;
        else
            _2317 <= _168;
    end
    assign _2321 = 8'b01011000;
    assign _2322 = _817 == _2321;
    assign _2323 = _814 & _2322;
    assign _2327 = _2323 ? _258 : _2326;
    assign _2329 = _805 ? _4707 : _2327;
    assign _169 = _2329;
    always @(posedge _791) begin
        if (_789)
            _2326 <= _4707;
        else
            _2326 <= _169;
    end
    assign _2330 = 8'b01010111;
    assign _2331 = _817 == _2330;
    assign _2332 = _814 & _2331;
    assign _2336 = _2332 ? _258 : _2335;
    assign _2338 = _805 ? _4707 : _2336;
    assign _170 = _2338;
    always @(posedge _791) begin
        if (_789)
            _2335 <= _4707;
        else
            _2335 <= _170;
    end
    assign _2339 = 8'b01010110;
    assign _2340 = _817 == _2339;
    assign _2341 = _814 & _2340;
    assign _2345 = _2341 ? _258 : _2344;
    assign _2347 = _805 ? _4707 : _2345;
    assign _171 = _2347;
    always @(posedge _791) begin
        if (_789)
            _2344 <= _4707;
        else
            _2344 <= _171;
    end
    assign _2348 = 8'b01010101;
    assign _2349 = _817 == _2348;
    assign _2350 = _814 & _2349;
    assign _2354 = _2350 ? _258 : _2353;
    assign _2356 = _805 ? _4707 : _2354;
    assign _172 = _2356;
    always @(posedge _791) begin
        if (_789)
            _2353 <= _4707;
        else
            _2353 <= _172;
    end
    assign _2357 = 8'b01010100;
    assign _2358 = _817 == _2357;
    assign _2359 = _814 & _2358;
    assign _2363 = _2359 ? _258 : _2362;
    assign _2365 = _805 ? _4707 : _2363;
    assign _173 = _2365;
    always @(posedge _791) begin
        if (_789)
            _2362 <= _4707;
        else
            _2362 <= _173;
    end
    assign _2366 = 8'b01010011;
    assign _2367 = _817 == _2366;
    assign _2368 = _814 & _2367;
    assign _2372 = _2368 ? _258 : _2371;
    assign _2374 = _805 ? _4707 : _2372;
    assign _174 = _2374;
    always @(posedge _791) begin
        if (_789)
            _2371 <= _4707;
        else
            _2371 <= _174;
    end
    assign _2375 = 8'b01010010;
    assign _2376 = _817 == _2375;
    assign _2377 = _814 & _2376;
    assign _2381 = _2377 ? _258 : _2380;
    assign _2383 = _805 ? _4707 : _2381;
    assign _175 = _2383;
    always @(posedge _791) begin
        if (_789)
            _2380 <= _4707;
        else
            _2380 <= _175;
    end
    assign _2384 = 8'b01010001;
    assign _2385 = _817 == _2384;
    assign _2386 = _814 & _2385;
    assign _2390 = _2386 ? _258 : _2389;
    assign _2392 = _805 ? _4707 : _2390;
    assign _176 = _2392;
    always @(posedge _791) begin
        if (_789)
            _2389 <= _4707;
        else
            _2389 <= _176;
    end
    assign _2393 = 8'b01010000;
    assign _2394 = _817 == _2393;
    assign _2395 = _814 & _2394;
    assign _2399 = _2395 ? _258 : _2398;
    assign _2401 = _805 ? _4707 : _2399;
    assign _177 = _2401;
    always @(posedge _791) begin
        if (_789)
            _2398 <= _4707;
        else
            _2398 <= _177;
    end
    assign _2402 = 8'b01001111;
    assign _2403 = _817 == _2402;
    assign _2404 = _814 & _2403;
    assign _2408 = _2404 ? _258 : _2407;
    assign _2410 = _805 ? _4707 : _2408;
    assign _178 = _2410;
    always @(posedge _791) begin
        if (_789)
            _2407 <= _4707;
        else
            _2407 <= _178;
    end
    assign _2411 = 8'b01001110;
    assign _2412 = _817 == _2411;
    assign _2413 = _814 & _2412;
    assign _2417 = _2413 ? _258 : _2416;
    assign _2419 = _805 ? _4707 : _2417;
    assign _179 = _2419;
    always @(posedge _791) begin
        if (_789)
            _2416 <= _4707;
        else
            _2416 <= _179;
    end
    assign _2420 = 8'b01001101;
    assign _2421 = _817 == _2420;
    assign _2422 = _814 & _2421;
    assign _2426 = _2422 ? _258 : _2425;
    assign _2428 = _805 ? _4707 : _2426;
    assign _180 = _2428;
    always @(posedge _791) begin
        if (_789)
            _2425 <= _4707;
        else
            _2425 <= _180;
    end
    assign _2429 = 8'b01001100;
    assign _2430 = _817 == _2429;
    assign _2431 = _814 & _2430;
    assign _2435 = _2431 ? _258 : _2434;
    assign _2437 = _805 ? _4707 : _2435;
    assign _181 = _2437;
    always @(posedge _791) begin
        if (_789)
            _2434 <= _4707;
        else
            _2434 <= _181;
    end
    assign _2438 = 8'b01001011;
    assign _2439 = _817 == _2438;
    assign _2440 = _814 & _2439;
    assign _2444 = _2440 ? _258 : _2443;
    assign _2446 = _805 ? _4707 : _2444;
    assign _182 = _2446;
    always @(posedge _791) begin
        if (_789)
            _2443 <= _4707;
        else
            _2443 <= _182;
    end
    assign _2447 = 8'b01001010;
    assign _2448 = _817 == _2447;
    assign _2449 = _814 & _2448;
    assign _2453 = _2449 ? _258 : _2452;
    assign _2455 = _805 ? _4707 : _2453;
    assign _183 = _2455;
    always @(posedge _791) begin
        if (_789)
            _2452 <= _4707;
        else
            _2452 <= _183;
    end
    assign _2456 = 8'b01001001;
    assign _2457 = _817 == _2456;
    assign _2458 = _814 & _2457;
    assign _2462 = _2458 ? _258 : _2461;
    assign _2464 = _805 ? _4707 : _2462;
    assign _184 = _2464;
    always @(posedge _791) begin
        if (_789)
            _2461 <= _4707;
        else
            _2461 <= _184;
    end
    assign _2465 = 8'b01001000;
    assign _2466 = _817 == _2465;
    assign _2467 = _814 & _2466;
    assign _2471 = _2467 ? _258 : _2470;
    assign _2473 = _805 ? _4707 : _2471;
    assign _185 = _2473;
    always @(posedge _791) begin
        if (_789)
            _2470 <= _4707;
        else
            _2470 <= _185;
    end
    assign _2474 = 8'b01000111;
    assign _2475 = _817 == _2474;
    assign _2476 = _814 & _2475;
    assign _2480 = _2476 ? _258 : _2479;
    assign _2482 = _805 ? _4707 : _2480;
    assign _186 = _2482;
    always @(posedge _791) begin
        if (_789)
            _2479 <= _4707;
        else
            _2479 <= _186;
    end
    assign _2483 = 8'b01000110;
    assign _2484 = _817 == _2483;
    assign _2485 = _814 & _2484;
    assign _2489 = _2485 ? _258 : _2488;
    assign _2491 = _805 ? _4707 : _2489;
    assign _187 = _2491;
    always @(posedge _791) begin
        if (_789)
            _2488 <= _4707;
        else
            _2488 <= _187;
    end
    assign _2492 = 8'b01000101;
    assign _2493 = _817 == _2492;
    assign _2494 = _814 & _2493;
    assign _2498 = _2494 ? _258 : _2497;
    assign _2500 = _805 ? _4707 : _2498;
    assign _188 = _2500;
    always @(posedge _791) begin
        if (_789)
            _2497 <= _4707;
        else
            _2497 <= _188;
    end
    assign _2501 = 8'b01000100;
    assign _2502 = _817 == _2501;
    assign _2503 = _814 & _2502;
    assign _2507 = _2503 ? _258 : _2506;
    assign _2509 = _805 ? _4707 : _2507;
    assign _189 = _2509;
    always @(posedge _791) begin
        if (_789)
            _2506 <= _4707;
        else
            _2506 <= _189;
    end
    assign _2510 = 8'b01000011;
    assign _2511 = _817 == _2510;
    assign _2512 = _814 & _2511;
    assign _2516 = _2512 ? _258 : _2515;
    assign _2518 = _805 ? _4707 : _2516;
    assign _190 = _2518;
    always @(posedge _791) begin
        if (_789)
            _2515 <= _4707;
        else
            _2515 <= _190;
    end
    assign _2519 = 8'b01000010;
    assign _2520 = _817 == _2519;
    assign _2521 = _814 & _2520;
    assign _2525 = _2521 ? _258 : _2524;
    assign _2527 = _805 ? _4707 : _2525;
    assign _191 = _2527;
    always @(posedge _791) begin
        if (_789)
            _2524 <= _4707;
        else
            _2524 <= _191;
    end
    assign _2528 = 8'b01000001;
    assign _2529 = _817 == _2528;
    assign _2530 = _814 & _2529;
    assign _2534 = _2530 ? _258 : _2533;
    assign _2536 = _805 ? _4707 : _2534;
    assign _192 = _2536;
    always @(posedge _791) begin
        if (_789)
            _2533 <= _4707;
        else
            _2533 <= _192;
    end
    assign _2537 = 8'b01000000;
    assign _2538 = _817 == _2537;
    assign _2539 = _814 & _2538;
    assign _2543 = _2539 ? _258 : _2542;
    assign _2545 = _805 ? _4707 : _2543;
    assign _193 = _2545;
    always @(posedge _791) begin
        if (_789)
            _2542 <= _4707;
        else
            _2542 <= _193;
    end
    assign _2546 = 8'b00111111;
    assign _2547 = _817 == _2546;
    assign _2548 = _814 & _2547;
    assign _2552 = _2548 ? _258 : _2551;
    assign _2554 = _805 ? _4707 : _2552;
    assign _194 = _2554;
    always @(posedge _791) begin
        if (_789)
            _2551 <= _4707;
        else
            _2551 <= _194;
    end
    assign _2555 = 8'b00111110;
    assign _2556 = _817 == _2555;
    assign _2557 = _814 & _2556;
    assign _2561 = _2557 ? _258 : _2560;
    assign _2563 = _805 ? _4707 : _2561;
    assign _195 = _2563;
    always @(posedge _791) begin
        if (_789)
            _2560 <= _4707;
        else
            _2560 <= _195;
    end
    assign _2564 = 8'b00111101;
    assign _2565 = _817 == _2564;
    assign _2566 = _814 & _2565;
    assign _2570 = _2566 ? _258 : _2569;
    assign _2572 = _805 ? _4707 : _2570;
    assign _196 = _2572;
    always @(posedge _791) begin
        if (_789)
            _2569 <= _4707;
        else
            _2569 <= _196;
    end
    assign _2573 = 8'b00111100;
    assign _2574 = _817 == _2573;
    assign _2575 = _814 & _2574;
    assign _2579 = _2575 ? _258 : _2578;
    assign _2581 = _805 ? _4707 : _2579;
    assign _197 = _2581;
    always @(posedge _791) begin
        if (_789)
            _2578 <= _4707;
        else
            _2578 <= _197;
    end
    assign _2582 = 8'b00111011;
    assign _2583 = _817 == _2582;
    assign _2584 = _814 & _2583;
    assign _2588 = _2584 ? _258 : _2587;
    assign _2590 = _805 ? _4707 : _2588;
    assign _198 = _2590;
    always @(posedge _791) begin
        if (_789)
            _2587 <= _4707;
        else
            _2587 <= _198;
    end
    assign _2591 = 8'b00111010;
    assign _2592 = _817 == _2591;
    assign _2593 = _814 & _2592;
    assign _2597 = _2593 ? _258 : _2596;
    assign _2599 = _805 ? _4707 : _2597;
    assign _199 = _2599;
    always @(posedge _791) begin
        if (_789)
            _2596 <= _4707;
        else
            _2596 <= _199;
    end
    assign _2600 = 8'b00111001;
    assign _2601 = _817 == _2600;
    assign _2602 = _814 & _2601;
    assign _2606 = _2602 ? _258 : _2605;
    assign _2608 = _805 ? _4707 : _2606;
    assign _200 = _2608;
    always @(posedge _791) begin
        if (_789)
            _2605 <= _4707;
        else
            _2605 <= _200;
    end
    assign _2609 = 8'b00111000;
    assign _2610 = _817 == _2609;
    assign _2611 = _814 & _2610;
    assign _2615 = _2611 ? _258 : _2614;
    assign _2617 = _805 ? _4707 : _2615;
    assign _201 = _2617;
    always @(posedge _791) begin
        if (_789)
            _2614 <= _4707;
        else
            _2614 <= _201;
    end
    assign _2618 = 8'b00110111;
    assign _2619 = _817 == _2618;
    assign _2620 = _814 & _2619;
    assign _2624 = _2620 ? _258 : _2623;
    assign _2626 = _805 ? _4707 : _2624;
    assign _202 = _2626;
    always @(posedge _791) begin
        if (_789)
            _2623 <= _4707;
        else
            _2623 <= _202;
    end
    assign _2627 = 8'b00110110;
    assign _2628 = _817 == _2627;
    assign _2629 = _814 & _2628;
    assign _2633 = _2629 ? _258 : _2632;
    assign _2635 = _805 ? _4707 : _2633;
    assign _203 = _2635;
    always @(posedge _791) begin
        if (_789)
            _2632 <= _4707;
        else
            _2632 <= _203;
    end
    assign _2636 = 8'b00110101;
    assign _2637 = _817 == _2636;
    assign _2638 = _814 & _2637;
    assign _2642 = _2638 ? _258 : _2641;
    assign _2644 = _805 ? _4707 : _2642;
    assign _204 = _2644;
    always @(posedge _791) begin
        if (_789)
            _2641 <= _4707;
        else
            _2641 <= _204;
    end
    assign _2645 = 8'b00110100;
    assign _2646 = _817 == _2645;
    assign _2647 = _814 & _2646;
    assign _2651 = _2647 ? _258 : _2650;
    assign _2653 = _805 ? _4707 : _2651;
    assign _205 = _2653;
    always @(posedge _791) begin
        if (_789)
            _2650 <= _4707;
        else
            _2650 <= _205;
    end
    assign _2654 = 8'b00110011;
    assign _2655 = _817 == _2654;
    assign _2656 = _814 & _2655;
    assign _2660 = _2656 ? _258 : _2659;
    assign _2662 = _805 ? _4707 : _2660;
    assign _206 = _2662;
    always @(posedge _791) begin
        if (_789)
            _2659 <= _4707;
        else
            _2659 <= _206;
    end
    assign _2663 = 8'b00110010;
    assign _2664 = _817 == _2663;
    assign _2665 = _814 & _2664;
    assign _2669 = _2665 ? _258 : _2668;
    assign _2671 = _805 ? _4707 : _2669;
    assign _207 = _2671;
    always @(posedge _791) begin
        if (_789)
            _2668 <= _4707;
        else
            _2668 <= _207;
    end
    assign _2672 = 8'b00110001;
    assign _2673 = _817 == _2672;
    assign _2674 = _814 & _2673;
    assign _2678 = _2674 ? _258 : _2677;
    assign _2680 = _805 ? _4707 : _2678;
    assign _208 = _2680;
    always @(posedge _791) begin
        if (_789)
            _2677 <= _4707;
        else
            _2677 <= _208;
    end
    assign _2681 = 8'b00110000;
    assign _2682 = _817 == _2681;
    assign _2683 = _814 & _2682;
    assign _2687 = _2683 ? _258 : _2686;
    assign _2689 = _805 ? _4707 : _2687;
    assign _209 = _2689;
    always @(posedge _791) begin
        if (_789)
            _2686 <= _4707;
        else
            _2686 <= _209;
    end
    assign _2690 = 8'b00101111;
    assign _2691 = _817 == _2690;
    assign _2692 = _814 & _2691;
    assign _2696 = _2692 ? _258 : _2695;
    assign _2698 = _805 ? _4707 : _2696;
    assign _210 = _2698;
    always @(posedge _791) begin
        if (_789)
            _2695 <= _4707;
        else
            _2695 <= _210;
    end
    assign _2699 = 8'b00101110;
    assign _2700 = _817 == _2699;
    assign _2701 = _814 & _2700;
    assign _2705 = _2701 ? _258 : _2704;
    assign _2707 = _805 ? _4707 : _2705;
    assign _211 = _2707;
    always @(posedge _791) begin
        if (_789)
            _2704 <= _4707;
        else
            _2704 <= _211;
    end
    assign _2708 = 8'b00101101;
    assign _2709 = _817 == _2708;
    assign _2710 = _814 & _2709;
    assign _2714 = _2710 ? _258 : _2713;
    assign _2716 = _805 ? _4707 : _2714;
    assign _212 = _2716;
    always @(posedge _791) begin
        if (_789)
            _2713 <= _4707;
        else
            _2713 <= _212;
    end
    assign _2717 = 8'b00101100;
    assign _2718 = _817 == _2717;
    assign _2719 = _814 & _2718;
    assign _2723 = _2719 ? _258 : _2722;
    assign _2725 = _805 ? _4707 : _2723;
    assign _213 = _2725;
    always @(posedge _791) begin
        if (_789)
            _2722 <= _4707;
        else
            _2722 <= _213;
    end
    assign _2726 = 8'b00101011;
    assign _2727 = _817 == _2726;
    assign _2728 = _814 & _2727;
    assign _2732 = _2728 ? _258 : _2731;
    assign _2734 = _805 ? _4707 : _2732;
    assign _214 = _2734;
    always @(posedge _791) begin
        if (_789)
            _2731 <= _4707;
        else
            _2731 <= _214;
    end
    assign _2735 = 8'b00101010;
    assign _2736 = _817 == _2735;
    assign _2737 = _814 & _2736;
    assign _2741 = _2737 ? _258 : _2740;
    assign _2743 = _805 ? _4707 : _2741;
    assign _215 = _2743;
    always @(posedge _791) begin
        if (_789)
            _2740 <= _4707;
        else
            _2740 <= _215;
    end
    assign _2744 = 8'b00101001;
    assign _2745 = _817 == _2744;
    assign _2746 = _814 & _2745;
    assign _2750 = _2746 ? _258 : _2749;
    assign _2752 = _805 ? _4707 : _2750;
    assign _216 = _2752;
    always @(posedge _791) begin
        if (_789)
            _2749 <= _4707;
        else
            _2749 <= _216;
    end
    assign _2753 = 8'b00101000;
    assign _2754 = _817 == _2753;
    assign _2755 = _814 & _2754;
    assign _2759 = _2755 ? _258 : _2758;
    assign _2761 = _805 ? _4707 : _2759;
    assign _217 = _2761;
    always @(posedge _791) begin
        if (_789)
            _2758 <= _4707;
        else
            _2758 <= _217;
    end
    assign _2762 = 8'b00100111;
    assign _2763 = _817 == _2762;
    assign _2764 = _814 & _2763;
    assign _2768 = _2764 ? _258 : _2767;
    assign _2770 = _805 ? _4707 : _2768;
    assign _218 = _2770;
    always @(posedge _791) begin
        if (_789)
            _2767 <= _4707;
        else
            _2767 <= _218;
    end
    assign _2771 = 8'b00100110;
    assign _2772 = _817 == _2771;
    assign _2773 = _814 & _2772;
    assign _2777 = _2773 ? _258 : _2776;
    assign _2779 = _805 ? _4707 : _2777;
    assign _219 = _2779;
    always @(posedge _791) begin
        if (_789)
            _2776 <= _4707;
        else
            _2776 <= _219;
    end
    assign _2780 = 8'b00100101;
    assign _2781 = _817 == _2780;
    assign _2782 = _814 & _2781;
    assign _2786 = _2782 ? _258 : _2785;
    assign _2788 = _805 ? _4707 : _2786;
    assign _220 = _2788;
    always @(posedge _791) begin
        if (_789)
            _2785 <= _4707;
        else
            _2785 <= _220;
    end
    assign _2789 = 8'b00100100;
    assign _2790 = _817 == _2789;
    assign _2791 = _814 & _2790;
    assign _2795 = _2791 ? _258 : _2794;
    assign _2797 = _805 ? _4707 : _2795;
    assign _221 = _2797;
    always @(posedge _791) begin
        if (_789)
            _2794 <= _4707;
        else
            _2794 <= _221;
    end
    assign _2798 = 8'b00100011;
    assign _2799 = _817 == _2798;
    assign _2800 = _814 & _2799;
    assign _2804 = _2800 ? _258 : _2803;
    assign _2806 = _805 ? _4707 : _2804;
    assign _222 = _2806;
    always @(posedge _791) begin
        if (_789)
            _2803 <= _4707;
        else
            _2803 <= _222;
    end
    assign _2807 = 8'b00100010;
    assign _2808 = _817 == _2807;
    assign _2809 = _814 & _2808;
    assign _2813 = _2809 ? _258 : _2812;
    assign _2815 = _805 ? _4707 : _2813;
    assign _223 = _2815;
    always @(posedge _791) begin
        if (_789)
            _2812 <= _4707;
        else
            _2812 <= _223;
    end
    assign _2816 = 8'b00100001;
    assign _2817 = _817 == _2816;
    assign _2818 = _814 & _2817;
    assign _2822 = _2818 ? _258 : _2821;
    assign _2824 = _805 ? _4707 : _2822;
    assign _224 = _2824;
    always @(posedge _791) begin
        if (_789)
            _2821 <= _4707;
        else
            _2821 <= _224;
    end
    assign _2825 = 8'b00100000;
    assign _2826 = _817 == _2825;
    assign _2827 = _814 & _2826;
    assign _2831 = _2827 ? _258 : _2830;
    assign _2833 = _805 ? _4707 : _2831;
    assign _225 = _2833;
    always @(posedge _791) begin
        if (_789)
            _2830 <= _4707;
        else
            _2830 <= _225;
    end
    assign _2834 = 8'b00011111;
    assign _2835 = _817 == _2834;
    assign _2836 = _814 & _2835;
    assign _2840 = _2836 ? _258 : _2839;
    assign _2842 = _805 ? _4707 : _2840;
    assign _226 = _2842;
    always @(posedge _791) begin
        if (_789)
            _2839 <= _4707;
        else
            _2839 <= _226;
    end
    assign _2843 = 8'b00011110;
    assign _2844 = _817 == _2843;
    assign _2845 = _814 & _2844;
    assign _2849 = _2845 ? _258 : _2848;
    assign _2851 = _805 ? _4707 : _2849;
    assign _227 = _2851;
    always @(posedge _791) begin
        if (_789)
            _2848 <= _4707;
        else
            _2848 <= _227;
    end
    assign _2852 = 8'b00011101;
    assign _2853 = _817 == _2852;
    assign _2854 = _814 & _2853;
    assign _2858 = _2854 ? _258 : _2857;
    assign _2860 = _805 ? _4707 : _2858;
    assign _228 = _2860;
    always @(posedge _791) begin
        if (_789)
            _2857 <= _4707;
        else
            _2857 <= _228;
    end
    assign _2861 = 8'b00011100;
    assign _2862 = _817 == _2861;
    assign _2863 = _814 & _2862;
    assign _2867 = _2863 ? _258 : _2866;
    assign _2869 = _805 ? _4707 : _2867;
    assign _229 = _2869;
    always @(posedge _791) begin
        if (_789)
            _2866 <= _4707;
        else
            _2866 <= _229;
    end
    assign _2870 = 8'b00011011;
    assign _2871 = _817 == _2870;
    assign _2872 = _814 & _2871;
    assign _2876 = _2872 ? _258 : _2875;
    assign _2878 = _805 ? _4707 : _2876;
    assign _230 = _2878;
    always @(posedge _791) begin
        if (_789)
            _2875 <= _4707;
        else
            _2875 <= _230;
    end
    assign _2879 = 8'b00011010;
    assign _2880 = _817 == _2879;
    assign _2881 = _814 & _2880;
    assign _2885 = _2881 ? _258 : _2884;
    assign _2887 = _805 ? _4707 : _2885;
    assign _231 = _2887;
    always @(posedge _791) begin
        if (_789)
            _2884 <= _4707;
        else
            _2884 <= _231;
    end
    assign _2888 = 8'b00011001;
    assign _2889 = _817 == _2888;
    assign _2890 = _814 & _2889;
    assign _2894 = _2890 ? _258 : _2893;
    assign _2896 = _805 ? _4707 : _2894;
    assign _232 = _2896;
    always @(posedge _791) begin
        if (_789)
            _2893 <= _4707;
        else
            _2893 <= _232;
    end
    assign _2897 = 8'b00011000;
    assign _2898 = _817 == _2897;
    assign _2899 = _814 & _2898;
    assign _2903 = _2899 ? _258 : _2902;
    assign _2905 = _805 ? _4707 : _2903;
    assign _233 = _2905;
    always @(posedge _791) begin
        if (_789)
            _2902 <= _4707;
        else
            _2902 <= _233;
    end
    assign _2906 = 8'b00010111;
    assign _2907 = _817 == _2906;
    assign _2908 = _814 & _2907;
    assign _2912 = _2908 ? _258 : _2911;
    assign _2914 = _805 ? _4707 : _2912;
    assign _234 = _2914;
    always @(posedge _791) begin
        if (_789)
            _2911 <= _4707;
        else
            _2911 <= _234;
    end
    assign _2915 = 8'b00010110;
    assign _2916 = _817 == _2915;
    assign _2917 = _814 & _2916;
    assign _2921 = _2917 ? _258 : _2920;
    assign _2923 = _805 ? _4707 : _2921;
    assign _235 = _2923;
    always @(posedge _791) begin
        if (_789)
            _2920 <= _4707;
        else
            _2920 <= _235;
    end
    assign _2924 = 8'b00010101;
    assign _2925 = _817 == _2924;
    assign _2926 = _814 & _2925;
    assign _2930 = _2926 ? _258 : _2929;
    assign _2932 = _805 ? _4707 : _2930;
    assign _236 = _2932;
    always @(posedge _791) begin
        if (_789)
            _2929 <= _4707;
        else
            _2929 <= _236;
    end
    assign _2933 = 8'b00010100;
    assign _2934 = _817 == _2933;
    assign _2935 = _814 & _2934;
    assign _2939 = _2935 ? _258 : _2938;
    assign _2941 = _805 ? _4707 : _2939;
    assign _237 = _2941;
    always @(posedge _791) begin
        if (_789)
            _2938 <= _4707;
        else
            _2938 <= _237;
    end
    assign _2942 = 8'b00010011;
    assign _2943 = _817 == _2942;
    assign _2944 = _814 & _2943;
    assign _2948 = _2944 ? _258 : _2947;
    assign _2950 = _805 ? _4707 : _2948;
    assign _238 = _2950;
    always @(posedge _791) begin
        if (_789)
            _2947 <= _4707;
        else
            _2947 <= _238;
    end
    assign _2951 = 8'b00010010;
    assign _2952 = _817 == _2951;
    assign _2953 = _814 & _2952;
    assign _2957 = _2953 ? _258 : _2956;
    assign _2959 = _805 ? _4707 : _2957;
    assign _239 = _2959;
    always @(posedge _791) begin
        if (_789)
            _2956 <= _4707;
        else
            _2956 <= _239;
    end
    assign _2960 = 8'b00010001;
    assign _2961 = _817 == _2960;
    assign _2962 = _814 & _2961;
    assign _2966 = _2962 ? _258 : _2965;
    assign _2968 = _805 ? _4707 : _2966;
    assign _240 = _2968;
    always @(posedge _791) begin
        if (_789)
            _2965 <= _4707;
        else
            _2965 <= _240;
    end
    assign _2969 = 8'b00010000;
    assign _2970 = _817 == _2969;
    assign _2971 = _814 & _2970;
    assign _2975 = _2971 ? _258 : _2974;
    assign _2977 = _805 ? _4707 : _2975;
    assign _241 = _2977;
    always @(posedge _791) begin
        if (_789)
            _2974 <= _4707;
        else
            _2974 <= _241;
    end
    assign _2978 = 8'b00001111;
    assign _2979 = _817 == _2978;
    assign _2980 = _814 & _2979;
    assign _2984 = _2980 ? _258 : _2983;
    assign _2986 = _805 ? _4707 : _2984;
    assign _242 = _2986;
    always @(posedge _791) begin
        if (_789)
            _2983 <= _4707;
        else
            _2983 <= _242;
    end
    assign _2987 = 8'b00001110;
    assign _2988 = _817 == _2987;
    assign _2989 = _814 & _2988;
    assign _2993 = _2989 ? _258 : _2992;
    assign _2995 = _805 ? _4707 : _2993;
    assign _243 = _2995;
    always @(posedge _791) begin
        if (_789)
            _2992 <= _4707;
        else
            _2992 <= _243;
    end
    assign _2996 = 8'b00001101;
    assign _2997 = _817 == _2996;
    assign _2998 = _814 & _2997;
    assign _3002 = _2998 ? _258 : _3001;
    assign _3004 = _805 ? _4707 : _3002;
    assign _244 = _3004;
    always @(posedge _791) begin
        if (_789)
            _3001 <= _4707;
        else
            _3001 <= _244;
    end
    assign _3005 = 8'b00001100;
    assign _3006 = _817 == _3005;
    assign _3007 = _814 & _3006;
    assign _3011 = _3007 ? _258 : _3010;
    assign _3013 = _805 ? _4707 : _3011;
    assign _245 = _3013;
    always @(posedge _791) begin
        if (_789)
            _3010 <= _4707;
        else
            _3010 <= _245;
    end
    assign _3014 = 8'b00001011;
    assign _3015 = _817 == _3014;
    assign _3016 = _814 & _3015;
    assign _3020 = _3016 ? _258 : _3019;
    assign _3022 = _805 ? _4707 : _3020;
    assign _246 = _3022;
    always @(posedge _791) begin
        if (_789)
            _3019 <= _4707;
        else
            _3019 <= _246;
    end
    assign _3023 = 8'b00001010;
    assign _3024 = _817 == _3023;
    assign _3025 = _814 & _3024;
    assign _3029 = _3025 ? _258 : _3028;
    assign _3031 = _805 ? _4707 : _3029;
    assign _247 = _3031;
    always @(posedge _791) begin
        if (_789)
            _3028 <= _4707;
        else
            _3028 <= _247;
    end
    assign _3032 = 8'b00001001;
    assign _3033 = _817 == _3032;
    assign _3034 = _814 & _3033;
    assign _3038 = _3034 ? _258 : _3037;
    assign _3040 = _805 ? _4707 : _3038;
    assign _248 = _3040;
    always @(posedge _791) begin
        if (_789)
            _3037 <= _4707;
        else
            _3037 <= _248;
    end
    assign _3041 = 8'b00001000;
    assign _3042 = _817 == _3041;
    assign _3043 = _814 & _3042;
    assign _3047 = _3043 ? _258 : _3046;
    assign _3049 = _805 ? _4707 : _3047;
    assign _249 = _3049;
    always @(posedge _791) begin
        if (_789)
            _3046 <= _4707;
        else
            _3046 <= _249;
    end
    assign _3050 = 8'b00000111;
    assign _3051 = _817 == _3050;
    assign _3052 = _814 & _3051;
    assign _3056 = _3052 ? _258 : _3055;
    assign _3058 = _805 ? _4707 : _3056;
    assign _250 = _3058;
    always @(posedge _791) begin
        if (_789)
            _3055 <= _4707;
        else
            _3055 <= _250;
    end
    assign _3059 = 8'b00000110;
    assign _3060 = _817 == _3059;
    assign _3061 = _814 & _3060;
    assign _3065 = _3061 ? _258 : _3064;
    assign _3067 = _805 ? _4707 : _3065;
    assign _251 = _3067;
    always @(posedge _791) begin
        if (_789)
            _3064 <= _4707;
        else
            _3064 <= _251;
    end
    assign _3068 = 8'b00000101;
    assign _3069 = _817 == _3068;
    assign _3070 = _814 & _3069;
    assign _3074 = _3070 ? _258 : _3073;
    assign _3076 = _805 ? _4707 : _3074;
    assign _252 = _3076;
    always @(posedge _791) begin
        if (_789)
            _3073 <= _4707;
        else
            _3073 <= _252;
    end
    assign _3077 = 8'b00000100;
    assign _3078 = _817 == _3077;
    assign _3079 = _814 & _3078;
    assign _3083 = _3079 ? _258 : _3082;
    assign _3085 = _805 ? _4707 : _3083;
    assign _253 = _3085;
    always @(posedge _791) begin
        if (_789)
            _3082 <= _4707;
        else
            _3082 <= _253;
    end
    assign _3086 = 8'b00000011;
    assign _3087 = _817 == _3086;
    assign _3088 = _814 & _3087;
    assign _3092 = _3088 ? _258 : _3091;
    assign _3094 = _805 ? _4707 : _3092;
    assign _254 = _3094;
    always @(posedge _791) begin
        if (_789)
            _3091 <= _4707;
        else
            _3091 <= _254;
    end
    assign _3095 = 8'b00000010;
    assign _3096 = _817 == _3095;
    assign _3097 = _814 & _3096;
    assign _3101 = _3097 ? _258 : _3100;
    assign _3103 = _805 ? _4707 : _3101;
    assign _255 = _3103;
    always @(posedge _791) begin
        if (_789)
            _3100 <= _4707;
        else
            _3100 <= _255;
    end
    assign _3104 = 8'b00000001;
    assign _3105 = _817 == _3104;
    assign _3106 = _814 & _3105;
    assign _3110 = _3106 ? _258 : _3109;
    assign _3112 = _805 ? _4707 : _3110;
    assign _256 = _3112;
    always @(posedge _791) begin
        if (_789)
            _3109 <= _4707;
        else
            _3109 <= _256;
    end
    assign _258 = x0_value;
    assign _3118 = 8'b00000000;
    assign _3116 = _3114 + _3104;
    assign _3114 = _805 ? _3118 : _817;
    assign _3117 = _814 ? _3116 : _3114;
    assign _259 = _3117;
    always @(posedge _791) begin
        if (_789)
            _817 <= _3118;
        else
            _817 <= _259;
    end
    assign _3119 = _817 == _3118;
    assign _3120 = _814 & _3119;
    assign _3124 = _3120 ? _258 : _3123;
    assign _3126 = _805 ? _4707 : _3124;
    assign _260 = _3126;
    always @(posedge _791) begin
        if (_789)
            _3123 <= _4707;
        else
            _3123 <= _260;
    end
    always @* begin
        case (_785)
        0:
            _4705 <= _3123;
        1:
            _4705 <= _3109;
        2:
            _4705 <= _3100;
        3:
            _4705 <= _3091;
        4:
            _4705 <= _3082;
        5:
            _4705 <= _3073;
        6:
            _4705 <= _3064;
        7:
            _4705 <= _3055;
        8:
            _4705 <= _3046;
        9:
            _4705 <= _3037;
        10:
            _4705 <= _3028;
        11:
            _4705 <= _3019;
        12:
            _4705 <= _3010;
        13:
            _4705 <= _3001;
        14:
            _4705 <= _2992;
        15:
            _4705 <= _2983;
        16:
            _4705 <= _2974;
        17:
            _4705 <= _2965;
        18:
            _4705 <= _2956;
        19:
            _4705 <= _2947;
        20:
            _4705 <= _2938;
        21:
            _4705 <= _2929;
        22:
            _4705 <= _2920;
        23:
            _4705 <= _2911;
        24:
            _4705 <= _2902;
        25:
            _4705 <= _2893;
        26:
            _4705 <= _2884;
        27:
            _4705 <= _2875;
        28:
            _4705 <= _2866;
        29:
            _4705 <= _2857;
        30:
            _4705 <= _2848;
        31:
            _4705 <= _2839;
        32:
            _4705 <= _2830;
        33:
            _4705 <= _2821;
        34:
            _4705 <= _2812;
        35:
            _4705 <= _2803;
        36:
            _4705 <= _2794;
        37:
            _4705 <= _2785;
        38:
            _4705 <= _2776;
        39:
            _4705 <= _2767;
        40:
            _4705 <= _2758;
        41:
            _4705 <= _2749;
        42:
            _4705 <= _2740;
        43:
            _4705 <= _2731;
        44:
            _4705 <= _2722;
        45:
            _4705 <= _2713;
        46:
            _4705 <= _2704;
        47:
            _4705 <= _2695;
        48:
            _4705 <= _2686;
        49:
            _4705 <= _2677;
        50:
            _4705 <= _2668;
        51:
            _4705 <= _2659;
        52:
            _4705 <= _2650;
        53:
            _4705 <= _2641;
        54:
            _4705 <= _2632;
        55:
            _4705 <= _2623;
        56:
            _4705 <= _2614;
        57:
            _4705 <= _2605;
        58:
            _4705 <= _2596;
        59:
            _4705 <= _2587;
        60:
            _4705 <= _2578;
        61:
            _4705 <= _2569;
        62:
            _4705 <= _2560;
        63:
            _4705 <= _2551;
        64:
            _4705 <= _2542;
        65:
            _4705 <= _2533;
        66:
            _4705 <= _2524;
        67:
            _4705 <= _2515;
        68:
            _4705 <= _2506;
        69:
            _4705 <= _2497;
        70:
            _4705 <= _2488;
        71:
            _4705 <= _2479;
        72:
            _4705 <= _2470;
        73:
            _4705 <= _2461;
        74:
            _4705 <= _2452;
        75:
            _4705 <= _2443;
        76:
            _4705 <= _2434;
        77:
            _4705 <= _2425;
        78:
            _4705 <= _2416;
        79:
            _4705 <= _2407;
        80:
            _4705 <= _2398;
        81:
            _4705 <= _2389;
        82:
            _4705 <= _2380;
        83:
            _4705 <= _2371;
        84:
            _4705 <= _2362;
        85:
            _4705 <= _2353;
        86:
            _4705 <= _2344;
        87:
            _4705 <= _2335;
        88:
            _4705 <= _2326;
        89:
            _4705 <= _2317;
        90:
            _4705 <= _2308;
        91:
            _4705 <= _2299;
        92:
            _4705 <= _2290;
        93:
            _4705 <= _2281;
        94:
            _4705 <= _2272;
        95:
            _4705 <= _2263;
        96:
            _4705 <= _2254;
        97:
            _4705 <= _2245;
        98:
            _4705 <= _2236;
        99:
            _4705 <= _2227;
        100:
            _4705 <= _2218;
        101:
            _4705 <= _2209;
        102:
            _4705 <= _2200;
        103:
            _4705 <= _2191;
        104:
            _4705 <= _2182;
        105:
            _4705 <= _2173;
        106:
            _4705 <= _2164;
        107:
            _4705 <= _2155;
        108:
            _4705 <= _2146;
        109:
            _4705 <= _2137;
        110:
            _4705 <= _2128;
        111:
            _4705 <= _2119;
        112:
            _4705 <= _2110;
        113:
            _4705 <= _2101;
        114:
            _4705 <= _2092;
        115:
            _4705 <= _2083;
        116:
            _4705 <= _2074;
        117:
            _4705 <= _2065;
        118:
            _4705 <= _2056;
        119:
            _4705 <= _2047;
        120:
            _4705 <= _2038;
        121:
            _4705 <= _2029;
        122:
            _4705 <= _2020;
        123:
            _4705 <= _2011;
        124:
            _4705 <= _2002;
        125:
            _4705 <= _1993;
        126:
            _4705 <= _1984;
        127:
            _4705 <= _1975;
        128:
            _4705 <= _1966;
        129:
            _4705 <= _1957;
        130:
            _4705 <= _1948;
        131:
            _4705 <= _1939;
        132:
            _4705 <= _1930;
        133:
            _4705 <= _1921;
        134:
            _4705 <= _1912;
        135:
            _4705 <= _1903;
        136:
            _4705 <= _1894;
        137:
            _4705 <= _1885;
        138:
            _4705 <= _1876;
        139:
            _4705 <= _1867;
        140:
            _4705 <= _1858;
        141:
            _4705 <= _1849;
        142:
            _4705 <= _1840;
        143:
            _4705 <= _1831;
        144:
            _4705 <= _1822;
        145:
            _4705 <= _1813;
        146:
            _4705 <= _1804;
        147:
            _4705 <= _1795;
        148:
            _4705 <= _1786;
        149:
            _4705 <= _1777;
        150:
            _4705 <= _1768;
        151:
            _4705 <= _1759;
        152:
            _4705 <= _1750;
        153:
            _4705 <= _1741;
        154:
            _4705 <= _1732;
        155:
            _4705 <= _1723;
        156:
            _4705 <= _1714;
        157:
            _4705 <= _1705;
        158:
            _4705 <= _1696;
        159:
            _4705 <= _1687;
        160:
            _4705 <= _1678;
        161:
            _4705 <= _1669;
        162:
            _4705 <= _1660;
        163:
            _4705 <= _1651;
        164:
            _4705 <= _1642;
        165:
            _4705 <= _1633;
        166:
            _4705 <= _1624;
        167:
            _4705 <= _1615;
        168:
            _4705 <= _1606;
        169:
            _4705 <= _1597;
        170:
            _4705 <= _1588;
        171:
            _4705 <= _1579;
        172:
            _4705 <= _1570;
        173:
            _4705 <= _1561;
        174:
            _4705 <= _1552;
        175:
            _4705 <= _1543;
        176:
            _4705 <= _1534;
        177:
            _4705 <= _1525;
        178:
            _4705 <= _1516;
        179:
            _4705 <= _1507;
        180:
            _4705 <= _1498;
        181:
            _4705 <= _1489;
        182:
            _4705 <= _1480;
        183:
            _4705 <= _1471;
        184:
            _4705 <= _1462;
        185:
            _4705 <= _1453;
        186:
            _4705 <= _1444;
        187:
            _4705 <= _1435;
        188:
            _4705 <= _1426;
        189:
            _4705 <= _1417;
        190:
            _4705 <= _1408;
        191:
            _4705 <= _1399;
        192:
            _4705 <= _1390;
        193:
            _4705 <= _1381;
        194:
            _4705 <= _1372;
        195:
            _4705 <= _1363;
        196:
            _4705 <= _1354;
        197:
            _4705 <= _1345;
        198:
            _4705 <= _1336;
        199:
            _4705 <= _1327;
        200:
            _4705 <= _1318;
        201:
            _4705 <= _1309;
        202:
            _4705 <= _1300;
        203:
            _4705 <= _1291;
        204:
            _4705 <= _1282;
        205:
            _4705 <= _1273;
        206:
            _4705 <= _1264;
        207:
            _4705 <= _1255;
        208:
            _4705 <= _1246;
        209:
            _4705 <= _1237;
        210:
            _4705 <= _1228;
        211:
            _4705 <= _1219;
        212:
            _4705 <= _1210;
        213:
            _4705 <= _1201;
        214:
            _4705 <= _1192;
        215:
            _4705 <= _1183;
        216:
            _4705 <= _1174;
        217:
            _4705 <= _1165;
        218:
            _4705 <= _1156;
        219:
            _4705 <= _1147;
        220:
            _4705 <= _1138;
        221:
            _4705 <= _1129;
        222:
            _4705 <= _1120;
        223:
            _4705 <= _1111;
        224:
            _4705 <= _1102;
        225:
            _4705 <= _1093;
        226:
            _4705 <= _1084;
        227:
            _4705 <= _1075;
        228:
            _4705 <= _1066;
        229:
            _4705 <= _1057;
        230:
            _4705 <= _1048;
        231:
            _4705 <= _1039;
        232:
            _4705 <= _1030;
        233:
            _4705 <= _1021;
        234:
            _4705 <= _1012;
        235:
            _4705 <= _1003;
        236:
            _4705 <= _994;
        237:
            _4705 <= _985;
        238:
            _4705 <= _976;
        239:
            _4705 <= _967;
        240:
            _4705 <= _958;
        241:
            _4705 <= _949;
        242:
            _4705 <= _940;
        243:
            _4705 <= _931;
        244:
            _4705 <= _922;
        245:
            _4705 <= _913;
        246:
            _4705 <= _904;
        247:
            _4705 <= _895;
        248:
            _4705 <= _886;
        249:
            _4705 <= _877;
        250:
            _4705 <= _868;
        251:
            _4705 <= _859;
        252:
            _4705 <= _850;
        253:
            _4705 <= _841;
        254:
            _4705 <= _832;
        default:
            _4705 <= _823;
        endcase
    end
    assign _4706 = { _4707,
                     _4705 };
    assign _4710 = _4706 * _4709;
    assign _4711 = _4710[63:0];
    assign _4703 = _805 ? _4700 : _4701;
    assign _4712 = _4698 ? _4711 : _4703;
    assign _261 = _4712;
    always @(posedge _791) begin
        if (_789)
            _4701 <= _4700;
        else
            _4701 <= _261;
    end
    assign _4718 = 16'b0000000000000000;
    assign _5251 = _4719 < _5245;
    assign _5252 = _5251 ? _5245 : _4719;
    assign _5253 = _5250 ? _5249 : _5252;
    assign _5254 = _5246 ? _5249 : _5253;
    assign _4721 = _805 ? _4718 : _4719;
    assign _4723 = _4716 ? _4718 : _4721;
    assign _5255 = _4714 ? _5254 : _4723;
    assign _263 = _5255;
    always @(posedge _791) begin
        if (_789)
            _4719 <= _4718;
        else
            _4719 <= _263;
    end
    assign _5282 = 48'b000000000000000000000000000000000000000000000000;
    assign _5283 = { _5282,
                     _4719 };
    assign _5250 = _5249 < _5245;
    assign _5260 = _5250 ? _5245 : _5249;
    assign _5261 = _5246 ? _4726 : _5260;
    assign _5257 = _805 ? _4718 : _5249;
    assign _5259 = _4716 ? _4718 : _5257;
    assign _5262 = _4714 ? _5261 : _5259;
    assign _264 = _5262;
    always @(posedge _791) begin
        if (_789)
            _5249 <= _4718;
        else
            _5249 <= _264;
    end
    assign _5279 = { _5282,
                     _5249 };
    always @* begin
        case (_4729)
        0:
            _5244 <= _3925;
        1:
            _5244 <= _3928;
        2:
            _5244 <= _3931;
        3:
            _5244 <= _3934;
        4:
            _5244 <= _3937;
        5:
            _5244 <= _3940;
        6:
            _5244 <= _3943;
        7:
            _5244 <= _3946;
        8:
            _5244 <= _3949;
        9:
            _5244 <= _3952;
        10:
            _5244 <= _3955;
        11:
            _5244 <= _3958;
        12:
            _5244 <= _3961;
        13:
            _5244 <= _3964;
        14:
            _5244 <= _3967;
        15:
            _5244 <= _3970;
        16:
            _5244 <= _3973;
        17:
            _5244 <= _3976;
        18:
            _5244 <= _3979;
        19:
            _5244 <= _3982;
        20:
            _5244 <= _3985;
        21:
            _5244 <= _3988;
        22:
            _5244 <= _3991;
        23:
            _5244 <= _3994;
        24:
            _5244 <= _3997;
        25:
            _5244 <= _4000;
        26:
            _5244 <= _4003;
        27:
            _5244 <= _4006;
        28:
            _5244 <= _4009;
        29:
            _5244 <= _4012;
        30:
            _5244 <= _4015;
        31:
            _5244 <= _4018;
        32:
            _5244 <= _4021;
        33:
            _5244 <= _4024;
        34:
            _5244 <= _4027;
        35:
            _5244 <= _4030;
        36:
            _5244 <= _4033;
        37:
            _5244 <= _4036;
        38:
            _5244 <= _4039;
        39:
            _5244 <= _4042;
        40:
            _5244 <= _4045;
        41:
            _5244 <= _4048;
        42:
            _5244 <= _4051;
        43:
            _5244 <= _4054;
        44:
            _5244 <= _4057;
        45:
            _5244 <= _4060;
        46:
            _5244 <= _4063;
        47:
            _5244 <= _4066;
        48:
            _5244 <= _4069;
        49:
            _5244 <= _4072;
        50:
            _5244 <= _4075;
        51:
            _5244 <= _4078;
        52:
            _5244 <= _4081;
        53:
            _5244 <= _4084;
        54:
            _5244 <= _4087;
        55:
            _5244 <= _4090;
        56:
            _5244 <= _4093;
        57:
            _5244 <= _4096;
        58:
            _5244 <= _4099;
        59:
            _5244 <= _4102;
        60:
            _5244 <= _4105;
        61:
            _5244 <= _4108;
        62:
            _5244 <= _4111;
        63:
            _5244 <= _4114;
        64:
            _5244 <= _4117;
        65:
            _5244 <= _4120;
        66:
            _5244 <= _4123;
        67:
            _5244 <= _4126;
        68:
            _5244 <= _4129;
        69:
            _5244 <= _4132;
        70:
            _5244 <= _4135;
        71:
            _5244 <= _4138;
        72:
            _5244 <= _4141;
        73:
            _5244 <= _4144;
        74:
            _5244 <= _4147;
        75:
            _5244 <= _4150;
        76:
            _5244 <= _4153;
        77:
            _5244 <= _4156;
        78:
            _5244 <= _4159;
        79:
            _5244 <= _4162;
        80:
            _5244 <= _4165;
        81:
            _5244 <= _4168;
        82:
            _5244 <= _4171;
        83:
            _5244 <= _4174;
        84:
            _5244 <= _4177;
        85:
            _5244 <= _4180;
        86:
            _5244 <= _4183;
        87:
            _5244 <= _4186;
        88:
            _5244 <= _4189;
        89:
            _5244 <= _4192;
        90:
            _5244 <= _4195;
        91:
            _5244 <= _4198;
        92:
            _5244 <= _4201;
        93:
            _5244 <= _4204;
        94:
            _5244 <= _4207;
        95:
            _5244 <= _4210;
        96:
            _5244 <= _4213;
        97:
            _5244 <= _4216;
        98:
            _5244 <= _4219;
        99:
            _5244 <= _4222;
        100:
            _5244 <= _4225;
        101:
            _5244 <= _4228;
        102:
            _5244 <= _4231;
        103:
            _5244 <= _4234;
        104:
            _5244 <= _4237;
        105:
            _5244 <= _4240;
        106:
            _5244 <= _4243;
        107:
            _5244 <= _4246;
        108:
            _5244 <= _4249;
        109:
            _5244 <= _4252;
        110:
            _5244 <= _4255;
        111:
            _5244 <= _4258;
        112:
            _5244 <= _4261;
        113:
            _5244 <= _4264;
        114:
            _5244 <= _4267;
        115:
            _5244 <= _4270;
        116:
            _5244 <= _4273;
        117:
            _5244 <= _4276;
        118:
            _5244 <= _4279;
        119:
            _5244 <= _4282;
        120:
            _5244 <= _4285;
        121:
            _5244 <= _4288;
        122:
            _5244 <= _4291;
        123:
            _5244 <= _4294;
        124:
            _5244 <= _4297;
        125:
            _5244 <= _4300;
        126:
            _5244 <= _4303;
        127:
            _5244 <= _4306;
        128:
            _5244 <= _4309;
        129:
            _5244 <= _4312;
        130:
            _5244 <= _4315;
        131:
            _5244 <= _4318;
        132:
            _5244 <= _4321;
        133:
            _5244 <= _4324;
        134:
            _5244 <= _4327;
        135:
            _5244 <= _4330;
        136:
            _5244 <= _4333;
        137:
            _5244 <= _4336;
        138:
            _5244 <= _4339;
        139:
            _5244 <= _4342;
        140:
            _5244 <= _4345;
        141:
            _5244 <= _4348;
        142:
            _5244 <= _4351;
        143:
            _5244 <= _4354;
        144:
            _5244 <= _4357;
        145:
            _5244 <= _4360;
        146:
            _5244 <= _4363;
        147:
            _5244 <= _4366;
        148:
            _5244 <= _4369;
        149:
            _5244 <= _4372;
        150:
            _5244 <= _4375;
        151:
            _5244 <= _4378;
        152:
            _5244 <= _4381;
        153:
            _5244 <= _4384;
        154:
            _5244 <= _4387;
        155:
            _5244 <= _4390;
        156:
            _5244 <= _4393;
        157:
            _5244 <= _4396;
        158:
            _5244 <= _4399;
        159:
            _5244 <= _4402;
        160:
            _5244 <= _4405;
        161:
            _5244 <= _4408;
        162:
            _5244 <= _4411;
        163:
            _5244 <= _4414;
        164:
            _5244 <= _4417;
        165:
            _5244 <= _4420;
        166:
            _5244 <= _4423;
        167:
            _5244 <= _4426;
        168:
            _5244 <= _4429;
        169:
            _5244 <= _4432;
        170:
            _5244 <= _4435;
        171:
            _5244 <= _4438;
        172:
            _5244 <= _4441;
        173:
            _5244 <= _4444;
        174:
            _5244 <= _4447;
        175:
            _5244 <= _4450;
        176:
            _5244 <= _4453;
        177:
            _5244 <= _4456;
        178:
            _5244 <= _4459;
        179:
            _5244 <= _4462;
        180:
            _5244 <= _4465;
        181:
            _5244 <= _4468;
        182:
            _5244 <= _4471;
        183:
            _5244 <= _4474;
        184:
            _5244 <= _4477;
        185:
            _5244 <= _4480;
        186:
            _5244 <= _4483;
        187:
            _5244 <= _4486;
        188:
            _5244 <= _4489;
        189:
            _5244 <= _4492;
        190:
            _5244 <= _4495;
        191:
            _5244 <= _4498;
        192:
            _5244 <= _4501;
        193:
            _5244 <= _4504;
        194:
            _5244 <= _4507;
        195:
            _5244 <= _4510;
        196:
            _5244 <= _4513;
        197:
            _5244 <= _4516;
        198:
            _5244 <= _4519;
        199:
            _5244 <= _4522;
        200:
            _5244 <= _4525;
        201:
            _5244 <= _4528;
        202:
            _5244 <= _4531;
        203:
            _5244 <= _4534;
        204:
            _5244 <= _4537;
        205:
            _5244 <= _4540;
        206:
            _5244 <= _4543;
        207:
            _5244 <= _4546;
        208:
            _5244 <= _4549;
        209:
            _5244 <= _4552;
        210:
            _5244 <= _4555;
        211:
            _5244 <= _4558;
        212:
            _5244 <= _4561;
        213:
            _5244 <= _4564;
        214:
            _5244 <= _4567;
        215:
            _5244 <= _4570;
        216:
            _5244 <= _4573;
        217:
            _5244 <= _4576;
        218:
            _5244 <= _4579;
        219:
            _5244 <= _4582;
        220:
            _5244 <= _4585;
        221:
            _5244 <= _4588;
        222:
            _5244 <= _4591;
        223:
            _5244 <= _4594;
        224:
            _5244 <= _4597;
        225:
            _5244 <= _4600;
        226:
            _5244 <= _4603;
        227:
            _5244 <= _4606;
        228:
            _5244 <= _4609;
        229:
            _5244 <= _4612;
        230:
            _5244 <= _4615;
        231:
            _5244 <= _4618;
        232:
            _5244 <= _4621;
        233:
            _5244 <= _4624;
        234:
            _5244 <= _4627;
        235:
            _5244 <= _4630;
        236:
            _5244 <= _4633;
        237:
            _5244 <= _4636;
        238:
            _5244 <= _4639;
        239:
            _5244 <= _4642;
        240:
            _5244 <= _4645;
        241:
            _5244 <= _4648;
        242:
            _5244 <= _4651;
        243:
            _5244 <= _4654;
        244:
            _5244 <= _4657;
        245:
            _5244 <= _4660;
        246:
            _5244 <= _4663;
        247:
            _5244 <= _4666;
        248:
            _5244 <= _4669;
        249:
            _5244 <= _4672;
        250:
            _5244 <= _4675;
        251:
            _5244 <= _4678;
        252:
            _5244 <= _4681;
        253:
            _5244 <= _4684;
        254:
            _5244 <= _4687;
        default:
            _5244 <= _4690;
        endcase
    end
    assign _5241 = _3903 == _818;
    assign _5239 = _3900 == _827;
    assign _5237 = _3897 == _836;
    assign _5235 = _3894 == _845;
    assign _5233 = _3891 == _854;
    assign _5231 = _3888 == _863;
    assign _5229 = _3885 == _872;
    assign _5227 = _3882 == _881;
    assign _5225 = _3879 == _890;
    assign _5223 = _3876 == _899;
    assign _5221 = _3873 == _908;
    assign _5219 = _3870 == _917;
    assign _5217 = _3867 == _926;
    assign _5215 = _3864 == _935;
    assign _5213 = _3861 == _944;
    assign _5211 = _3858 == _953;
    assign _5209 = _3855 == _962;
    assign _5207 = _3852 == _971;
    assign _5205 = _3849 == _980;
    assign _5203 = _3846 == _989;
    assign _5201 = _3843 == _998;
    assign _5199 = _3840 == _1007;
    assign _5197 = _3837 == _1016;
    assign _5195 = _3834 == _1025;
    assign _5193 = _3831 == _1034;
    assign _5191 = _3828 == _1043;
    assign _5189 = _3825 == _1052;
    assign _5187 = _3822 == _1061;
    assign _5185 = _3819 == _1070;
    assign _5183 = _3816 == _1079;
    assign _5181 = _3813 == _1088;
    assign _5179 = _3810 == _1097;
    assign _5177 = _3807 == _1106;
    assign _5175 = _3804 == _1115;
    assign _5173 = _3801 == _1124;
    assign _5171 = _3798 == _1133;
    assign _5169 = _3795 == _1142;
    assign _5167 = _3792 == _1151;
    assign _5165 = _3789 == _1160;
    assign _5163 = _3786 == _1169;
    assign _5161 = _3783 == _1178;
    assign _5159 = _3780 == _1187;
    assign _5157 = _3777 == _1196;
    assign _5155 = _3774 == _1205;
    assign _5153 = _3771 == _1214;
    assign _5151 = _3768 == _1223;
    assign _5149 = _3765 == _1232;
    assign _5147 = _3762 == _1241;
    assign _5145 = _3759 == _1250;
    assign _5143 = _3756 == _1259;
    assign _5141 = _3753 == _1268;
    assign _5139 = _3750 == _1277;
    assign _5137 = _3747 == _1286;
    assign _5135 = _3744 == _1295;
    assign _5133 = _3741 == _1304;
    assign _5131 = _3738 == _1313;
    assign _5129 = _3735 == _1322;
    assign _5127 = _3732 == _1331;
    assign _5125 = _3729 == _1340;
    assign _5123 = _3726 == _1349;
    assign _5121 = _3723 == _1358;
    assign _5119 = _3720 == _1367;
    assign _5117 = _3717 == _1376;
    assign _5115 = _3714 == _1385;
    assign _5113 = _3711 == _1394;
    assign _5111 = _3708 == _1403;
    assign _5109 = _3705 == _1412;
    assign _5107 = _3702 == _1421;
    assign _5105 = _3699 == _1430;
    assign _5103 = _3696 == _1439;
    assign _5101 = _3693 == _1448;
    assign _5099 = _3690 == _1457;
    assign _5097 = _3687 == _1466;
    assign _5095 = _3684 == _1475;
    assign _5093 = _3681 == _1484;
    assign _5091 = _3678 == _1493;
    assign _5089 = _3675 == _1502;
    assign _5087 = _3672 == _1511;
    assign _5085 = _3669 == _1520;
    assign _5083 = _3666 == _1529;
    assign _5081 = _3663 == _1538;
    assign _5079 = _3660 == _1547;
    assign _5077 = _3657 == _1556;
    assign _5075 = _3654 == _1565;
    assign _5073 = _3651 == _1574;
    assign _5071 = _3648 == _1583;
    assign _5069 = _3645 == _1592;
    assign _5067 = _3642 == _1601;
    assign _5065 = _3639 == _1610;
    assign _5063 = _3636 == _1619;
    assign _5061 = _3633 == _1628;
    assign _5059 = _3630 == _1637;
    assign _5057 = _3627 == _1646;
    assign _5055 = _3624 == _1655;
    assign _5053 = _3621 == _1664;
    assign _5051 = _3618 == _1673;
    assign _5049 = _3615 == _1682;
    assign _5047 = _3612 == _1691;
    assign _5045 = _3609 == _1700;
    assign _5043 = _3606 == _1709;
    assign _5041 = _3603 == _1718;
    assign _5039 = _3600 == _1727;
    assign _5037 = _3597 == _1736;
    assign _5035 = _3594 == _1745;
    assign _5033 = _3591 == _1754;
    assign _5031 = _3588 == _1763;
    assign _5029 = _3585 == _1772;
    assign _5027 = _3582 == _1781;
    assign _5025 = _3579 == _1790;
    assign _5023 = _3576 == _1799;
    assign _5021 = _3573 == _1808;
    assign _5019 = _3570 == _1817;
    assign _5017 = _3567 == _1826;
    assign _5015 = _3564 == _1835;
    assign _5013 = _3561 == _1844;
    assign _5011 = _3558 == _1853;
    assign _5009 = _3555 == _1862;
    assign _5007 = _3552 == _1871;
    assign _5005 = _3549 == _1880;
    assign _5003 = _3546 == _1889;
    assign _5001 = _3543 == _1898;
    assign _4999 = _3540 == _1907;
    assign _4997 = _3537 == _1916;
    assign _4995 = _3534 == _1925;
    assign _4993 = _3531 == _1934;
    assign _4991 = _3528 == _1943;
    assign _4989 = _3525 == _1952;
    assign _4987 = _3522 == _1961;
    assign _4985 = _3519 == _1970;
    assign _4983 = _3516 == _1979;
    assign _4981 = _3513 == _1988;
    assign _4979 = _3510 == _1997;
    assign _4977 = _3507 == _2006;
    assign _4975 = _3504 == _2015;
    assign _4973 = _3501 == _2024;
    assign _4971 = _3498 == _2033;
    assign _4969 = _3495 == _2042;
    assign _4967 = _3492 == _2051;
    assign _4965 = _3489 == _2060;
    assign _4963 = _3486 == _2069;
    assign _4961 = _3483 == _2078;
    assign _4959 = _3480 == _2087;
    assign _4957 = _3477 == _2096;
    assign _4955 = _3474 == _2105;
    assign _4953 = _3471 == _2114;
    assign _4951 = _3468 == _2123;
    assign _4949 = _3465 == _2132;
    assign _4947 = _3462 == _2141;
    assign _4945 = _3459 == _2150;
    assign _4943 = _3456 == _2159;
    assign _4941 = _3453 == _2168;
    assign _4939 = _3450 == _2177;
    assign _4937 = _3447 == _2186;
    assign _4935 = _3444 == _2195;
    assign _4933 = _3441 == _2204;
    assign _4931 = _3438 == _2213;
    assign _4929 = _3435 == _2222;
    assign _4927 = _3432 == _2231;
    assign _4925 = _3429 == _2240;
    assign _4923 = _3426 == _2249;
    assign _4921 = _3423 == _2258;
    assign _4919 = _3420 == _2267;
    assign _4917 = _3417 == _2276;
    assign _4915 = _3414 == _2285;
    assign _4913 = _3411 == _2294;
    assign _4911 = _3408 == _2303;
    assign _4909 = _3405 == _2312;
    assign _4907 = _3402 == _2321;
    assign _4905 = _3399 == _2330;
    assign _4903 = _3396 == _2339;
    assign _4901 = _3393 == _2348;
    assign _4899 = _3390 == _2357;
    assign _4897 = _3387 == _2366;
    assign _4895 = _3384 == _2375;
    assign _4893 = _3381 == _2384;
    assign _4891 = _3378 == _2393;
    assign _4889 = _3375 == _2402;
    assign _4887 = _3372 == _2411;
    assign _4885 = _3369 == _2420;
    assign _4883 = _3366 == _2429;
    assign _4881 = _3363 == _2438;
    assign _4879 = _3360 == _2447;
    assign _4877 = _3357 == _2456;
    assign _4875 = _3354 == _2465;
    assign _4873 = _3351 == _2474;
    assign _4871 = _3348 == _2483;
    assign _4869 = _3345 == _2492;
    assign _4867 = _3342 == _2501;
    assign _4865 = _3339 == _2510;
    assign _4863 = _3336 == _2519;
    assign _4861 = _3333 == _2528;
    assign _4859 = _3330 == _2537;
    assign _4857 = _3327 == _2546;
    assign _4855 = _3324 == _2555;
    assign _4853 = _3321 == _2564;
    assign _4851 = _3318 == _2573;
    assign _4849 = _3315 == _2582;
    assign _4847 = _3312 == _2591;
    assign _4845 = _3309 == _2600;
    assign _4843 = _3306 == _2609;
    assign _4841 = _3303 == _2618;
    assign _4839 = _3300 == _2627;
    assign _4837 = _3297 == _2636;
    assign _4835 = _3294 == _2645;
    assign _4833 = _3291 == _2654;
    assign _4831 = _3288 == _2663;
    assign _4829 = _3285 == _2672;
    assign _4827 = _3282 == _2681;
    assign _4825 = _3279 == _2690;
    assign _4823 = _3276 == _2699;
    assign _4821 = _3273 == _2708;
    assign _4819 = _3270 == _2717;
    assign _4817 = _3267 == _2726;
    assign _4815 = _3264 == _2735;
    assign _4813 = _3261 == _2744;
    assign _4811 = _3258 == _2753;
    assign _4809 = _3255 == _2762;
    assign _4807 = _3252 == _2771;
    assign _4805 = _3249 == _2780;
    assign _4803 = _3246 == _2789;
    assign _4801 = _3243 == _2798;
    assign _4799 = _3240 == _2807;
    assign _4797 = _3237 == _2816;
    assign _4795 = _3234 == _2825;
    assign _4793 = _3231 == _2834;
    assign _4791 = _3228 == _2843;
    assign _4789 = _3225 == _2852;
    assign _4787 = _3222 == _2861;
    assign _4785 = _3219 == _2870;
    assign _4783 = _3216 == _2879;
    assign _4781 = _3213 == _2888;
    assign _4779 = _3210 == _2897;
    assign _4777 = _3207 == _2906;
    assign _4775 = _3204 == _2915;
    assign _4773 = _3201 == _2924;
    assign _4771 = _3198 == _2933;
    assign _4769 = _3195 == _2942;
    assign _4767 = _3192 == _2951;
    assign _4765 = _3189 == _2960;
    assign _4763 = _3186 == _2969;
    assign _4761 = _3183 == _2978;
    assign _4759 = _3180 == _2987;
    assign _4757 = _3177 == _2996;
    assign _4755 = _3174 == _3005;
    assign _4753 = _3171 == _3014;
    assign _4751 = _3168 == _3023;
    assign _4749 = _3165 == _3032;
    assign _4747 = _3162 == _3041;
    assign _4745 = _3159 == _3050;
    assign _4743 = _3156 == _3059;
    assign _4741 = _3153 == _3068;
    assign _4739 = _3150 == _3077;
    assign _4737 = _3147 == _3086;
    assign _4735 = _3144 == _3095;
    assign _4733 = _3141 == _3104;
    assign _4731 = _3138 == _3118;
    always @* begin
        case (_4729)
        0:
            _5242 <= _4731;
        1:
            _5242 <= _4733;
        2:
            _5242 <= _4735;
        3:
            _5242 <= _4737;
        4:
            _5242 <= _4739;
        5:
            _5242 <= _4741;
        6:
            _5242 <= _4743;
        7:
            _5242 <= _4745;
        8:
            _5242 <= _4747;
        9:
            _5242 <= _4749;
        10:
            _5242 <= _4751;
        11:
            _5242 <= _4753;
        12:
            _5242 <= _4755;
        13:
            _5242 <= _4757;
        14:
            _5242 <= _4759;
        15:
            _5242 <= _4761;
        16:
            _5242 <= _4763;
        17:
            _5242 <= _4765;
        18:
            _5242 <= _4767;
        19:
            _5242 <= _4769;
        20:
            _5242 <= _4771;
        21:
            _5242 <= _4773;
        22:
            _5242 <= _4775;
        23:
            _5242 <= _4777;
        24:
            _5242 <= _4779;
        25:
            _5242 <= _4781;
        26:
            _5242 <= _4783;
        27:
            _5242 <= _4785;
        28:
            _5242 <= _4787;
        29:
            _5242 <= _4789;
        30:
            _5242 <= _4791;
        31:
            _5242 <= _4793;
        32:
            _5242 <= _4795;
        33:
            _5242 <= _4797;
        34:
            _5242 <= _4799;
        35:
            _5242 <= _4801;
        36:
            _5242 <= _4803;
        37:
            _5242 <= _4805;
        38:
            _5242 <= _4807;
        39:
            _5242 <= _4809;
        40:
            _5242 <= _4811;
        41:
            _5242 <= _4813;
        42:
            _5242 <= _4815;
        43:
            _5242 <= _4817;
        44:
            _5242 <= _4819;
        45:
            _5242 <= _4821;
        46:
            _5242 <= _4823;
        47:
            _5242 <= _4825;
        48:
            _5242 <= _4827;
        49:
            _5242 <= _4829;
        50:
            _5242 <= _4831;
        51:
            _5242 <= _4833;
        52:
            _5242 <= _4835;
        53:
            _5242 <= _4837;
        54:
            _5242 <= _4839;
        55:
            _5242 <= _4841;
        56:
            _5242 <= _4843;
        57:
            _5242 <= _4845;
        58:
            _5242 <= _4847;
        59:
            _5242 <= _4849;
        60:
            _5242 <= _4851;
        61:
            _5242 <= _4853;
        62:
            _5242 <= _4855;
        63:
            _5242 <= _4857;
        64:
            _5242 <= _4859;
        65:
            _5242 <= _4861;
        66:
            _5242 <= _4863;
        67:
            _5242 <= _4865;
        68:
            _5242 <= _4867;
        69:
            _5242 <= _4869;
        70:
            _5242 <= _4871;
        71:
            _5242 <= _4873;
        72:
            _5242 <= _4875;
        73:
            _5242 <= _4877;
        74:
            _5242 <= _4879;
        75:
            _5242 <= _4881;
        76:
            _5242 <= _4883;
        77:
            _5242 <= _4885;
        78:
            _5242 <= _4887;
        79:
            _5242 <= _4889;
        80:
            _5242 <= _4891;
        81:
            _5242 <= _4893;
        82:
            _5242 <= _4895;
        83:
            _5242 <= _4897;
        84:
            _5242 <= _4899;
        85:
            _5242 <= _4901;
        86:
            _5242 <= _4903;
        87:
            _5242 <= _4905;
        88:
            _5242 <= _4907;
        89:
            _5242 <= _4909;
        90:
            _5242 <= _4911;
        91:
            _5242 <= _4913;
        92:
            _5242 <= _4915;
        93:
            _5242 <= _4917;
        94:
            _5242 <= _4919;
        95:
            _5242 <= _4921;
        96:
            _5242 <= _4923;
        97:
            _5242 <= _4925;
        98:
            _5242 <= _4927;
        99:
            _5242 <= _4929;
        100:
            _5242 <= _4931;
        101:
            _5242 <= _4933;
        102:
            _5242 <= _4935;
        103:
            _5242 <= _4937;
        104:
            _5242 <= _4939;
        105:
            _5242 <= _4941;
        106:
            _5242 <= _4943;
        107:
            _5242 <= _4945;
        108:
            _5242 <= _4947;
        109:
            _5242 <= _4949;
        110:
            _5242 <= _4951;
        111:
            _5242 <= _4953;
        112:
            _5242 <= _4955;
        113:
            _5242 <= _4957;
        114:
            _5242 <= _4959;
        115:
            _5242 <= _4961;
        116:
            _5242 <= _4963;
        117:
            _5242 <= _4965;
        118:
            _5242 <= _4967;
        119:
            _5242 <= _4969;
        120:
            _5242 <= _4971;
        121:
            _5242 <= _4973;
        122:
            _5242 <= _4975;
        123:
            _5242 <= _4977;
        124:
            _5242 <= _4979;
        125:
            _5242 <= _4981;
        126:
            _5242 <= _4983;
        127:
            _5242 <= _4985;
        128:
            _5242 <= _4987;
        129:
            _5242 <= _4989;
        130:
            _5242 <= _4991;
        131:
            _5242 <= _4993;
        132:
            _5242 <= _4995;
        133:
            _5242 <= _4997;
        134:
            _5242 <= _4999;
        135:
            _5242 <= _5001;
        136:
            _5242 <= _5003;
        137:
            _5242 <= _5005;
        138:
            _5242 <= _5007;
        139:
            _5242 <= _5009;
        140:
            _5242 <= _5011;
        141:
            _5242 <= _5013;
        142:
            _5242 <= _5015;
        143:
            _5242 <= _5017;
        144:
            _5242 <= _5019;
        145:
            _5242 <= _5021;
        146:
            _5242 <= _5023;
        147:
            _5242 <= _5025;
        148:
            _5242 <= _5027;
        149:
            _5242 <= _5029;
        150:
            _5242 <= _5031;
        151:
            _5242 <= _5033;
        152:
            _5242 <= _5035;
        153:
            _5242 <= _5037;
        154:
            _5242 <= _5039;
        155:
            _5242 <= _5041;
        156:
            _5242 <= _5043;
        157:
            _5242 <= _5045;
        158:
            _5242 <= _5047;
        159:
            _5242 <= _5049;
        160:
            _5242 <= _5051;
        161:
            _5242 <= _5053;
        162:
            _5242 <= _5055;
        163:
            _5242 <= _5057;
        164:
            _5242 <= _5059;
        165:
            _5242 <= _5061;
        166:
            _5242 <= _5063;
        167:
            _5242 <= _5065;
        168:
            _5242 <= _5067;
        169:
            _5242 <= _5069;
        170:
            _5242 <= _5071;
        171:
            _5242 <= _5073;
        172:
            _5242 <= _5075;
        173:
            _5242 <= _5077;
        174:
            _5242 <= _5079;
        175:
            _5242 <= _5081;
        176:
            _5242 <= _5083;
        177:
            _5242 <= _5085;
        178:
            _5242 <= _5087;
        179:
            _5242 <= _5089;
        180:
            _5242 <= _5091;
        181:
            _5242 <= _5093;
        182:
            _5242 <= _5095;
        183:
            _5242 <= _5097;
        184:
            _5242 <= _5099;
        185:
            _5242 <= _5101;
        186:
            _5242 <= _5103;
        187:
            _5242 <= _5105;
        188:
            _5242 <= _5107;
        189:
            _5242 <= _5109;
        190:
            _5242 <= _5111;
        191:
            _5242 <= _5113;
        192:
            _5242 <= _5115;
        193:
            _5242 <= _5117;
        194:
            _5242 <= _5119;
        195:
            _5242 <= _5121;
        196:
            _5242 <= _5123;
        197:
            _5242 <= _5125;
        198:
            _5242 <= _5127;
        199:
            _5242 <= _5129;
        200:
            _5242 <= _5131;
        201:
            _5242 <= _5133;
        202:
            _5242 <= _5135;
        203:
            _5242 <= _5137;
        204:
            _5242 <= _5139;
        205:
            _5242 <= _5141;
        206:
            _5242 <= _5143;
        207:
            _5242 <= _5145;
        208:
            _5242 <= _5147;
        209:
            _5242 <= _5149;
        210:
            _5242 <= _5151;
        211:
            _5242 <= _5153;
        212:
            _5242 <= _5155;
        213:
            _5242 <= _5157;
        214:
            _5242 <= _5159;
        215:
            _5242 <= _5161;
        216:
            _5242 <= _5163;
        217:
            _5242 <= _5165;
        218:
            _5242 <= _5167;
        219:
            _5242 <= _5169;
        220:
            _5242 <= _5171;
        221:
            _5242 <= _5173;
        222:
            _5242 <= _5175;
        223:
            _5242 <= _5177;
        224:
            _5242 <= _5179;
        225:
            _5242 <= _5181;
        226:
            _5242 <= _5183;
        227:
            _5242 <= _5185;
        228:
            _5242 <= _5187;
        229:
            _5242 <= _5189;
        230:
            _5242 <= _5191;
        231:
            _5242 <= _5193;
        232:
            _5242 <= _5195;
        233:
            _5242 <= _5197;
        234:
            _5242 <= _5199;
        235:
            _5242 <= _5201;
        236:
            _5242 <= _5203;
        237:
            _5242 <= _5205;
        238:
            _5242 <= _5207;
        239:
            _5242 <= _5209;
        240:
            _5242 <= _5211;
        241:
            _5242 <= _5213;
        242:
            _5242 <= _5215;
        243:
            _5242 <= _5217;
        244:
            _5242 <= _5219;
        245:
            _5242 <= _5221;
        246:
            _5242 <= _5223;
        247:
            _5242 <= _5225;
        248:
            _5242 <= _5227;
        249:
            _5242 <= _5229;
        250:
            _5242 <= _5231;
        251:
            _5242 <= _5233;
        252:
            _5242 <= _5235;
        253:
            _5242 <= _5237;
        254:
            _5242 <= _5239;
        default:
            _5242 <= _5241;
        endcase
    end
    assign _5245 = _5242 ? _5244 : _4718;
    assign _5246 = _4726 < _5245;
    assign _5267 = _5246 ? _5245 : _4726;
    assign _5264 = _805 ? _4718 : _4726;
    assign _5266 = _4716 ? _4718 : _5264;
    assign _5268 = _4714 ? _5267 : _5266;
    assign _265 = _5268;
    always @(posedge _791) begin
        if (_789)
            _4726 <= _4718;
        else
            _4726 <= _265;
    end
    assign _5277 = { _5282,
                     _4726 };
    assign _5280 = _5277 * _5279;
    assign _5281 = _5280[63:0];
    assign _5284 = _5281 * _5283;
    assign _5285 = _5284[63:0];
    assign _5275 = _805 ? _4700 : _5273;
    assign _5286 = _5270 ? _5285 : _5275;
    assign _266 = _5286;
    always @(posedge _791) begin
        if (_789)
            _5273 <= _4700;
        else
            _5273 <= _266;
    end
    assign _5288 = _811 == _5287;
    assign _809 = 3'b000;
    assign _5287 = 3'b110;
    assign _11990 = _3132 & _3135;
    assign _11991 = _11990 & _793;
    assign _11992 = _11991 ? _5287 : _811;
    assign _4696 = { _3118,
                     _787 };
    assign _4694 = _3920 ? _4691 : _4693;
    assign _4697 = _4694 == _4696;
    assign _11940 = 16'b0000000000000001;
    assign _5306 = _5304 == _818;
    assign _5300 = ~ _3920;
    assign _5301 = _3135 & _5300;
    assign _5307 = _5301 & _5306;
    assign _5308 = _5307 ? _4693 : _4690;
    assign _5298 = _5296 == _818;
    assign _5299 = _5293 & _5298;
    assign _5310 = _5299 ? _11940 : _5308;
    assign _5312 = _805 ? _4718 : _5310;
    assign _270 = _5312;
    always @(posedge _791) begin
        if (_789)
            _4690 <= _4718;
        else
            _4690 <= _270;
    end
    assign _5319 = _5304 == _827;
    assign _5316 = ~ _3920;
    assign _5317 = _3135 & _5316;
    assign _5320 = _5317 & _5319;
    assign _5321 = _5320 ? _4693 : _4687;
    assign _5314 = _5296 == _827;
    assign _5315 = _5293 & _5314;
    assign _5323 = _5315 ? _11940 : _5321;
    assign _5325 = _805 ? _4718 : _5323;
    assign _271 = _5325;
    always @(posedge _791) begin
        if (_789)
            _4687 <= _4718;
        else
            _4687 <= _271;
    end
    assign _5332 = _5304 == _836;
    assign _5329 = ~ _3920;
    assign _5330 = _3135 & _5329;
    assign _5333 = _5330 & _5332;
    assign _5334 = _5333 ? _4693 : _4684;
    assign _5327 = _5296 == _836;
    assign _5328 = _5293 & _5327;
    assign _5336 = _5328 ? _11940 : _5334;
    assign _5338 = _805 ? _4718 : _5336;
    assign _272 = _5338;
    always @(posedge _791) begin
        if (_789)
            _4684 <= _4718;
        else
            _4684 <= _272;
    end
    assign _5345 = _5304 == _845;
    assign _5342 = ~ _3920;
    assign _5343 = _3135 & _5342;
    assign _5346 = _5343 & _5345;
    assign _5347 = _5346 ? _4693 : _4681;
    assign _5340 = _5296 == _845;
    assign _5341 = _5293 & _5340;
    assign _5349 = _5341 ? _11940 : _5347;
    assign _5351 = _805 ? _4718 : _5349;
    assign _273 = _5351;
    always @(posedge _791) begin
        if (_789)
            _4681 <= _4718;
        else
            _4681 <= _273;
    end
    assign _5358 = _5304 == _854;
    assign _5355 = ~ _3920;
    assign _5356 = _3135 & _5355;
    assign _5359 = _5356 & _5358;
    assign _5360 = _5359 ? _4693 : _4678;
    assign _5353 = _5296 == _854;
    assign _5354 = _5293 & _5353;
    assign _5362 = _5354 ? _11940 : _5360;
    assign _5364 = _805 ? _4718 : _5362;
    assign _274 = _5364;
    always @(posedge _791) begin
        if (_789)
            _4678 <= _4718;
        else
            _4678 <= _274;
    end
    assign _5371 = _5304 == _863;
    assign _5368 = ~ _3920;
    assign _5369 = _3135 & _5368;
    assign _5372 = _5369 & _5371;
    assign _5373 = _5372 ? _4693 : _4675;
    assign _5366 = _5296 == _863;
    assign _5367 = _5293 & _5366;
    assign _5375 = _5367 ? _11940 : _5373;
    assign _5377 = _805 ? _4718 : _5375;
    assign _275 = _5377;
    always @(posedge _791) begin
        if (_789)
            _4675 <= _4718;
        else
            _4675 <= _275;
    end
    assign _5384 = _5304 == _872;
    assign _5381 = ~ _3920;
    assign _5382 = _3135 & _5381;
    assign _5385 = _5382 & _5384;
    assign _5386 = _5385 ? _4693 : _4672;
    assign _5379 = _5296 == _872;
    assign _5380 = _5293 & _5379;
    assign _5388 = _5380 ? _11940 : _5386;
    assign _5390 = _805 ? _4718 : _5388;
    assign _276 = _5390;
    always @(posedge _791) begin
        if (_789)
            _4672 <= _4718;
        else
            _4672 <= _276;
    end
    assign _5397 = _5304 == _881;
    assign _5394 = ~ _3920;
    assign _5395 = _3135 & _5394;
    assign _5398 = _5395 & _5397;
    assign _5399 = _5398 ? _4693 : _4669;
    assign _5392 = _5296 == _881;
    assign _5393 = _5293 & _5392;
    assign _5401 = _5393 ? _11940 : _5399;
    assign _5403 = _805 ? _4718 : _5401;
    assign _277 = _5403;
    always @(posedge _791) begin
        if (_789)
            _4669 <= _4718;
        else
            _4669 <= _277;
    end
    assign _5410 = _5304 == _890;
    assign _5407 = ~ _3920;
    assign _5408 = _3135 & _5407;
    assign _5411 = _5408 & _5410;
    assign _5412 = _5411 ? _4693 : _4666;
    assign _5405 = _5296 == _890;
    assign _5406 = _5293 & _5405;
    assign _5414 = _5406 ? _11940 : _5412;
    assign _5416 = _805 ? _4718 : _5414;
    assign _278 = _5416;
    always @(posedge _791) begin
        if (_789)
            _4666 <= _4718;
        else
            _4666 <= _278;
    end
    assign _5423 = _5304 == _899;
    assign _5420 = ~ _3920;
    assign _5421 = _3135 & _5420;
    assign _5424 = _5421 & _5423;
    assign _5425 = _5424 ? _4693 : _4663;
    assign _5418 = _5296 == _899;
    assign _5419 = _5293 & _5418;
    assign _5427 = _5419 ? _11940 : _5425;
    assign _5429 = _805 ? _4718 : _5427;
    assign _279 = _5429;
    always @(posedge _791) begin
        if (_789)
            _4663 <= _4718;
        else
            _4663 <= _279;
    end
    assign _5436 = _5304 == _908;
    assign _5433 = ~ _3920;
    assign _5434 = _3135 & _5433;
    assign _5437 = _5434 & _5436;
    assign _5438 = _5437 ? _4693 : _4660;
    assign _5431 = _5296 == _908;
    assign _5432 = _5293 & _5431;
    assign _5440 = _5432 ? _11940 : _5438;
    assign _5442 = _805 ? _4718 : _5440;
    assign _280 = _5442;
    always @(posedge _791) begin
        if (_789)
            _4660 <= _4718;
        else
            _4660 <= _280;
    end
    assign _5449 = _5304 == _917;
    assign _5446 = ~ _3920;
    assign _5447 = _3135 & _5446;
    assign _5450 = _5447 & _5449;
    assign _5451 = _5450 ? _4693 : _4657;
    assign _5444 = _5296 == _917;
    assign _5445 = _5293 & _5444;
    assign _5453 = _5445 ? _11940 : _5451;
    assign _5455 = _805 ? _4718 : _5453;
    assign _281 = _5455;
    always @(posedge _791) begin
        if (_789)
            _4657 <= _4718;
        else
            _4657 <= _281;
    end
    assign _5462 = _5304 == _926;
    assign _5459 = ~ _3920;
    assign _5460 = _3135 & _5459;
    assign _5463 = _5460 & _5462;
    assign _5464 = _5463 ? _4693 : _4654;
    assign _5457 = _5296 == _926;
    assign _5458 = _5293 & _5457;
    assign _5466 = _5458 ? _11940 : _5464;
    assign _5468 = _805 ? _4718 : _5466;
    assign _282 = _5468;
    always @(posedge _791) begin
        if (_789)
            _4654 <= _4718;
        else
            _4654 <= _282;
    end
    assign _5475 = _5304 == _935;
    assign _5472 = ~ _3920;
    assign _5473 = _3135 & _5472;
    assign _5476 = _5473 & _5475;
    assign _5477 = _5476 ? _4693 : _4651;
    assign _5470 = _5296 == _935;
    assign _5471 = _5293 & _5470;
    assign _5479 = _5471 ? _11940 : _5477;
    assign _5481 = _805 ? _4718 : _5479;
    assign _283 = _5481;
    always @(posedge _791) begin
        if (_789)
            _4651 <= _4718;
        else
            _4651 <= _283;
    end
    assign _5488 = _5304 == _944;
    assign _5485 = ~ _3920;
    assign _5486 = _3135 & _5485;
    assign _5489 = _5486 & _5488;
    assign _5490 = _5489 ? _4693 : _4648;
    assign _5483 = _5296 == _944;
    assign _5484 = _5293 & _5483;
    assign _5492 = _5484 ? _11940 : _5490;
    assign _5494 = _805 ? _4718 : _5492;
    assign _284 = _5494;
    always @(posedge _791) begin
        if (_789)
            _4648 <= _4718;
        else
            _4648 <= _284;
    end
    assign _5501 = _5304 == _953;
    assign _5498 = ~ _3920;
    assign _5499 = _3135 & _5498;
    assign _5502 = _5499 & _5501;
    assign _5503 = _5502 ? _4693 : _4645;
    assign _5496 = _5296 == _953;
    assign _5497 = _5293 & _5496;
    assign _5505 = _5497 ? _11940 : _5503;
    assign _5507 = _805 ? _4718 : _5505;
    assign _285 = _5507;
    always @(posedge _791) begin
        if (_789)
            _4645 <= _4718;
        else
            _4645 <= _285;
    end
    assign _5514 = _5304 == _962;
    assign _5511 = ~ _3920;
    assign _5512 = _3135 & _5511;
    assign _5515 = _5512 & _5514;
    assign _5516 = _5515 ? _4693 : _4642;
    assign _5509 = _5296 == _962;
    assign _5510 = _5293 & _5509;
    assign _5518 = _5510 ? _11940 : _5516;
    assign _5520 = _805 ? _4718 : _5518;
    assign _286 = _5520;
    always @(posedge _791) begin
        if (_789)
            _4642 <= _4718;
        else
            _4642 <= _286;
    end
    assign _5527 = _5304 == _971;
    assign _5524 = ~ _3920;
    assign _5525 = _3135 & _5524;
    assign _5528 = _5525 & _5527;
    assign _5529 = _5528 ? _4693 : _4639;
    assign _5522 = _5296 == _971;
    assign _5523 = _5293 & _5522;
    assign _5531 = _5523 ? _11940 : _5529;
    assign _5533 = _805 ? _4718 : _5531;
    assign _287 = _5533;
    always @(posedge _791) begin
        if (_789)
            _4639 <= _4718;
        else
            _4639 <= _287;
    end
    assign _5540 = _5304 == _980;
    assign _5537 = ~ _3920;
    assign _5538 = _3135 & _5537;
    assign _5541 = _5538 & _5540;
    assign _5542 = _5541 ? _4693 : _4636;
    assign _5535 = _5296 == _980;
    assign _5536 = _5293 & _5535;
    assign _5544 = _5536 ? _11940 : _5542;
    assign _5546 = _805 ? _4718 : _5544;
    assign _288 = _5546;
    always @(posedge _791) begin
        if (_789)
            _4636 <= _4718;
        else
            _4636 <= _288;
    end
    assign _5553 = _5304 == _989;
    assign _5550 = ~ _3920;
    assign _5551 = _3135 & _5550;
    assign _5554 = _5551 & _5553;
    assign _5555 = _5554 ? _4693 : _4633;
    assign _5548 = _5296 == _989;
    assign _5549 = _5293 & _5548;
    assign _5557 = _5549 ? _11940 : _5555;
    assign _5559 = _805 ? _4718 : _5557;
    assign _289 = _5559;
    always @(posedge _791) begin
        if (_789)
            _4633 <= _4718;
        else
            _4633 <= _289;
    end
    assign _5566 = _5304 == _998;
    assign _5563 = ~ _3920;
    assign _5564 = _3135 & _5563;
    assign _5567 = _5564 & _5566;
    assign _5568 = _5567 ? _4693 : _4630;
    assign _5561 = _5296 == _998;
    assign _5562 = _5293 & _5561;
    assign _5570 = _5562 ? _11940 : _5568;
    assign _5572 = _805 ? _4718 : _5570;
    assign _290 = _5572;
    always @(posedge _791) begin
        if (_789)
            _4630 <= _4718;
        else
            _4630 <= _290;
    end
    assign _5579 = _5304 == _1007;
    assign _5576 = ~ _3920;
    assign _5577 = _3135 & _5576;
    assign _5580 = _5577 & _5579;
    assign _5581 = _5580 ? _4693 : _4627;
    assign _5574 = _5296 == _1007;
    assign _5575 = _5293 & _5574;
    assign _5583 = _5575 ? _11940 : _5581;
    assign _5585 = _805 ? _4718 : _5583;
    assign _291 = _5585;
    always @(posedge _791) begin
        if (_789)
            _4627 <= _4718;
        else
            _4627 <= _291;
    end
    assign _5592 = _5304 == _1016;
    assign _5589 = ~ _3920;
    assign _5590 = _3135 & _5589;
    assign _5593 = _5590 & _5592;
    assign _5594 = _5593 ? _4693 : _4624;
    assign _5587 = _5296 == _1016;
    assign _5588 = _5293 & _5587;
    assign _5596 = _5588 ? _11940 : _5594;
    assign _5598 = _805 ? _4718 : _5596;
    assign _292 = _5598;
    always @(posedge _791) begin
        if (_789)
            _4624 <= _4718;
        else
            _4624 <= _292;
    end
    assign _5605 = _5304 == _1025;
    assign _5602 = ~ _3920;
    assign _5603 = _3135 & _5602;
    assign _5606 = _5603 & _5605;
    assign _5607 = _5606 ? _4693 : _4621;
    assign _5600 = _5296 == _1025;
    assign _5601 = _5293 & _5600;
    assign _5609 = _5601 ? _11940 : _5607;
    assign _5611 = _805 ? _4718 : _5609;
    assign _293 = _5611;
    always @(posedge _791) begin
        if (_789)
            _4621 <= _4718;
        else
            _4621 <= _293;
    end
    assign _5618 = _5304 == _1034;
    assign _5615 = ~ _3920;
    assign _5616 = _3135 & _5615;
    assign _5619 = _5616 & _5618;
    assign _5620 = _5619 ? _4693 : _4618;
    assign _5613 = _5296 == _1034;
    assign _5614 = _5293 & _5613;
    assign _5622 = _5614 ? _11940 : _5620;
    assign _5624 = _805 ? _4718 : _5622;
    assign _294 = _5624;
    always @(posedge _791) begin
        if (_789)
            _4618 <= _4718;
        else
            _4618 <= _294;
    end
    assign _5631 = _5304 == _1043;
    assign _5628 = ~ _3920;
    assign _5629 = _3135 & _5628;
    assign _5632 = _5629 & _5631;
    assign _5633 = _5632 ? _4693 : _4615;
    assign _5626 = _5296 == _1043;
    assign _5627 = _5293 & _5626;
    assign _5635 = _5627 ? _11940 : _5633;
    assign _5637 = _805 ? _4718 : _5635;
    assign _295 = _5637;
    always @(posedge _791) begin
        if (_789)
            _4615 <= _4718;
        else
            _4615 <= _295;
    end
    assign _5644 = _5304 == _1052;
    assign _5641 = ~ _3920;
    assign _5642 = _3135 & _5641;
    assign _5645 = _5642 & _5644;
    assign _5646 = _5645 ? _4693 : _4612;
    assign _5639 = _5296 == _1052;
    assign _5640 = _5293 & _5639;
    assign _5648 = _5640 ? _11940 : _5646;
    assign _5650 = _805 ? _4718 : _5648;
    assign _296 = _5650;
    always @(posedge _791) begin
        if (_789)
            _4612 <= _4718;
        else
            _4612 <= _296;
    end
    assign _5657 = _5304 == _1061;
    assign _5654 = ~ _3920;
    assign _5655 = _3135 & _5654;
    assign _5658 = _5655 & _5657;
    assign _5659 = _5658 ? _4693 : _4609;
    assign _5652 = _5296 == _1061;
    assign _5653 = _5293 & _5652;
    assign _5661 = _5653 ? _11940 : _5659;
    assign _5663 = _805 ? _4718 : _5661;
    assign _297 = _5663;
    always @(posedge _791) begin
        if (_789)
            _4609 <= _4718;
        else
            _4609 <= _297;
    end
    assign _5670 = _5304 == _1070;
    assign _5667 = ~ _3920;
    assign _5668 = _3135 & _5667;
    assign _5671 = _5668 & _5670;
    assign _5672 = _5671 ? _4693 : _4606;
    assign _5665 = _5296 == _1070;
    assign _5666 = _5293 & _5665;
    assign _5674 = _5666 ? _11940 : _5672;
    assign _5676 = _805 ? _4718 : _5674;
    assign _298 = _5676;
    always @(posedge _791) begin
        if (_789)
            _4606 <= _4718;
        else
            _4606 <= _298;
    end
    assign _5683 = _5304 == _1079;
    assign _5680 = ~ _3920;
    assign _5681 = _3135 & _5680;
    assign _5684 = _5681 & _5683;
    assign _5685 = _5684 ? _4693 : _4603;
    assign _5678 = _5296 == _1079;
    assign _5679 = _5293 & _5678;
    assign _5687 = _5679 ? _11940 : _5685;
    assign _5689 = _805 ? _4718 : _5687;
    assign _299 = _5689;
    always @(posedge _791) begin
        if (_789)
            _4603 <= _4718;
        else
            _4603 <= _299;
    end
    assign _5696 = _5304 == _1088;
    assign _5693 = ~ _3920;
    assign _5694 = _3135 & _5693;
    assign _5697 = _5694 & _5696;
    assign _5698 = _5697 ? _4693 : _4600;
    assign _5691 = _5296 == _1088;
    assign _5692 = _5293 & _5691;
    assign _5700 = _5692 ? _11940 : _5698;
    assign _5702 = _805 ? _4718 : _5700;
    assign _300 = _5702;
    always @(posedge _791) begin
        if (_789)
            _4600 <= _4718;
        else
            _4600 <= _300;
    end
    assign _5709 = _5304 == _1097;
    assign _5706 = ~ _3920;
    assign _5707 = _3135 & _5706;
    assign _5710 = _5707 & _5709;
    assign _5711 = _5710 ? _4693 : _4597;
    assign _5704 = _5296 == _1097;
    assign _5705 = _5293 & _5704;
    assign _5713 = _5705 ? _11940 : _5711;
    assign _5715 = _805 ? _4718 : _5713;
    assign _301 = _5715;
    always @(posedge _791) begin
        if (_789)
            _4597 <= _4718;
        else
            _4597 <= _301;
    end
    assign _5722 = _5304 == _1106;
    assign _5719 = ~ _3920;
    assign _5720 = _3135 & _5719;
    assign _5723 = _5720 & _5722;
    assign _5724 = _5723 ? _4693 : _4594;
    assign _5717 = _5296 == _1106;
    assign _5718 = _5293 & _5717;
    assign _5726 = _5718 ? _11940 : _5724;
    assign _5728 = _805 ? _4718 : _5726;
    assign _302 = _5728;
    always @(posedge _791) begin
        if (_789)
            _4594 <= _4718;
        else
            _4594 <= _302;
    end
    assign _5735 = _5304 == _1115;
    assign _5732 = ~ _3920;
    assign _5733 = _3135 & _5732;
    assign _5736 = _5733 & _5735;
    assign _5737 = _5736 ? _4693 : _4591;
    assign _5730 = _5296 == _1115;
    assign _5731 = _5293 & _5730;
    assign _5739 = _5731 ? _11940 : _5737;
    assign _5741 = _805 ? _4718 : _5739;
    assign _303 = _5741;
    always @(posedge _791) begin
        if (_789)
            _4591 <= _4718;
        else
            _4591 <= _303;
    end
    assign _5748 = _5304 == _1124;
    assign _5745 = ~ _3920;
    assign _5746 = _3135 & _5745;
    assign _5749 = _5746 & _5748;
    assign _5750 = _5749 ? _4693 : _4588;
    assign _5743 = _5296 == _1124;
    assign _5744 = _5293 & _5743;
    assign _5752 = _5744 ? _11940 : _5750;
    assign _5754 = _805 ? _4718 : _5752;
    assign _304 = _5754;
    always @(posedge _791) begin
        if (_789)
            _4588 <= _4718;
        else
            _4588 <= _304;
    end
    assign _5761 = _5304 == _1133;
    assign _5758 = ~ _3920;
    assign _5759 = _3135 & _5758;
    assign _5762 = _5759 & _5761;
    assign _5763 = _5762 ? _4693 : _4585;
    assign _5756 = _5296 == _1133;
    assign _5757 = _5293 & _5756;
    assign _5765 = _5757 ? _11940 : _5763;
    assign _5767 = _805 ? _4718 : _5765;
    assign _305 = _5767;
    always @(posedge _791) begin
        if (_789)
            _4585 <= _4718;
        else
            _4585 <= _305;
    end
    assign _5774 = _5304 == _1142;
    assign _5771 = ~ _3920;
    assign _5772 = _3135 & _5771;
    assign _5775 = _5772 & _5774;
    assign _5776 = _5775 ? _4693 : _4582;
    assign _5769 = _5296 == _1142;
    assign _5770 = _5293 & _5769;
    assign _5778 = _5770 ? _11940 : _5776;
    assign _5780 = _805 ? _4718 : _5778;
    assign _306 = _5780;
    always @(posedge _791) begin
        if (_789)
            _4582 <= _4718;
        else
            _4582 <= _306;
    end
    assign _5787 = _5304 == _1151;
    assign _5784 = ~ _3920;
    assign _5785 = _3135 & _5784;
    assign _5788 = _5785 & _5787;
    assign _5789 = _5788 ? _4693 : _4579;
    assign _5782 = _5296 == _1151;
    assign _5783 = _5293 & _5782;
    assign _5791 = _5783 ? _11940 : _5789;
    assign _5793 = _805 ? _4718 : _5791;
    assign _307 = _5793;
    always @(posedge _791) begin
        if (_789)
            _4579 <= _4718;
        else
            _4579 <= _307;
    end
    assign _5800 = _5304 == _1160;
    assign _5797 = ~ _3920;
    assign _5798 = _3135 & _5797;
    assign _5801 = _5798 & _5800;
    assign _5802 = _5801 ? _4693 : _4576;
    assign _5795 = _5296 == _1160;
    assign _5796 = _5293 & _5795;
    assign _5804 = _5796 ? _11940 : _5802;
    assign _5806 = _805 ? _4718 : _5804;
    assign _308 = _5806;
    always @(posedge _791) begin
        if (_789)
            _4576 <= _4718;
        else
            _4576 <= _308;
    end
    assign _5813 = _5304 == _1169;
    assign _5810 = ~ _3920;
    assign _5811 = _3135 & _5810;
    assign _5814 = _5811 & _5813;
    assign _5815 = _5814 ? _4693 : _4573;
    assign _5808 = _5296 == _1169;
    assign _5809 = _5293 & _5808;
    assign _5817 = _5809 ? _11940 : _5815;
    assign _5819 = _805 ? _4718 : _5817;
    assign _309 = _5819;
    always @(posedge _791) begin
        if (_789)
            _4573 <= _4718;
        else
            _4573 <= _309;
    end
    assign _5826 = _5304 == _1178;
    assign _5823 = ~ _3920;
    assign _5824 = _3135 & _5823;
    assign _5827 = _5824 & _5826;
    assign _5828 = _5827 ? _4693 : _4570;
    assign _5821 = _5296 == _1178;
    assign _5822 = _5293 & _5821;
    assign _5830 = _5822 ? _11940 : _5828;
    assign _5832 = _805 ? _4718 : _5830;
    assign _310 = _5832;
    always @(posedge _791) begin
        if (_789)
            _4570 <= _4718;
        else
            _4570 <= _310;
    end
    assign _5839 = _5304 == _1187;
    assign _5836 = ~ _3920;
    assign _5837 = _3135 & _5836;
    assign _5840 = _5837 & _5839;
    assign _5841 = _5840 ? _4693 : _4567;
    assign _5834 = _5296 == _1187;
    assign _5835 = _5293 & _5834;
    assign _5843 = _5835 ? _11940 : _5841;
    assign _5845 = _805 ? _4718 : _5843;
    assign _311 = _5845;
    always @(posedge _791) begin
        if (_789)
            _4567 <= _4718;
        else
            _4567 <= _311;
    end
    assign _5852 = _5304 == _1196;
    assign _5849 = ~ _3920;
    assign _5850 = _3135 & _5849;
    assign _5853 = _5850 & _5852;
    assign _5854 = _5853 ? _4693 : _4564;
    assign _5847 = _5296 == _1196;
    assign _5848 = _5293 & _5847;
    assign _5856 = _5848 ? _11940 : _5854;
    assign _5858 = _805 ? _4718 : _5856;
    assign _312 = _5858;
    always @(posedge _791) begin
        if (_789)
            _4564 <= _4718;
        else
            _4564 <= _312;
    end
    assign _5865 = _5304 == _1205;
    assign _5862 = ~ _3920;
    assign _5863 = _3135 & _5862;
    assign _5866 = _5863 & _5865;
    assign _5867 = _5866 ? _4693 : _4561;
    assign _5860 = _5296 == _1205;
    assign _5861 = _5293 & _5860;
    assign _5869 = _5861 ? _11940 : _5867;
    assign _5871 = _805 ? _4718 : _5869;
    assign _313 = _5871;
    always @(posedge _791) begin
        if (_789)
            _4561 <= _4718;
        else
            _4561 <= _313;
    end
    assign _5878 = _5304 == _1214;
    assign _5875 = ~ _3920;
    assign _5876 = _3135 & _5875;
    assign _5879 = _5876 & _5878;
    assign _5880 = _5879 ? _4693 : _4558;
    assign _5873 = _5296 == _1214;
    assign _5874 = _5293 & _5873;
    assign _5882 = _5874 ? _11940 : _5880;
    assign _5884 = _805 ? _4718 : _5882;
    assign _314 = _5884;
    always @(posedge _791) begin
        if (_789)
            _4558 <= _4718;
        else
            _4558 <= _314;
    end
    assign _5891 = _5304 == _1223;
    assign _5888 = ~ _3920;
    assign _5889 = _3135 & _5888;
    assign _5892 = _5889 & _5891;
    assign _5893 = _5892 ? _4693 : _4555;
    assign _5886 = _5296 == _1223;
    assign _5887 = _5293 & _5886;
    assign _5895 = _5887 ? _11940 : _5893;
    assign _5897 = _805 ? _4718 : _5895;
    assign _315 = _5897;
    always @(posedge _791) begin
        if (_789)
            _4555 <= _4718;
        else
            _4555 <= _315;
    end
    assign _5904 = _5304 == _1232;
    assign _5901 = ~ _3920;
    assign _5902 = _3135 & _5901;
    assign _5905 = _5902 & _5904;
    assign _5906 = _5905 ? _4693 : _4552;
    assign _5899 = _5296 == _1232;
    assign _5900 = _5293 & _5899;
    assign _5908 = _5900 ? _11940 : _5906;
    assign _5910 = _805 ? _4718 : _5908;
    assign _316 = _5910;
    always @(posedge _791) begin
        if (_789)
            _4552 <= _4718;
        else
            _4552 <= _316;
    end
    assign _5917 = _5304 == _1241;
    assign _5914 = ~ _3920;
    assign _5915 = _3135 & _5914;
    assign _5918 = _5915 & _5917;
    assign _5919 = _5918 ? _4693 : _4549;
    assign _5912 = _5296 == _1241;
    assign _5913 = _5293 & _5912;
    assign _5921 = _5913 ? _11940 : _5919;
    assign _5923 = _805 ? _4718 : _5921;
    assign _317 = _5923;
    always @(posedge _791) begin
        if (_789)
            _4549 <= _4718;
        else
            _4549 <= _317;
    end
    assign _5930 = _5304 == _1250;
    assign _5927 = ~ _3920;
    assign _5928 = _3135 & _5927;
    assign _5931 = _5928 & _5930;
    assign _5932 = _5931 ? _4693 : _4546;
    assign _5925 = _5296 == _1250;
    assign _5926 = _5293 & _5925;
    assign _5934 = _5926 ? _11940 : _5932;
    assign _5936 = _805 ? _4718 : _5934;
    assign _318 = _5936;
    always @(posedge _791) begin
        if (_789)
            _4546 <= _4718;
        else
            _4546 <= _318;
    end
    assign _5943 = _5304 == _1259;
    assign _5940 = ~ _3920;
    assign _5941 = _3135 & _5940;
    assign _5944 = _5941 & _5943;
    assign _5945 = _5944 ? _4693 : _4543;
    assign _5938 = _5296 == _1259;
    assign _5939 = _5293 & _5938;
    assign _5947 = _5939 ? _11940 : _5945;
    assign _5949 = _805 ? _4718 : _5947;
    assign _319 = _5949;
    always @(posedge _791) begin
        if (_789)
            _4543 <= _4718;
        else
            _4543 <= _319;
    end
    assign _5956 = _5304 == _1268;
    assign _5953 = ~ _3920;
    assign _5954 = _3135 & _5953;
    assign _5957 = _5954 & _5956;
    assign _5958 = _5957 ? _4693 : _4540;
    assign _5951 = _5296 == _1268;
    assign _5952 = _5293 & _5951;
    assign _5960 = _5952 ? _11940 : _5958;
    assign _5962 = _805 ? _4718 : _5960;
    assign _320 = _5962;
    always @(posedge _791) begin
        if (_789)
            _4540 <= _4718;
        else
            _4540 <= _320;
    end
    assign _5969 = _5304 == _1277;
    assign _5966 = ~ _3920;
    assign _5967 = _3135 & _5966;
    assign _5970 = _5967 & _5969;
    assign _5971 = _5970 ? _4693 : _4537;
    assign _5964 = _5296 == _1277;
    assign _5965 = _5293 & _5964;
    assign _5973 = _5965 ? _11940 : _5971;
    assign _5975 = _805 ? _4718 : _5973;
    assign _321 = _5975;
    always @(posedge _791) begin
        if (_789)
            _4537 <= _4718;
        else
            _4537 <= _321;
    end
    assign _5982 = _5304 == _1286;
    assign _5979 = ~ _3920;
    assign _5980 = _3135 & _5979;
    assign _5983 = _5980 & _5982;
    assign _5984 = _5983 ? _4693 : _4534;
    assign _5977 = _5296 == _1286;
    assign _5978 = _5293 & _5977;
    assign _5986 = _5978 ? _11940 : _5984;
    assign _5988 = _805 ? _4718 : _5986;
    assign _322 = _5988;
    always @(posedge _791) begin
        if (_789)
            _4534 <= _4718;
        else
            _4534 <= _322;
    end
    assign _5995 = _5304 == _1295;
    assign _5992 = ~ _3920;
    assign _5993 = _3135 & _5992;
    assign _5996 = _5993 & _5995;
    assign _5997 = _5996 ? _4693 : _4531;
    assign _5990 = _5296 == _1295;
    assign _5991 = _5293 & _5990;
    assign _5999 = _5991 ? _11940 : _5997;
    assign _6001 = _805 ? _4718 : _5999;
    assign _323 = _6001;
    always @(posedge _791) begin
        if (_789)
            _4531 <= _4718;
        else
            _4531 <= _323;
    end
    assign _6008 = _5304 == _1304;
    assign _6005 = ~ _3920;
    assign _6006 = _3135 & _6005;
    assign _6009 = _6006 & _6008;
    assign _6010 = _6009 ? _4693 : _4528;
    assign _6003 = _5296 == _1304;
    assign _6004 = _5293 & _6003;
    assign _6012 = _6004 ? _11940 : _6010;
    assign _6014 = _805 ? _4718 : _6012;
    assign _324 = _6014;
    always @(posedge _791) begin
        if (_789)
            _4528 <= _4718;
        else
            _4528 <= _324;
    end
    assign _6021 = _5304 == _1313;
    assign _6018 = ~ _3920;
    assign _6019 = _3135 & _6018;
    assign _6022 = _6019 & _6021;
    assign _6023 = _6022 ? _4693 : _4525;
    assign _6016 = _5296 == _1313;
    assign _6017 = _5293 & _6016;
    assign _6025 = _6017 ? _11940 : _6023;
    assign _6027 = _805 ? _4718 : _6025;
    assign _325 = _6027;
    always @(posedge _791) begin
        if (_789)
            _4525 <= _4718;
        else
            _4525 <= _325;
    end
    assign _6034 = _5304 == _1322;
    assign _6031 = ~ _3920;
    assign _6032 = _3135 & _6031;
    assign _6035 = _6032 & _6034;
    assign _6036 = _6035 ? _4693 : _4522;
    assign _6029 = _5296 == _1322;
    assign _6030 = _5293 & _6029;
    assign _6038 = _6030 ? _11940 : _6036;
    assign _6040 = _805 ? _4718 : _6038;
    assign _326 = _6040;
    always @(posedge _791) begin
        if (_789)
            _4522 <= _4718;
        else
            _4522 <= _326;
    end
    assign _6047 = _5304 == _1331;
    assign _6044 = ~ _3920;
    assign _6045 = _3135 & _6044;
    assign _6048 = _6045 & _6047;
    assign _6049 = _6048 ? _4693 : _4519;
    assign _6042 = _5296 == _1331;
    assign _6043 = _5293 & _6042;
    assign _6051 = _6043 ? _11940 : _6049;
    assign _6053 = _805 ? _4718 : _6051;
    assign _327 = _6053;
    always @(posedge _791) begin
        if (_789)
            _4519 <= _4718;
        else
            _4519 <= _327;
    end
    assign _6060 = _5304 == _1340;
    assign _6057 = ~ _3920;
    assign _6058 = _3135 & _6057;
    assign _6061 = _6058 & _6060;
    assign _6062 = _6061 ? _4693 : _4516;
    assign _6055 = _5296 == _1340;
    assign _6056 = _5293 & _6055;
    assign _6064 = _6056 ? _11940 : _6062;
    assign _6066 = _805 ? _4718 : _6064;
    assign _328 = _6066;
    always @(posedge _791) begin
        if (_789)
            _4516 <= _4718;
        else
            _4516 <= _328;
    end
    assign _6073 = _5304 == _1349;
    assign _6070 = ~ _3920;
    assign _6071 = _3135 & _6070;
    assign _6074 = _6071 & _6073;
    assign _6075 = _6074 ? _4693 : _4513;
    assign _6068 = _5296 == _1349;
    assign _6069 = _5293 & _6068;
    assign _6077 = _6069 ? _11940 : _6075;
    assign _6079 = _805 ? _4718 : _6077;
    assign _329 = _6079;
    always @(posedge _791) begin
        if (_789)
            _4513 <= _4718;
        else
            _4513 <= _329;
    end
    assign _6086 = _5304 == _1358;
    assign _6083 = ~ _3920;
    assign _6084 = _3135 & _6083;
    assign _6087 = _6084 & _6086;
    assign _6088 = _6087 ? _4693 : _4510;
    assign _6081 = _5296 == _1358;
    assign _6082 = _5293 & _6081;
    assign _6090 = _6082 ? _11940 : _6088;
    assign _6092 = _805 ? _4718 : _6090;
    assign _330 = _6092;
    always @(posedge _791) begin
        if (_789)
            _4510 <= _4718;
        else
            _4510 <= _330;
    end
    assign _6099 = _5304 == _1367;
    assign _6096 = ~ _3920;
    assign _6097 = _3135 & _6096;
    assign _6100 = _6097 & _6099;
    assign _6101 = _6100 ? _4693 : _4507;
    assign _6094 = _5296 == _1367;
    assign _6095 = _5293 & _6094;
    assign _6103 = _6095 ? _11940 : _6101;
    assign _6105 = _805 ? _4718 : _6103;
    assign _331 = _6105;
    always @(posedge _791) begin
        if (_789)
            _4507 <= _4718;
        else
            _4507 <= _331;
    end
    assign _6112 = _5304 == _1376;
    assign _6109 = ~ _3920;
    assign _6110 = _3135 & _6109;
    assign _6113 = _6110 & _6112;
    assign _6114 = _6113 ? _4693 : _4504;
    assign _6107 = _5296 == _1376;
    assign _6108 = _5293 & _6107;
    assign _6116 = _6108 ? _11940 : _6114;
    assign _6118 = _805 ? _4718 : _6116;
    assign _332 = _6118;
    always @(posedge _791) begin
        if (_789)
            _4504 <= _4718;
        else
            _4504 <= _332;
    end
    assign _6125 = _5304 == _1385;
    assign _6122 = ~ _3920;
    assign _6123 = _3135 & _6122;
    assign _6126 = _6123 & _6125;
    assign _6127 = _6126 ? _4693 : _4501;
    assign _6120 = _5296 == _1385;
    assign _6121 = _5293 & _6120;
    assign _6129 = _6121 ? _11940 : _6127;
    assign _6131 = _805 ? _4718 : _6129;
    assign _333 = _6131;
    always @(posedge _791) begin
        if (_789)
            _4501 <= _4718;
        else
            _4501 <= _333;
    end
    assign _6138 = _5304 == _1394;
    assign _6135 = ~ _3920;
    assign _6136 = _3135 & _6135;
    assign _6139 = _6136 & _6138;
    assign _6140 = _6139 ? _4693 : _4498;
    assign _6133 = _5296 == _1394;
    assign _6134 = _5293 & _6133;
    assign _6142 = _6134 ? _11940 : _6140;
    assign _6144 = _805 ? _4718 : _6142;
    assign _334 = _6144;
    always @(posedge _791) begin
        if (_789)
            _4498 <= _4718;
        else
            _4498 <= _334;
    end
    assign _6151 = _5304 == _1403;
    assign _6148 = ~ _3920;
    assign _6149 = _3135 & _6148;
    assign _6152 = _6149 & _6151;
    assign _6153 = _6152 ? _4693 : _4495;
    assign _6146 = _5296 == _1403;
    assign _6147 = _5293 & _6146;
    assign _6155 = _6147 ? _11940 : _6153;
    assign _6157 = _805 ? _4718 : _6155;
    assign _335 = _6157;
    always @(posedge _791) begin
        if (_789)
            _4495 <= _4718;
        else
            _4495 <= _335;
    end
    assign _6164 = _5304 == _1412;
    assign _6161 = ~ _3920;
    assign _6162 = _3135 & _6161;
    assign _6165 = _6162 & _6164;
    assign _6166 = _6165 ? _4693 : _4492;
    assign _6159 = _5296 == _1412;
    assign _6160 = _5293 & _6159;
    assign _6168 = _6160 ? _11940 : _6166;
    assign _6170 = _805 ? _4718 : _6168;
    assign _336 = _6170;
    always @(posedge _791) begin
        if (_789)
            _4492 <= _4718;
        else
            _4492 <= _336;
    end
    assign _6177 = _5304 == _1421;
    assign _6174 = ~ _3920;
    assign _6175 = _3135 & _6174;
    assign _6178 = _6175 & _6177;
    assign _6179 = _6178 ? _4693 : _4489;
    assign _6172 = _5296 == _1421;
    assign _6173 = _5293 & _6172;
    assign _6181 = _6173 ? _11940 : _6179;
    assign _6183 = _805 ? _4718 : _6181;
    assign _337 = _6183;
    always @(posedge _791) begin
        if (_789)
            _4489 <= _4718;
        else
            _4489 <= _337;
    end
    assign _6190 = _5304 == _1430;
    assign _6187 = ~ _3920;
    assign _6188 = _3135 & _6187;
    assign _6191 = _6188 & _6190;
    assign _6192 = _6191 ? _4693 : _4486;
    assign _6185 = _5296 == _1430;
    assign _6186 = _5293 & _6185;
    assign _6194 = _6186 ? _11940 : _6192;
    assign _6196 = _805 ? _4718 : _6194;
    assign _338 = _6196;
    always @(posedge _791) begin
        if (_789)
            _4486 <= _4718;
        else
            _4486 <= _338;
    end
    assign _6203 = _5304 == _1439;
    assign _6200 = ~ _3920;
    assign _6201 = _3135 & _6200;
    assign _6204 = _6201 & _6203;
    assign _6205 = _6204 ? _4693 : _4483;
    assign _6198 = _5296 == _1439;
    assign _6199 = _5293 & _6198;
    assign _6207 = _6199 ? _11940 : _6205;
    assign _6209 = _805 ? _4718 : _6207;
    assign _339 = _6209;
    always @(posedge _791) begin
        if (_789)
            _4483 <= _4718;
        else
            _4483 <= _339;
    end
    assign _6216 = _5304 == _1448;
    assign _6213 = ~ _3920;
    assign _6214 = _3135 & _6213;
    assign _6217 = _6214 & _6216;
    assign _6218 = _6217 ? _4693 : _4480;
    assign _6211 = _5296 == _1448;
    assign _6212 = _5293 & _6211;
    assign _6220 = _6212 ? _11940 : _6218;
    assign _6222 = _805 ? _4718 : _6220;
    assign _340 = _6222;
    always @(posedge _791) begin
        if (_789)
            _4480 <= _4718;
        else
            _4480 <= _340;
    end
    assign _6229 = _5304 == _1457;
    assign _6226 = ~ _3920;
    assign _6227 = _3135 & _6226;
    assign _6230 = _6227 & _6229;
    assign _6231 = _6230 ? _4693 : _4477;
    assign _6224 = _5296 == _1457;
    assign _6225 = _5293 & _6224;
    assign _6233 = _6225 ? _11940 : _6231;
    assign _6235 = _805 ? _4718 : _6233;
    assign _341 = _6235;
    always @(posedge _791) begin
        if (_789)
            _4477 <= _4718;
        else
            _4477 <= _341;
    end
    assign _6242 = _5304 == _1466;
    assign _6239 = ~ _3920;
    assign _6240 = _3135 & _6239;
    assign _6243 = _6240 & _6242;
    assign _6244 = _6243 ? _4693 : _4474;
    assign _6237 = _5296 == _1466;
    assign _6238 = _5293 & _6237;
    assign _6246 = _6238 ? _11940 : _6244;
    assign _6248 = _805 ? _4718 : _6246;
    assign _342 = _6248;
    always @(posedge _791) begin
        if (_789)
            _4474 <= _4718;
        else
            _4474 <= _342;
    end
    assign _6255 = _5304 == _1475;
    assign _6252 = ~ _3920;
    assign _6253 = _3135 & _6252;
    assign _6256 = _6253 & _6255;
    assign _6257 = _6256 ? _4693 : _4471;
    assign _6250 = _5296 == _1475;
    assign _6251 = _5293 & _6250;
    assign _6259 = _6251 ? _11940 : _6257;
    assign _6261 = _805 ? _4718 : _6259;
    assign _343 = _6261;
    always @(posedge _791) begin
        if (_789)
            _4471 <= _4718;
        else
            _4471 <= _343;
    end
    assign _6268 = _5304 == _1484;
    assign _6265 = ~ _3920;
    assign _6266 = _3135 & _6265;
    assign _6269 = _6266 & _6268;
    assign _6270 = _6269 ? _4693 : _4468;
    assign _6263 = _5296 == _1484;
    assign _6264 = _5293 & _6263;
    assign _6272 = _6264 ? _11940 : _6270;
    assign _6274 = _805 ? _4718 : _6272;
    assign _344 = _6274;
    always @(posedge _791) begin
        if (_789)
            _4468 <= _4718;
        else
            _4468 <= _344;
    end
    assign _6281 = _5304 == _1493;
    assign _6278 = ~ _3920;
    assign _6279 = _3135 & _6278;
    assign _6282 = _6279 & _6281;
    assign _6283 = _6282 ? _4693 : _4465;
    assign _6276 = _5296 == _1493;
    assign _6277 = _5293 & _6276;
    assign _6285 = _6277 ? _11940 : _6283;
    assign _6287 = _805 ? _4718 : _6285;
    assign _345 = _6287;
    always @(posedge _791) begin
        if (_789)
            _4465 <= _4718;
        else
            _4465 <= _345;
    end
    assign _6294 = _5304 == _1502;
    assign _6291 = ~ _3920;
    assign _6292 = _3135 & _6291;
    assign _6295 = _6292 & _6294;
    assign _6296 = _6295 ? _4693 : _4462;
    assign _6289 = _5296 == _1502;
    assign _6290 = _5293 & _6289;
    assign _6298 = _6290 ? _11940 : _6296;
    assign _6300 = _805 ? _4718 : _6298;
    assign _346 = _6300;
    always @(posedge _791) begin
        if (_789)
            _4462 <= _4718;
        else
            _4462 <= _346;
    end
    assign _6307 = _5304 == _1511;
    assign _6304 = ~ _3920;
    assign _6305 = _3135 & _6304;
    assign _6308 = _6305 & _6307;
    assign _6309 = _6308 ? _4693 : _4459;
    assign _6302 = _5296 == _1511;
    assign _6303 = _5293 & _6302;
    assign _6311 = _6303 ? _11940 : _6309;
    assign _6313 = _805 ? _4718 : _6311;
    assign _347 = _6313;
    always @(posedge _791) begin
        if (_789)
            _4459 <= _4718;
        else
            _4459 <= _347;
    end
    assign _6320 = _5304 == _1520;
    assign _6317 = ~ _3920;
    assign _6318 = _3135 & _6317;
    assign _6321 = _6318 & _6320;
    assign _6322 = _6321 ? _4693 : _4456;
    assign _6315 = _5296 == _1520;
    assign _6316 = _5293 & _6315;
    assign _6324 = _6316 ? _11940 : _6322;
    assign _6326 = _805 ? _4718 : _6324;
    assign _348 = _6326;
    always @(posedge _791) begin
        if (_789)
            _4456 <= _4718;
        else
            _4456 <= _348;
    end
    assign _6333 = _5304 == _1529;
    assign _6330 = ~ _3920;
    assign _6331 = _3135 & _6330;
    assign _6334 = _6331 & _6333;
    assign _6335 = _6334 ? _4693 : _4453;
    assign _6328 = _5296 == _1529;
    assign _6329 = _5293 & _6328;
    assign _6337 = _6329 ? _11940 : _6335;
    assign _6339 = _805 ? _4718 : _6337;
    assign _349 = _6339;
    always @(posedge _791) begin
        if (_789)
            _4453 <= _4718;
        else
            _4453 <= _349;
    end
    assign _6346 = _5304 == _1538;
    assign _6343 = ~ _3920;
    assign _6344 = _3135 & _6343;
    assign _6347 = _6344 & _6346;
    assign _6348 = _6347 ? _4693 : _4450;
    assign _6341 = _5296 == _1538;
    assign _6342 = _5293 & _6341;
    assign _6350 = _6342 ? _11940 : _6348;
    assign _6352 = _805 ? _4718 : _6350;
    assign _350 = _6352;
    always @(posedge _791) begin
        if (_789)
            _4450 <= _4718;
        else
            _4450 <= _350;
    end
    assign _6359 = _5304 == _1547;
    assign _6356 = ~ _3920;
    assign _6357 = _3135 & _6356;
    assign _6360 = _6357 & _6359;
    assign _6361 = _6360 ? _4693 : _4447;
    assign _6354 = _5296 == _1547;
    assign _6355 = _5293 & _6354;
    assign _6363 = _6355 ? _11940 : _6361;
    assign _6365 = _805 ? _4718 : _6363;
    assign _351 = _6365;
    always @(posedge _791) begin
        if (_789)
            _4447 <= _4718;
        else
            _4447 <= _351;
    end
    assign _6372 = _5304 == _1556;
    assign _6369 = ~ _3920;
    assign _6370 = _3135 & _6369;
    assign _6373 = _6370 & _6372;
    assign _6374 = _6373 ? _4693 : _4444;
    assign _6367 = _5296 == _1556;
    assign _6368 = _5293 & _6367;
    assign _6376 = _6368 ? _11940 : _6374;
    assign _6378 = _805 ? _4718 : _6376;
    assign _352 = _6378;
    always @(posedge _791) begin
        if (_789)
            _4444 <= _4718;
        else
            _4444 <= _352;
    end
    assign _6385 = _5304 == _1565;
    assign _6382 = ~ _3920;
    assign _6383 = _3135 & _6382;
    assign _6386 = _6383 & _6385;
    assign _6387 = _6386 ? _4693 : _4441;
    assign _6380 = _5296 == _1565;
    assign _6381 = _5293 & _6380;
    assign _6389 = _6381 ? _11940 : _6387;
    assign _6391 = _805 ? _4718 : _6389;
    assign _353 = _6391;
    always @(posedge _791) begin
        if (_789)
            _4441 <= _4718;
        else
            _4441 <= _353;
    end
    assign _6398 = _5304 == _1574;
    assign _6395 = ~ _3920;
    assign _6396 = _3135 & _6395;
    assign _6399 = _6396 & _6398;
    assign _6400 = _6399 ? _4693 : _4438;
    assign _6393 = _5296 == _1574;
    assign _6394 = _5293 & _6393;
    assign _6402 = _6394 ? _11940 : _6400;
    assign _6404 = _805 ? _4718 : _6402;
    assign _354 = _6404;
    always @(posedge _791) begin
        if (_789)
            _4438 <= _4718;
        else
            _4438 <= _354;
    end
    assign _6411 = _5304 == _1583;
    assign _6408 = ~ _3920;
    assign _6409 = _3135 & _6408;
    assign _6412 = _6409 & _6411;
    assign _6413 = _6412 ? _4693 : _4435;
    assign _6406 = _5296 == _1583;
    assign _6407 = _5293 & _6406;
    assign _6415 = _6407 ? _11940 : _6413;
    assign _6417 = _805 ? _4718 : _6415;
    assign _355 = _6417;
    always @(posedge _791) begin
        if (_789)
            _4435 <= _4718;
        else
            _4435 <= _355;
    end
    assign _6424 = _5304 == _1592;
    assign _6421 = ~ _3920;
    assign _6422 = _3135 & _6421;
    assign _6425 = _6422 & _6424;
    assign _6426 = _6425 ? _4693 : _4432;
    assign _6419 = _5296 == _1592;
    assign _6420 = _5293 & _6419;
    assign _6428 = _6420 ? _11940 : _6426;
    assign _6430 = _805 ? _4718 : _6428;
    assign _356 = _6430;
    always @(posedge _791) begin
        if (_789)
            _4432 <= _4718;
        else
            _4432 <= _356;
    end
    assign _6437 = _5304 == _1601;
    assign _6434 = ~ _3920;
    assign _6435 = _3135 & _6434;
    assign _6438 = _6435 & _6437;
    assign _6439 = _6438 ? _4693 : _4429;
    assign _6432 = _5296 == _1601;
    assign _6433 = _5293 & _6432;
    assign _6441 = _6433 ? _11940 : _6439;
    assign _6443 = _805 ? _4718 : _6441;
    assign _357 = _6443;
    always @(posedge _791) begin
        if (_789)
            _4429 <= _4718;
        else
            _4429 <= _357;
    end
    assign _6450 = _5304 == _1610;
    assign _6447 = ~ _3920;
    assign _6448 = _3135 & _6447;
    assign _6451 = _6448 & _6450;
    assign _6452 = _6451 ? _4693 : _4426;
    assign _6445 = _5296 == _1610;
    assign _6446 = _5293 & _6445;
    assign _6454 = _6446 ? _11940 : _6452;
    assign _6456 = _805 ? _4718 : _6454;
    assign _358 = _6456;
    always @(posedge _791) begin
        if (_789)
            _4426 <= _4718;
        else
            _4426 <= _358;
    end
    assign _6463 = _5304 == _1619;
    assign _6460 = ~ _3920;
    assign _6461 = _3135 & _6460;
    assign _6464 = _6461 & _6463;
    assign _6465 = _6464 ? _4693 : _4423;
    assign _6458 = _5296 == _1619;
    assign _6459 = _5293 & _6458;
    assign _6467 = _6459 ? _11940 : _6465;
    assign _6469 = _805 ? _4718 : _6467;
    assign _359 = _6469;
    always @(posedge _791) begin
        if (_789)
            _4423 <= _4718;
        else
            _4423 <= _359;
    end
    assign _6476 = _5304 == _1628;
    assign _6473 = ~ _3920;
    assign _6474 = _3135 & _6473;
    assign _6477 = _6474 & _6476;
    assign _6478 = _6477 ? _4693 : _4420;
    assign _6471 = _5296 == _1628;
    assign _6472 = _5293 & _6471;
    assign _6480 = _6472 ? _11940 : _6478;
    assign _6482 = _805 ? _4718 : _6480;
    assign _360 = _6482;
    always @(posedge _791) begin
        if (_789)
            _4420 <= _4718;
        else
            _4420 <= _360;
    end
    assign _6489 = _5304 == _1637;
    assign _6486 = ~ _3920;
    assign _6487 = _3135 & _6486;
    assign _6490 = _6487 & _6489;
    assign _6491 = _6490 ? _4693 : _4417;
    assign _6484 = _5296 == _1637;
    assign _6485 = _5293 & _6484;
    assign _6493 = _6485 ? _11940 : _6491;
    assign _6495 = _805 ? _4718 : _6493;
    assign _361 = _6495;
    always @(posedge _791) begin
        if (_789)
            _4417 <= _4718;
        else
            _4417 <= _361;
    end
    assign _6502 = _5304 == _1646;
    assign _6499 = ~ _3920;
    assign _6500 = _3135 & _6499;
    assign _6503 = _6500 & _6502;
    assign _6504 = _6503 ? _4693 : _4414;
    assign _6497 = _5296 == _1646;
    assign _6498 = _5293 & _6497;
    assign _6506 = _6498 ? _11940 : _6504;
    assign _6508 = _805 ? _4718 : _6506;
    assign _362 = _6508;
    always @(posedge _791) begin
        if (_789)
            _4414 <= _4718;
        else
            _4414 <= _362;
    end
    assign _6515 = _5304 == _1655;
    assign _6512 = ~ _3920;
    assign _6513 = _3135 & _6512;
    assign _6516 = _6513 & _6515;
    assign _6517 = _6516 ? _4693 : _4411;
    assign _6510 = _5296 == _1655;
    assign _6511 = _5293 & _6510;
    assign _6519 = _6511 ? _11940 : _6517;
    assign _6521 = _805 ? _4718 : _6519;
    assign _363 = _6521;
    always @(posedge _791) begin
        if (_789)
            _4411 <= _4718;
        else
            _4411 <= _363;
    end
    assign _6528 = _5304 == _1664;
    assign _6525 = ~ _3920;
    assign _6526 = _3135 & _6525;
    assign _6529 = _6526 & _6528;
    assign _6530 = _6529 ? _4693 : _4408;
    assign _6523 = _5296 == _1664;
    assign _6524 = _5293 & _6523;
    assign _6532 = _6524 ? _11940 : _6530;
    assign _6534 = _805 ? _4718 : _6532;
    assign _364 = _6534;
    always @(posedge _791) begin
        if (_789)
            _4408 <= _4718;
        else
            _4408 <= _364;
    end
    assign _6541 = _5304 == _1673;
    assign _6538 = ~ _3920;
    assign _6539 = _3135 & _6538;
    assign _6542 = _6539 & _6541;
    assign _6543 = _6542 ? _4693 : _4405;
    assign _6536 = _5296 == _1673;
    assign _6537 = _5293 & _6536;
    assign _6545 = _6537 ? _11940 : _6543;
    assign _6547 = _805 ? _4718 : _6545;
    assign _365 = _6547;
    always @(posedge _791) begin
        if (_789)
            _4405 <= _4718;
        else
            _4405 <= _365;
    end
    assign _6554 = _5304 == _1682;
    assign _6551 = ~ _3920;
    assign _6552 = _3135 & _6551;
    assign _6555 = _6552 & _6554;
    assign _6556 = _6555 ? _4693 : _4402;
    assign _6549 = _5296 == _1682;
    assign _6550 = _5293 & _6549;
    assign _6558 = _6550 ? _11940 : _6556;
    assign _6560 = _805 ? _4718 : _6558;
    assign _366 = _6560;
    always @(posedge _791) begin
        if (_789)
            _4402 <= _4718;
        else
            _4402 <= _366;
    end
    assign _6567 = _5304 == _1691;
    assign _6564 = ~ _3920;
    assign _6565 = _3135 & _6564;
    assign _6568 = _6565 & _6567;
    assign _6569 = _6568 ? _4693 : _4399;
    assign _6562 = _5296 == _1691;
    assign _6563 = _5293 & _6562;
    assign _6571 = _6563 ? _11940 : _6569;
    assign _6573 = _805 ? _4718 : _6571;
    assign _367 = _6573;
    always @(posedge _791) begin
        if (_789)
            _4399 <= _4718;
        else
            _4399 <= _367;
    end
    assign _6580 = _5304 == _1700;
    assign _6577 = ~ _3920;
    assign _6578 = _3135 & _6577;
    assign _6581 = _6578 & _6580;
    assign _6582 = _6581 ? _4693 : _4396;
    assign _6575 = _5296 == _1700;
    assign _6576 = _5293 & _6575;
    assign _6584 = _6576 ? _11940 : _6582;
    assign _6586 = _805 ? _4718 : _6584;
    assign _368 = _6586;
    always @(posedge _791) begin
        if (_789)
            _4396 <= _4718;
        else
            _4396 <= _368;
    end
    assign _6593 = _5304 == _1709;
    assign _6590 = ~ _3920;
    assign _6591 = _3135 & _6590;
    assign _6594 = _6591 & _6593;
    assign _6595 = _6594 ? _4693 : _4393;
    assign _6588 = _5296 == _1709;
    assign _6589 = _5293 & _6588;
    assign _6597 = _6589 ? _11940 : _6595;
    assign _6599 = _805 ? _4718 : _6597;
    assign _369 = _6599;
    always @(posedge _791) begin
        if (_789)
            _4393 <= _4718;
        else
            _4393 <= _369;
    end
    assign _6606 = _5304 == _1718;
    assign _6603 = ~ _3920;
    assign _6604 = _3135 & _6603;
    assign _6607 = _6604 & _6606;
    assign _6608 = _6607 ? _4693 : _4390;
    assign _6601 = _5296 == _1718;
    assign _6602 = _5293 & _6601;
    assign _6610 = _6602 ? _11940 : _6608;
    assign _6612 = _805 ? _4718 : _6610;
    assign _370 = _6612;
    always @(posedge _791) begin
        if (_789)
            _4390 <= _4718;
        else
            _4390 <= _370;
    end
    assign _6619 = _5304 == _1727;
    assign _6616 = ~ _3920;
    assign _6617 = _3135 & _6616;
    assign _6620 = _6617 & _6619;
    assign _6621 = _6620 ? _4693 : _4387;
    assign _6614 = _5296 == _1727;
    assign _6615 = _5293 & _6614;
    assign _6623 = _6615 ? _11940 : _6621;
    assign _6625 = _805 ? _4718 : _6623;
    assign _371 = _6625;
    always @(posedge _791) begin
        if (_789)
            _4387 <= _4718;
        else
            _4387 <= _371;
    end
    assign _6632 = _5304 == _1736;
    assign _6629 = ~ _3920;
    assign _6630 = _3135 & _6629;
    assign _6633 = _6630 & _6632;
    assign _6634 = _6633 ? _4693 : _4384;
    assign _6627 = _5296 == _1736;
    assign _6628 = _5293 & _6627;
    assign _6636 = _6628 ? _11940 : _6634;
    assign _6638 = _805 ? _4718 : _6636;
    assign _372 = _6638;
    always @(posedge _791) begin
        if (_789)
            _4384 <= _4718;
        else
            _4384 <= _372;
    end
    assign _6645 = _5304 == _1745;
    assign _6642 = ~ _3920;
    assign _6643 = _3135 & _6642;
    assign _6646 = _6643 & _6645;
    assign _6647 = _6646 ? _4693 : _4381;
    assign _6640 = _5296 == _1745;
    assign _6641 = _5293 & _6640;
    assign _6649 = _6641 ? _11940 : _6647;
    assign _6651 = _805 ? _4718 : _6649;
    assign _373 = _6651;
    always @(posedge _791) begin
        if (_789)
            _4381 <= _4718;
        else
            _4381 <= _373;
    end
    assign _6658 = _5304 == _1754;
    assign _6655 = ~ _3920;
    assign _6656 = _3135 & _6655;
    assign _6659 = _6656 & _6658;
    assign _6660 = _6659 ? _4693 : _4378;
    assign _6653 = _5296 == _1754;
    assign _6654 = _5293 & _6653;
    assign _6662 = _6654 ? _11940 : _6660;
    assign _6664 = _805 ? _4718 : _6662;
    assign _374 = _6664;
    always @(posedge _791) begin
        if (_789)
            _4378 <= _4718;
        else
            _4378 <= _374;
    end
    assign _6671 = _5304 == _1763;
    assign _6668 = ~ _3920;
    assign _6669 = _3135 & _6668;
    assign _6672 = _6669 & _6671;
    assign _6673 = _6672 ? _4693 : _4375;
    assign _6666 = _5296 == _1763;
    assign _6667 = _5293 & _6666;
    assign _6675 = _6667 ? _11940 : _6673;
    assign _6677 = _805 ? _4718 : _6675;
    assign _375 = _6677;
    always @(posedge _791) begin
        if (_789)
            _4375 <= _4718;
        else
            _4375 <= _375;
    end
    assign _6684 = _5304 == _1772;
    assign _6681 = ~ _3920;
    assign _6682 = _3135 & _6681;
    assign _6685 = _6682 & _6684;
    assign _6686 = _6685 ? _4693 : _4372;
    assign _6679 = _5296 == _1772;
    assign _6680 = _5293 & _6679;
    assign _6688 = _6680 ? _11940 : _6686;
    assign _6690 = _805 ? _4718 : _6688;
    assign _376 = _6690;
    always @(posedge _791) begin
        if (_789)
            _4372 <= _4718;
        else
            _4372 <= _376;
    end
    assign _6697 = _5304 == _1781;
    assign _6694 = ~ _3920;
    assign _6695 = _3135 & _6694;
    assign _6698 = _6695 & _6697;
    assign _6699 = _6698 ? _4693 : _4369;
    assign _6692 = _5296 == _1781;
    assign _6693 = _5293 & _6692;
    assign _6701 = _6693 ? _11940 : _6699;
    assign _6703 = _805 ? _4718 : _6701;
    assign _377 = _6703;
    always @(posedge _791) begin
        if (_789)
            _4369 <= _4718;
        else
            _4369 <= _377;
    end
    assign _6710 = _5304 == _1790;
    assign _6707 = ~ _3920;
    assign _6708 = _3135 & _6707;
    assign _6711 = _6708 & _6710;
    assign _6712 = _6711 ? _4693 : _4366;
    assign _6705 = _5296 == _1790;
    assign _6706 = _5293 & _6705;
    assign _6714 = _6706 ? _11940 : _6712;
    assign _6716 = _805 ? _4718 : _6714;
    assign _378 = _6716;
    always @(posedge _791) begin
        if (_789)
            _4366 <= _4718;
        else
            _4366 <= _378;
    end
    assign _6723 = _5304 == _1799;
    assign _6720 = ~ _3920;
    assign _6721 = _3135 & _6720;
    assign _6724 = _6721 & _6723;
    assign _6725 = _6724 ? _4693 : _4363;
    assign _6718 = _5296 == _1799;
    assign _6719 = _5293 & _6718;
    assign _6727 = _6719 ? _11940 : _6725;
    assign _6729 = _805 ? _4718 : _6727;
    assign _379 = _6729;
    always @(posedge _791) begin
        if (_789)
            _4363 <= _4718;
        else
            _4363 <= _379;
    end
    assign _6736 = _5304 == _1808;
    assign _6733 = ~ _3920;
    assign _6734 = _3135 & _6733;
    assign _6737 = _6734 & _6736;
    assign _6738 = _6737 ? _4693 : _4360;
    assign _6731 = _5296 == _1808;
    assign _6732 = _5293 & _6731;
    assign _6740 = _6732 ? _11940 : _6738;
    assign _6742 = _805 ? _4718 : _6740;
    assign _380 = _6742;
    always @(posedge _791) begin
        if (_789)
            _4360 <= _4718;
        else
            _4360 <= _380;
    end
    assign _6749 = _5304 == _1817;
    assign _6746 = ~ _3920;
    assign _6747 = _3135 & _6746;
    assign _6750 = _6747 & _6749;
    assign _6751 = _6750 ? _4693 : _4357;
    assign _6744 = _5296 == _1817;
    assign _6745 = _5293 & _6744;
    assign _6753 = _6745 ? _11940 : _6751;
    assign _6755 = _805 ? _4718 : _6753;
    assign _381 = _6755;
    always @(posedge _791) begin
        if (_789)
            _4357 <= _4718;
        else
            _4357 <= _381;
    end
    assign _6762 = _5304 == _1826;
    assign _6759 = ~ _3920;
    assign _6760 = _3135 & _6759;
    assign _6763 = _6760 & _6762;
    assign _6764 = _6763 ? _4693 : _4354;
    assign _6757 = _5296 == _1826;
    assign _6758 = _5293 & _6757;
    assign _6766 = _6758 ? _11940 : _6764;
    assign _6768 = _805 ? _4718 : _6766;
    assign _382 = _6768;
    always @(posedge _791) begin
        if (_789)
            _4354 <= _4718;
        else
            _4354 <= _382;
    end
    assign _6775 = _5304 == _1835;
    assign _6772 = ~ _3920;
    assign _6773 = _3135 & _6772;
    assign _6776 = _6773 & _6775;
    assign _6777 = _6776 ? _4693 : _4351;
    assign _6770 = _5296 == _1835;
    assign _6771 = _5293 & _6770;
    assign _6779 = _6771 ? _11940 : _6777;
    assign _6781 = _805 ? _4718 : _6779;
    assign _383 = _6781;
    always @(posedge _791) begin
        if (_789)
            _4351 <= _4718;
        else
            _4351 <= _383;
    end
    assign _6788 = _5304 == _1844;
    assign _6785 = ~ _3920;
    assign _6786 = _3135 & _6785;
    assign _6789 = _6786 & _6788;
    assign _6790 = _6789 ? _4693 : _4348;
    assign _6783 = _5296 == _1844;
    assign _6784 = _5293 & _6783;
    assign _6792 = _6784 ? _11940 : _6790;
    assign _6794 = _805 ? _4718 : _6792;
    assign _384 = _6794;
    always @(posedge _791) begin
        if (_789)
            _4348 <= _4718;
        else
            _4348 <= _384;
    end
    assign _6801 = _5304 == _1853;
    assign _6798 = ~ _3920;
    assign _6799 = _3135 & _6798;
    assign _6802 = _6799 & _6801;
    assign _6803 = _6802 ? _4693 : _4345;
    assign _6796 = _5296 == _1853;
    assign _6797 = _5293 & _6796;
    assign _6805 = _6797 ? _11940 : _6803;
    assign _6807 = _805 ? _4718 : _6805;
    assign _385 = _6807;
    always @(posedge _791) begin
        if (_789)
            _4345 <= _4718;
        else
            _4345 <= _385;
    end
    assign _6814 = _5304 == _1862;
    assign _6811 = ~ _3920;
    assign _6812 = _3135 & _6811;
    assign _6815 = _6812 & _6814;
    assign _6816 = _6815 ? _4693 : _4342;
    assign _6809 = _5296 == _1862;
    assign _6810 = _5293 & _6809;
    assign _6818 = _6810 ? _11940 : _6816;
    assign _6820 = _805 ? _4718 : _6818;
    assign _386 = _6820;
    always @(posedge _791) begin
        if (_789)
            _4342 <= _4718;
        else
            _4342 <= _386;
    end
    assign _6827 = _5304 == _1871;
    assign _6824 = ~ _3920;
    assign _6825 = _3135 & _6824;
    assign _6828 = _6825 & _6827;
    assign _6829 = _6828 ? _4693 : _4339;
    assign _6822 = _5296 == _1871;
    assign _6823 = _5293 & _6822;
    assign _6831 = _6823 ? _11940 : _6829;
    assign _6833 = _805 ? _4718 : _6831;
    assign _387 = _6833;
    always @(posedge _791) begin
        if (_789)
            _4339 <= _4718;
        else
            _4339 <= _387;
    end
    assign _6840 = _5304 == _1880;
    assign _6837 = ~ _3920;
    assign _6838 = _3135 & _6837;
    assign _6841 = _6838 & _6840;
    assign _6842 = _6841 ? _4693 : _4336;
    assign _6835 = _5296 == _1880;
    assign _6836 = _5293 & _6835;
    assign _6844 = _6836 ? _11940 : _6842;
    assign _6846 = _805 ? _4718 : _6844;
    assign _388 = _6846;
    always @(posedge _791) begin
        if (_789)
            _4336 <= _4718;
        else
            _4336 <= _388;
    end
    assign _6853 = _5304 == _1889;
    assign _6850 = ~ _3920;
    assign _6851 = _3135 & _6850;
    assign _6854 = _6851 & _6853;
    assign _6855 = _6854 ? _4693 : _4333;
    assign _6848 = _5296 == _1889;
    assign _6849 = _5293 & _6848;
    assign _6857 = _6849 ? _11940 : _6855;
    assign _6859 = _805 ? _4718 : _6857;
    assign _389 = _6859;
    always @(posedge _791) begin
        if (_789)
            _4333 <= _4718;
        else
            _4333 <= _389;
    end
    assign _6866 = _5304 == _1898;
    assign _6863 = ~ _3920;
    assign _6864 = _3135 & _6863;
    assign _6867 = _6864 & _6866;
    assign _6868 = _6867 ? _4693 : _4330;
    assign _6861 = _5296 == _1898;
    assign _6862 = _5293 & _6861;
    assign _6870 = _6862 ? _11940 : _6868;
    assign _6872 = _805 ? _4718 : _6870;
    assign _390 = _6872;
    always @(posedge _791) begin
        if (_789)
            _4330 <= _4718;
        else
            _4330 <= _390;
    end
    assign _6879 = _5304 == _1907;
    assign _6876 = ~ _3920;
    assign _6877 = _3135 & _6876;
    assign _6880 = _6877 & _6879;
    assign _6881 = _6880 ? _4693 : _4327;
    assign _6874 = _5296 == _1907;
    assign _6875 = _5293 & _6874;
    assign _6883 = _6875 ? _11940 : _6881;
    assign _6885 = _805 ? _4718 : _6883;
    assign _391 = _6885;
    always @(posedge _791) begin
        if (_789)
            _4327 <= _4718;
        else
            _4327 <= _391;
    end
    assign _6892 = _5304 == _1916;
    assign _6889 = ~ _3920;
    assign _6890 = _3135 & _6889;
    assign _6893 = _6890 & _6892;
    assign _6894 = _6893 ? _4693 : _4324;
    assign _6887 = _5296 == _1916;
    assign _6888 = _5293 & _6887;
    assign _6896 = _6888 ? _11940 : _6894;
    assign _6898 = _805 ? _4718 : _6896;
    assign _392 = _6898;
    always @(posedge _791) begin
        if (_789)
            _4324 <= _4718;
        else
            _4324 <= _392;
    end
    assign _6905 = _5304 == _1925;
    assign _6902 = ~ _3920;
    assign _6903 = _3135 & _6902;
    assign _6906 = _6903 & _6905;
    assign _6907 = _6906 ? _4693 : _4321;
    assign _6900 = _5296 == _1925;
    assign _6901 = _5293 & _6900;
    assign _6909 = _6901 ? _11940 : _6907;
    assign _6911 = _805 ? _4718 : _6909;
    assign _393 = _6911;
    always @(posedge _791) begin
        if (_789)
            _4321 <= _4718;
        else
            _4321 <= _393;
    end
    assign _6918 = _5304 == _1934;
    assign _6915 = ~ _3920;
    assign _6916 = _3135 & _6915;
    assign _6919 = _6916 & _6918;
    assign _6920 = _6919 ? _4693 : _4318;
    assign _6913 = _5296 == _1934;
    assign _6914 = _5293 & _6913;
    assign _6922 = _6914 ? _11940 : _6920;
    assign _6924 = _805 ? _4718 : _6922;
    assign _394 = _6924;
    always @(posedge _791) begin
        if (_789)
            _4318 <= _4718;
        else
            _4318 <= _394;
    end
    assign _6931 = _5304 == _1943;
    assign _6928 = ~ _3920;
    assign _6929 = _3135 & _6928;
    assign _6932 = _6929 & _6931;
    assign _6933 = _6932 ? _4693 : _4315;
    assign _6926 = _5296 == _1943;
    assign _6927 = _5293 & _6926;
    assign _6935 = _6927 ? _11940 : _6933;
    assign _6937 = _805 ? _4718 : _6935;
    assign _395 = _6937;
    always @(posedge _791) begin
        if (_789)
            _4315 <= _4718;
        else
            _4315 <= _395;
    end
    assign _6944 = _5304 == _1952;
    assign _6941 = ~ _3920;
    assign _6942 = _3135 & _6941;
    assign _6945 = _6942 & _6944;
    assign _6946 = _6945 ? _4693 : _4312;
    assign _6939 = _5296 == _1952;
    assign _6940 = _5293 & _6939;
    assign _6948 = _6940 ? _11940 : _6946;
    assign _6950 = _805 ? _4718 : _6948;
    assign _396 = _6950;
    always @(posedge _791) begin
        if (_789)
            _4312 <= _4718;
        else
            _4312 <= _396;
    end
    assign _6957 = _5304 == _1961;
    assign _6954 = ~ _3920;
    assign _6955 = _3135 & _6954;
    assign _6958 = _6955 & _6957;
    assign _6959 = _6958 ? _4693 : _4309;
    assign _6952 = _5296 == _1961;
    assign _6953 = _5293 & _6952;
    assign _6961 = _6953 ? _11940 : _6959;
    assign _6963 = _805 ? _4718 : _6961;
    assign _397 = _6963;
    always @(posedge _791) begin
        if (_789)
            _4309 <= _4718;
        else
            _4309 <= _397;
    end
    assign _6970 = _5304 == _1970;
    assign _6967 = ~ _3920;
    assign _6968 = _3135 & _6967;
    assign _6971 = _6968 & _6970;
    assign _6972 = _6971 ? _4693 : _4306;
    assign _6965 = _5296 == _1970;
    assign _6966 = _5293 & _6965;
    assign _6974 = _6966 ? _11940 : _6972;
    assign _6976 = _805 ? _4718 : _6974;
    assign _398 = _6976;
    always @(posedge _791) begin
        if (_789)
            _4306 <= _4718;
        else
            _4306 <= _398;
    end
    assign _6983 = _5304 == _1979;
    assign _6980 = ~ _3920;
    assign _6981 = _3135 & _6980;
    assign _6984 = _6981 & _6983;
    assign _6985 = _6984 ? _4693 : _4303;
    assign _6978 = _5296 == _1979;
    assign _6979 = _5293 & _6978;
    assign _6987 = _6979 ? _11940 : _6985;
    assign _6989 = _805 ? _4718 : _6987;
    assign _399 = _6989;
    always @(posedge _791) begin
        if (_789)
            _4303 <= _4718;
        else
            _4303 <= _399;
    end
    assign _6996 = _5304 == _1988;
    assign _6993 = ~ _3920;
    assign _6994 = _3135 & _6993;
    assign _6997 = _6994 & _6996;
    assign _6998 = _6997 ? _4693 : _4300;
    assign _6991 = _5296 == _1988;
    assign _6992 = _5293 & _6991;
    assign _7000 = _6992 ? _11940 : _6998;
    assign _7002 = _805 ? _4718 : _7000;
    assign _400 = _7002;
    always @(posedge _791) begin
        if (_789)
            _4300 <= _4718;
        else
            _4300 <= _400;
    end
    assign _7009 = _5304 == _1997;
    assign _7006 = ~ _3920;
    assign _7007 = _3135 & _7006;
    assign _7010 = _7007 & _7009;
    assign _7011 = _7010 ? _4693 : _4297;
    assign _7004 = _5296 == _1997;
    assign _7005 = _5293 & _7004;
    assign _7013 = _7005 ? _11940 : _7011;
    assign _7015 = _805 ? _4718 : _7013;
    assign _401 = _7015;
    always @(posedge _791) begin
        if (_789)
            _4297 <= _4718;
        else
            _4297 <= _401;
    end
    assign _7022 = _5304 == _2006;
    assign _7019 = ~ _3920;
    assign _7020 = _3135 & _7019;
    assign _7023 = _7020 & _7022;
    assign _7024 = _7023 ? _4693 : _4294;
    assign _7017 = _5296 == _2006;
    assign _7018 = _5293 & _7017;
    assign _7026 = _7018 ? _11940 : _7024;
    assign _7028 = _805 ? _4718 : _7026;
    assign _402 = _7028;
    always @(posedge _791) begin
        if (_789)
            _4294 <= _4718;
        else
            _4294 <= _402;
    end
    assign _7035 = _5304 == _2015;
    assign _7032 = ~ _3920;
    assign _7033 = _3135 & _7032;
    assign _7036 = _7033 & _7035;
    assign _7037 = _7036 ? _4693 : _4291;
    assign _7030 = _5296 == _2015;
    assign _7031 = _5293 & _7030;
    assign _7039 = _7031 ? _11940 : _7037;
    assign _7041 = _805 ? _4718 : _7039;
    assign _403 = _7041;
    always @(posedge _791) begin
        if (_789)
            _4291 <= _4718;
        else
            _4291 <= _403;
    end
    assign _7048 = _5304 == _2024;
    assign _7045 = ~ _3920;
    assign _7046 = _3135 & _7045;
    assign _7049 = _7046 & _7048;
    assign _7050 = _7049 ? _4693 : _4288;
    assign _7043 = _5296 == _2024;
    assign _7044 = _5293 & _7043;
    assign _7052 = _7044 ? _11940 : _7050;
    assign _7054 = _805 ? _4718 : _7052;
    assign _404 = _7054;
    always @(posedge _791) begin
        if (_789)
            _4288 <= _4718;
        else
            _4288 <= _404;
    end
    assign _7061 = _5304 == _2033;
    assign _7058 = ~ _3920;
    assign _7059 = _3135 & _7058;
    assign _7062 = _7059 & _7061;
    assign _7063 = _7062 ? _4693 : _4285;
    assign _7056 = _5296 == _2033;
    assign _7057 = _5293 & _7056;
    assign _7065 = _7057 ? _11940 : _7063;
    assign _7067 = _805 ? _4718 : _7065;
    assign _405 = _7067;
    always @(posedge _791) begin
        if (_789)
            _4285 <= _4718;
        else
            _4285 <= _405;
    end
    assign _7074 = _5304 == _2042;
    assign _7071 = ~ _3920;
    assign _7072 = _3135 & _7071;
    assign _7075 = _7072 & _7074;
    assign _7076 = _7075 ? _4693 : _4282;
    assign _7069 = _5296 == _2042;
    assign _7070 = _5293 & _7069;
    assign _7078 = _7070 ? _11940 : _7076;
    assign _7080 = _805 ? _4718 : _7078;
    assign _406 = _7080;
    always @(posedge _791) begin
        if (_789)
            _4282 <= _4718;
        else
            _4282 <= _406;
    end
    assign _7087 = _5304 == _2051;
    assign _7084 = ~ _3920;
    assign _7085 = _3135 & _7084;
    assign _7088 = _7085 & _7087;
    assign _7089 = _7088 ? _4693 : _4279;
    assign _7082 = _5296 == _2051;
    assign _7083 = _5293 & _7082;
    assign _7091 = _7083 ? _11940 : _7089;
    assign _7093 = _805 ? _4718 : _7091;
    assign _407 = _7093;
    always @(posedge _791) begin
        if (_789)
            _4279 <= _4718;
        else
            _4279 <= _407;
    end
    assign _7100 = _5304 == _2060;
    assign _7097 = ~ _3920;
    assign _7098 = _3135 & _7097;
    assign _7101 = _7098 & _7100;
    assign _7102 = _7101 ? _4693 : _4276;
    assign _7095 = _5296 == _2060;
    assign _7096 = _5293 & _7095;
    assign _7104 = _7096 ? _11940 : _7102;
    assign _7106 = _805 ? _4718 : _7104;
    assign _408 = _7106;
    always @(posedge _791) begin
        if (_789)
            _4276 <= _4718;
        else
            _4276 <= _408;
    end
    assign _7113 = _5304 == _2069;
    assign _7110 = ~ _3920;
    assign _7111 = _3135 & _7110;
    assign _7114 = _7111 & _7113;
    assign _7115 = _7114 ? _4693 : _4273;
    assign _7108 = _5296 == _2069;
    assign _7109 = _5293 & _7108;
    assign _7117 = _7109 ? _11940 : _7115;
    assign _7119 = _805 ? _4718 : _7117;
    assign _409 = _7119;
    always @(posedge _791) begin
        if (_789)
            _4273 <= _4718;
        else
            _4273 <= _409;
    end
    assign _7126 = _5304 == _2078;
    assign _7123 = ~ _3920;
    assign _7124 = _3135 & _7123;
    assign _7127 = _7124 & _7126;
    assign _7128 = _7127 ? _4693 : _4270;
    assign _7121 = _5296 == _2078;
    assign _7122 = _5293 & _7121;
    assign _7130 = _7122 ? _11940 : _7128;
    assign _7132 = _805 ? _4718 : _7130;
    assign _410 = _7132;
    always @(posedge _791) begin
        if (_789)
            _4270 <= _4718;
        else
            _4270 <= _410;
    end
    assign _7139 = _5304 == _2087;
    assign _7136 = ~ _3920;
    assign _7137 = _3135 & _7136;
    assign _7140 = _7137 & _7139;
    assign _7141 = _7140 ? _4693 : _4267;
    assign _7134 = _5296 == _2087;
    assign _7135 = _5293 & _7134;
    assign _7143 = _7135 ? _11940 : _7141;
    assign _7145 = _805 ? _4718 : _7143;
    assign _411 = _7145;
    always @(posedge _791) begin
        if (_789)
            _4267 <= _4718;
        else
            _4267 <= _411;
    end
    assign _7152 = _5304 == _2096;
    assign _7149 = ~ _3920;
    assign _7150 = _3135 & _7149;
    assign _7153 = _7150 & _7152;
    assign _7154 = _7153 ? _4693 : _4264;
    assign _7147 = _5296 == _2096;
    assign _7148 = _5293 & _7147;
    assign _7156 = _7148 ? _11940 : _7154;
    assign _7158 = _805 ? _4718 : _7156;
    assign _412 = _7158;
    always @(posedge _791) begin
        if (_789)
            _4264 <= _4718;
        else
            _4264 <= _412;
    end
    assign _7165 = _5304 == _2105;
    assign _7162 = ~ _3920;
    assign _7163 = _3135 & _7162;
    assign _7166 = _7163 & _7165;
    assign _7167 = _7166 ? _4693 : _4261;
    assign _7160 = _5296 == _2105;
    assign _7161 = _5293 & _7160;
    assign _7169 = _7161 ? _11940 : _7167;
    assign _7171 = _805 ? _4718 : _7169;
    assign _413 = _7171;
    always @(posedge _791) begin
        if (_789)
            _4261 <= _4718;
        else
            _4261 <= _413;
    end
    assign _7178 = _5304 == _2114;
    assign _7175 = ~ _3920;
    assign _7176 = _3135 & _7175;
    assign _7179 = _7176 & _7178;
    assign _7180 = _7179 ? _4693 : _4258;
    assign _7173 = _5296 == _2114;
    assign _7174 = _5293 & _7173;
    assign _7182 = _7174 ? _11940 : _7180;
    assign _7184 = _805 ? _4718 : _7182;
    assign _414 = _7184;
    always @(posedge _791) begin
        if (_789)
            _4258 <= _4718;
        else
            _4258 <= _414;
    end
    assign _7191 = _5304 == _2123;
    assign _7188 = ~ _3920;
    assign _7189 = _3135 & _7188;
    assign _7192 = _7189 & _7191;
    assign _7193 = _7192 ? _4693 : _4255;
    assign _7186 = _5296 == _2123;
    assign _7187 = _5293 & _7186;
    assign _7195 = _7187 ? _11940 : _7193;
    assign _7197 = _805 ? _4718 : _7195;
    assign _415 = _7197;
    always @(posedge _791) begin
        if (_789)
            _4255 <= _4718;
        else
            _4255 <= _415;
    end
    assign _7204 = _5304 == _2132;
    assign _7201 = ~ _3920;
    assign _7202 = _3135 & _7201;
    assign _7205 = _7202 & _7204;
    assign _7206 = _7205 ? _4693 : _4252;
    assign _7199 = _5296 == _2132;
    assign _7200 = _5293 & _7199;
    assign _7208 = _7200 ? _11940 : _7206;
    assign _7210 = _805 ? _4718 : _7208;
    assign _416 = _7210;
    always @(posedge _791) begin
        if (_789)
            _4252 <= _4718;
        else
            _4252 <= _416;
    end
    assign _7217 = _5304 == _2141;
    assign _7214 = ~ _3920;
    assign _7215 = _3135 & _7214;
    assign _7218 = _7215 & _7217;
    assign _7219 = _7218 ? _4693 : _4249;
    assign _7212 = _5296 == _2141;
    assign _7213 = _5293 & _7212;
    assign _7221 = _7213 ? _11940 : _7219;
    assign _7223 = _805 ? _4718 : _7221;
    assign _417 = _7223;
    always @(posedge _791) begin
        if (_789)
            _4249 <= _4718;
        else
            _4249 <= _417;
    end
    assign _7230 = _5304 == _2150;
    assign _7227 = ~ _3920;
    assign _7228 = _3135 & _7227;
    assign _7231 = _7228 & _7230;
    assign _7232 = _7231 ? _4693 : _4246;
    assign _7225 = _5296 == _2150;
    assign _7226 = _5293 & _7225;
    assign _7234 = _7226 ? _11940 : _7232;
    assign _7236 = _805 ? _4718 : _7234;
    assign _418 = _7236;
    always @(posedge _791) begin
        if (_789)
            _4246 <= _4718;
        else
            _4246 <= _418;
    end
    assign _7243 = _5304 == _2159;
    assign _7240 = ~ _3920;
    assign _7241 = _3135 & _7240;
    assign _7244 = _7241 & _7243;
    assign _7245 = _7244 ? _4693 : _4243;
    assign _7238 = _5296 == _2159;
    assign _7239 = _5293 & _7238;
    assign _7247 = _7239 ? _11940 : _7245;
    assign _7249 = _805 ? _4718 : _7247;
    assign _419 = _7249;
    always @(posedge _791) begin
        if (_789)
            _4243 <= _4718;
        else
            _4243 <= _419;
    end
    assign _7256 = _5304 == _2168;
    assign _7253 = ~ _3920;
    assign _7254 = _3135 & _7253;
    assign _7257 = _7254 & _7256;
    assign _7258 = _7257 ? _4693 : _4240;
    assign _7251 = _5296 == _2168;
    assign _7252 = _5293 & _7251;
    assign _7260 = _7252 ? _11940 : _7258;
    assign _7262 = _805 ? _4718 : _7260;
    assign _420 = _7262;
    always @(posedge _791) begin
        if (_789)
            _4240 <= _4718;
        else
            _4240 <= _420;
    end
    assign _7269 = _5304 == _2177;
    assign _7266 = ~ _3920;
    assign _7267 = _3135 & _7266;
    assign _7270 = _7267 & _7269;
    assign _7271 = _7270 ? _4693 : _4237;
    assign _7264 = _5296 == _2177;
    assign _7265 = _5293 & _7264;
    assign _7273 = _7265 ? _11940 : _7271;
    assign _7275 = _805 ? _4718 : _7273;
    assign _421 = _7275;
    always @(posedge _791) begin
        if (_789)
            _4237 <= _4718;
        else
            _4237 <= _421;
    end
    assign _7282 = _5304 == _2186;
    assign _7279 = ~ _3920;
    assign _7280 = _3135 & _7279;
    assign _7283 = _7280 & _7282;
    assign _7284 = _7283 ? _4693 : _4234;
    assign _7277 = _5296 == _2186;
    assign _7278 = _5293 & _7277;
    assign _7286 = _7278 ? _11940 : _7284;
    assign _7288 = _805 ? _4718 : _7286;
    assign _422 = _7288;
    always @(posedge _791) begin
        if (_789)
            _4234 <= _4718;
        else
            _4234 <= _422;
    end
    assign _7295 = _5304 == _2195;
    assign _7292 = ~ _3920;
    assign _7293 = _3135 & _7292;
    assign _7296 = _7293 & _7295;
    assign _7297 = _7296 ? _4693 : _4231;
    assign _7290 = _5296 == _2195;
    assign _7291 = _5293 & _7290;
    assign _7299 = _7291 ? _11940 : _7297;
    assign _7301 = _805 ? _4718 : _7299;
    assign _423 = _7301;
    always @(posedge _791) begin
        if (_789)
            _4231 <= _4718;
        else
            _4231 <= _423;
    end
    assign _7308 = _5304 == _2204;
    assign _7305 = ~ _3920;
    assign _7306 = _3135 & _7305;
    assign _7309 = _7306 & _7308;
    assign _7310 = _7309 ? _4693 : _4228;
    assign _7303 = _5296 == _2204;
    assign _7304 = _5293 & _7303;
    assign _7312 = _7304 ? _11940 : _7310;
    assign _7314 = _805 ? _4718 : _7312;
    assign _424 = _7314;
    always @(posedge _791) begin
        if (_789)
            _4228 <= _4718;
        else
            _4228 <= _424;
    end
    assign _7321 = _5304 == _2213;
    assign _7318 = ~ _3920;
    assign _7319 = _3135 & _7318;
    assign _7322 = _7319 & _7321;
    assign _7323 = _7322 ? _4693 : _4225;
    assign _7316 = _5296 == _2213;
    assign _7317 = _5293 & _7316;
    assign _7325 = _7317 ? _11940 : _7323;
    assign _7327 = _805 ? _4718 : _7325;
    assign _425 = _7327;
    always @(posedge _791) begin
        if (_789)
            _4225 <= _4718;
        else
            _4225 <= _425;
    end
    assign _7334 = _5304 == _2222;
    assign _7331 = ~ _3920;
    assign _7332 = _3135 & _7331;
    assign _7335 = _7332 & _7334;
    assign _7336 = _7335 ? _4693 : _4222;
    assign _7329 = _5296 == _2222;
    assign _7330 = _5293 & _7329;
    assign _7338 = _7330 ? _11940 : _7336;
    assign _7340 = _805 ? _4718 : _7338;
    assign _426 = _7340;
    always @(posedge _791) begin
        if (_789)
            _4222 <= _4718;
        else
            _4222 <= _426;
    end
    assign _7347 = _5304 == _2231;
    assign _7344 = ~ _3920;
    assign _7345 = _3135 & _7344;
    assign _7348 = _7345 & _7347;
    assign _7349 = _7348 ? _4693 : _4219;
    assign _7342 = _5296 == _2231;
    assign _7343 = _5293 & _7342;
    assign _7351 = _7343 ? _11940 : _7349;
    assign _7353 = _805 ? _4718 : _7351;
    assign _427 = _7353;
    always @(posedge _791) begin
        if (_789)
            _4219 <= _4718;
        else
            _4219 <= _427;
    end
    assign _7360 = _5304 == _2240;
    assign _7357 = ~ _3920;
    assign _7358 = _3135 & _7357;
    assign _7361 = _7358 & _7360;
    assign _7362 = _7361 ? _4693 : _4216;
    assign _7355 = _5296 == _2240;
    assign _7356 = _5293 & _7355;
    assign _7364 = _7356 ? _11940 : _7362;
    assign _7366 = _805 ? _4718 : _7364;
    assign _428 = _7366;
    always @(posedge _791) begin
        if (_789)
            _4216 <= _4718;
        else
            _4216 <= _428;
    end
    assign _7373 = _5304 == _2249;
    assign _7370 = ~ _3920;
    assign _7371 = _3135 & _7370;
    assign _7374 = _7371 & _7373;
    assign _7375 = _7374 ? _4693 : _4213;
    assign _7368 = _5296 == _2249;
    assign _7369 = _5293 & _7368;
    assign _7377 = _7369 ? _11940 : _7375;
    assign _7379 = _805 ? _4718 : _7377;
    assign _429 = _7379;
    always @(posedge _791) begin
        if (_789)
            _4213 <= _4718;
        else
            _4213 <= _429;
    end
    assign _7386 = _5304 == _2258;
    assign _7383 = ~ _3920;
    assign _7384 = _3135 & _7383;
    assign _7387 = _7384 & _7386;
    assign _7388 = _7387 ? _4693 : _4210;
    assign _7381 = _5296 == _2258;
    assign _7382 = _5293 & _7381;
    assign _7390 = _7382 ? _11940 : _7388;
    assign _7392 = _805 ? _4718 : _7390;
    assign _430 = _7392;
    always @(posedge _791) begin
        if (_789)
            _4210 <= _4718;
        else
            _4210 <= _430;
    end
    assign _7399 = _5304 == _2267;
    assign _7396 = ~ _3920;
    assign _7397 = _3135 & _7396;
    assign _7400 = _7397 & _7399;
    assign _7401 = _7400 ? _4693 : _4207;
    assign _7394 = _5296 == _2267;
    assign _7395 = _5293 & _7394;
    assign _7403 = _7395 ? _11940 : _7401;
    assign _7405 = _805 ? _4718 : _7403;
    assign _431 = _7405;
    always @(posedge _791) begin
        if (_789)
            _4207 <= _4718;
        else
            _4207 <= _431;
    end
    assign _7412 = _5304 == _2276;
    assign _7409 = ~ _3920;
    assign _7410 = _3135 & _7409;
    assign _7413 = _7410 & _7412;
    assign _7414 = _7413 ? _4693 : _4204;
    assign _7407 = _5296 == _2276;
    assign _7408 = _5293 & _7407;
    assign _7416 = _7408 ? _11940 : _7414;
    assign _7418 = _805 ? _4718 : _7416;
    assign _432 = _7418;
    always @(posedge _791) begin
        if (_789)
            _4204 <= _4718;
        else
            _4204 <= _432;
    end
    assign _7425 = _5304 == _2285;
    assign _7422 = ~ _3920;
    assign _7423 = _3135 & _7422;
    assign _7426 = _7423 & _7425;
    assign _7427 = _7426 ? _4693 : _4201;
    assign _7420 = _5296 == _2285;
    assign _7421 = _5293 & _7420;
    assign _7429 = _7421 ? _11940 : _7427;
    assign _7431 = _805 ? _4718 : _7429;
    assign _433 = _7431;
    always @(posedge _791) begin
        if (_789)
            _4201 <= _4718;
        else
            _4201 <= _433;
    end
    assign _7438 = _5304 == _2294;
    assign _7435 = ~ _3920;
    assign _7436 = _3135 & _7435;
    assign _7439 = _7436 & _7438;
    assign _7440 = _7439 ? _4693 : _4198;
    assign _7433 = _5296 == _2294;
    assign _7434 = _5293 & _7433;
    assign _7442 = _7434 ? _11940 : _7440;
    assign _7444 = _805 ? _4718 : _7442;
    assign _434 = _7444;
    always @(posedge _791) begin
        if (_789)
            _4198 <= _4718;
        else
            _4198 <= _434;
    end
    assign _7451 = _5304 == _2303;
    assign _7448 = ~ _3920;
    assign _7449 = _3135 & _7448;
    assign _7452 = _7449 & _7451;
    assign _7453 = _7452 ? _4693 : _4195;
    assign _7446 = _5296 == _2303;
    assign _7447 = _5293 & _7446;
    assign _7455 = _7447 ? _11940 : _7453;
    assign _7457 = _805 ? _4718 : _7455;
    assign _435 = _7457;
    always @(posedge _791) begin
        if (_789)
            _4195 <= _4718;
        else
            _4195 <= _435;
    end
    assign _7464 = _5304 == _2312;
    assign _7461 = ~ _3920;
    assign _7462 = _3135 & _7461;
    assign _7465 = _7462 & _7464;
    assign _7466 = _7465 ? _4693 : _4192;
    assign _7459 = _5296 == _2312;
    assign _7460 = _5293 & _7459;
    assign _7468 = _7460 ? _11940 : _7466;
    assign _7470 = _805 ? _4718 : _7468;
    assign _436 = _7470;
    always @(posedge _791) begin
        if (_789)
            _4192 <= _4718;
        else
            _4192 <= _436;
    end
    assign _7477 = _5304 == _2321;
    assign _7474 = ~ _3920;
    assign _7475 = _3135 & _7474;
    assign _7478 = _7475 & _7477;
    assign _7479 = _7478 ? _4693 : _4189;
    assign _7472 = _5296 == _2321;
    assign _7473 = _5293 & _7472;
    assign _7481 = _7473 ? _11940 : _7479;
    assign _7483 = _805 ? _4718 : _7481;
    assign _437 = _7483;
    always @(posedge _791) begin
        if (_789)
            _4189 <= _4718;
        else
            _4189 <= _437;
    end
    assign _7490 = _5304 == _2330;
    assign _7487 = ~ _3920;
    assign _7488 = _3135 & _7487;
    assign _7491 = _7488 & _7490;
    assign _7492 = _7491 ? _4693 : _4186;
    assign _7485 = _5296 == _2330;
    assign _7486 = _5293 & _7485;
    assign _7494 = _7486 ? _11940 : _7492;
    assign _7496 = _805 ? _4718 : _7494;
    assign _438 = _7496;
    always @(posedge _791) begin
        if (_789)
            _4186 <= _4718;
        else
            _4186 <= _438;
    end
    assign _7503 = _5304 == _2339;
    assign _7500 = ~ _3920;
    assign _7501 = _3135 & _7500;
    assign _7504 = _7501 & _7503;
    assign _7505 = _7504 ? _4693 : _4183;
    assign _7498 = _5296 == _2339;
    assign _7499 = _5293 & _7498;
    assign _7507 = _7499 ? _11940 : _7505;
    assign _7509 = _805 ? _4718 : _7507;
    assign _439 = _7509;
    always @(posedge _791) begin
        if (_789)
            _4183 <= _4718;
        else
            _4183 <= _439;
    end
    assign _7516 = _5304 == _2348;
    assign _7513 = ~ _3920;
    assign _7514 = _3135 & _7513;
    assign _7517 = _7514 & _7516;
    assign _7518 = _7517 ? _4693 : _4180;
    assign _7511 = _5296 == _2348;
    assign _7512 = _5293 & _7511;
    assign _7520 = _7512 ? _11940 : _7518;
    assign _7522 = _805 ? _4718 : _7520;
    assign _440 = _7522;
    always @(posedge _791) begin
        if (_789)
            _4180 <= _4718;
        else
            _4180 <= _440;
    end
    assign _7529 = _5304 == _2357;
    assign _7526 = ~ _3920;
    assign _7527 = _3135 & _7526;
    assign _7530 = _7527 & _7529;
    assign _7531 = _7530 ? _4693 : _4177;
    assign _7524 = _5296 == _2357;
    assign _7525 = _5293 & _7524;
    assign _7533 = _7525 ? _11940 : _7531;
    assign _7535 = _805 ? _4718 : _7533;
    assign _441 = _7535;
    always @(posedge _791) begin
        if (_789)
            _4177 <= _4718;
        else
            _4177 <= _441;
    end
    assign _7542 = _5304 == _2366;
    assign _7539 = ~ _3920;
    assign _7540 = _3135 & _7539;
    assign _7543 = _7540 & _7542;
    assign _7544 = _7543 ? _4693 : _4174;
    assign _7537 = _5296 == _2366;
    assign _7538 = _5293 & _7537;
    assign _7546 = _7538 ? _11940 : _7544;
    assign _7548 = _805 ? _4718 : _7546;
    assign _442 = _7548;
    always @(posedge _791) begin
        if (_789)
            _4174 <= _4718;
        else
            _4174 <= _442;
    end
    assign _7555 = _5304 == _2375;
    assign _7552 = ~ _3920;
    assign _7553 = _3135 & _7552;
    assign _7556 = _7553 & _7555;
    assign _7557 = _7556 ? _4693 : _4171;
    assign _7550 = _5296 == _2375;
    assign _7551 = _5293 & _7550;
    assign _7559 = _7551 ? _11940 : _7557;
    assign _7561 = _805 ? _4718 : _7559;
    assign _443 = _7561;
    always @(posedge _791) begin
        if (_789)
            _4171 <= _4718;
        else
            _4171 <= _443;
    end
    assign _7568 = _5304 == _2384;
    assign _7565 = ~ _3920;
    assign _7566 = _3135 & _7565;
    assign _7569 = _7566 & _7568;
    assign _7570 = _7569 ? _4693 : _4168;
    assign _7563 = _5296 == _2384;
    assign _7564 = _5293 & _7563;
    assign _7572 = _7564 ? _11940 : _7570;
    assign _7574 = _805 ? _4718 : _7572;
    assign _444 = _7574;
    always @(posedge _791) begin
        if (_789)
            _4168 <= _4718;
        else
            _4168 <= _444;
    end
    assign _7581 = _5304 == _2393;
    assign _7578 = ~ _3920;
    assign _7579 = _3135 & _7578;
    assign _7582 = _7579 & _7581;
    assign _7583 = _7582 ? _4693 : _4165;
    assign _7576 = _5296 == _2393;
    assign _7577 = _5293 & _7576;
    assign _7585 = _7577 ? _11940 : _7583;
    assign _7587 = _805 ? _4718 : _7585;
    assign _445 = _7587;
    always @(posedge _791) begin
        if (_789)
            _4165 <= _4718;
        else
            _4165 <= _445;
    end
    assign _7594 = _5304 == _2402;
    assign _7591 = ~ _3920;
    assign _7592 = _3135 & _7591;
    assign _7595 = _7592 & _7594;
    assign _7596 = _7595 ? _4693 : _4162;
    assign _7589 = _5296 == _2402;
    assign _7590 = _5293 & _7589;
    assign _7598 = _7590 ? _11940 : _7596;
    assign _7600 = _805 ? _4718 : _7598;
    assign _446 = _7600;
    always @(posedge _791) begin
        if (_789)
            _4162 <= _4718;
        else
            _4162 <= _446;
    end
    assign _7607 = _5304 == _2411;
    assign _7604 = ~ _3920;
    assign _7605 = _3135 & _7604;
    assign _7608 = _7605 & _7607;
    assign _7609 = _7608 ? _4693 : _4159;
    assign _7602 = _5296 == _2411;
    assign _7603 = _5293 & _7602;
    assign _7611 = _7603 ? _11940 : _7609;
    assign _7613 = _805 ? _4718 : _7611;
    assign _447 = _7613;
    always @(posedge _791) begin
        if (_789)
            _4159 <= _4718;
        else
            _4159 <= _447;
    end
    assign _7620 = _5304 == _2420;
    assign _7617 = ~ _3920;
    assign _7618 = _3135 & _7617;
    assign _7621 = _7618 & _7620;
    assign _7622 = _7621 ? _4693 : _4156;
    assign _7615 = _5296 == _2420;
    assign _7616 = _5293 & _7615;
    assign _7624 = _7616 ? _11940 : _7622;
    assign _7626 = _805 ? _4718 : _7624;
    assign _448 = _7626;
    always @(posedge _791) begin
        if (_789)
            _4156 <= _4718;
        else
            _4156 <= _448;
    end
    assign _7633 = _5304 == _2429;
    assign _7630 = ~ _3920;
    assign _7631 = _3135 & _7630;
    assign _7634 = _7631 & _7633;
    assign _7635 = _7634 ? _4693 : _4153;
    assign _7628 = _5296 == _2429;
    assign _7629 = _5293 & _7628;
    assign _7637 = _7629 ? _11940 : _7635;
    assign _7639 = _805 ? _4718 : _7637;
    assign _449 = _7639;
    always @(posedge _791) begin
        if (_789)
            _4153 <= _4718;
        else
            _4153 <= _449;
    end
    assign _7646 = _5304 == _2438;
    assign _7643 = ~ _3920;
    assign _7644 = _3135 & _7643;
    assign _7647 = _7644 & _7646;
    assign _7648 = _7647 ? _4693 : _4150;
    assign _7641 = _5296 == _2438;
    assign _7642 = _5293 & _7641;
    assign _7650 = _7642 ? _11940 : _7648;
    assign _7652 = _805 ? _4718 : _7650;
    assign _450 = _7652;
    always @(posedge _791) begin
        if (_789)
            _4150 <= _4718;
        else
            _4150 <= _450;
    end
    assign _7659 = _5304 == _2447;
    assign _7656 = ~ _3920;
    assign _7657 = _3135 & _7656;
    assign _7660 = _7657 & _7659;
    assign _7661 = _7660 ? _4693 : _4147;
    assign _7654 = _5296 == _2447;
    assign _7655 = _5293 & _7654;
    assign _7663 = _7655 ? _11940 : _7661;
    assign _7665 = _805 ? _4718 : _7663;
    assign _451 = _7665;
    always @(posedge _791) begin
        if (_789)
            _4147 <= _4718;
        else
            _4147 <= _451;
    end
    assign _7672 = _5304 == _2456;
    assign _7669 = ~ _3920;
    assign _7670 = _3135 & _7669;
    assign _7673 = _7670 & _7672;
    assign _7674 = _7673 ? _4693 : _4144;
    assign _7667 = _5296 == _2456;
    assign _7668 = _5293 & _7667;
    assign _7676 = _7668 ? _11940 : _7674;
    assign _7678 = _805 ? _4718 : _7676;
    assign _452 = _7678;
    always @(posedge _791) begin
        if (_789)
            _4144 <= _4718;
        else
            _4144 <= _452;
    end
    assign _7685 = _5304 == _2465;
    assign _7682 = ~ _3920;
    assign _7683 = _3135 & _7682;
    assign _7686 = _7683 & _7685;
    assign _7687 = _7686 ? _4693 : _4141;
    assign _7680 = _5296 == _2465;
    assign _7681 = _5293 & _7680;
    assign _7689 = _7681 ? _11940 : _7687;
    assign _7691 = _805 ? _4718 : _7689;
    assign _453 = _7691;
    always @(posedge _791) begin
        if (_789)
            _4141 <= _4718;
        else
            _4141 <= _453;
    end
    assign _7698 = _5304 == _2474;
    assign _7695 = ~ _3920;
    assign _7696 = _3135 & _7695;
    assign _7699 = _7696 & _7698;
    assign _7700 = _7699 ? _4693 : _4138;
    assign _7693 = _5296 == _2474;
    assign _7694 = _5293 & _7693;
    assign _7702 = _7694 ? _11940 : _7700;
    assign _7704 = _805 ? _4718 : _7702;
    assign _454 = _7704;
    always @(posedge _791) begin
        if (_789)
            _4138 <= _4718;
        else
            _4138 <= _454;
    end
    assign _7711 = _5304 == _2483;
    assign _7708 = ~ _3920;
    assign _7709 = _3135 & _7708;
    assign _7712 = _7709 & _7711;
    assign _7713 = _7712 ? _4693 : _4135;
    assign _7706 = _5296 == _2483;
    assign _7707 = _5293 & _7706;
    assign _7715 = _7707 ? _11940 : _7713;
    assign _7717 = _805 ? _4718 : _7715;
    assign _455 = _7717;
    always @(posedge _791) begin
        if (_789)
            _4135 <= _4718;
        else
            _4135 <= _455;
    end
    assign _7724 = _5304 == _2492;
    assign _7721 = ~ _3920;
    assign _7722 = _3135 & _7721;
    assign _7725 = _7722 & _7724;
    assign _7726 = _7725 ? _4693 : _4132;
    assign _7719 = _5296 == _2492;
    assign _7720 = _5293 & _7719;
    assign _7728 = _7720 ? _11940 : _7726;
    assign _7730 = _805 ? _4718 : _7728;
    assign _456 = _7730;
    always @(posedge _791) begin
        if (_789)
            _4132 <= _4718;
        else
            _4132 <= _456;
    end
    assign _7737 = _5304 == _2501;
    assign _7734 = ~ _3920;
    assign _7735 = _3135 & _7734;
    assign _7738 = _7735 & _7737;
    assign _7739 = _7738 ? _4693 : _4129;
    assign _7732 = _5296 == _2501;
    assign _7733 = _5293 & _7732;
    assign _7741 = _7733 ? _11940 : _7739;
    assign _7743 = _805 ? _4718 : _7741;
    assign _457 = _7743;
    always @(posedge _791) begin
        if (_789)
            _4129 <= _4718;
        else
            _4129 <= _457;
    end
    assign _7750 = _5304 == _2510;
    assign _7747 = ~ _3920;
    assign _7748 = _3135 & _7747;
    assign _7751 = _7748 & _7750;
    assign _7752 = _7751 ? _4693 : _4126;
    assign _7745 = _5296 == _2510;
    assign _7746 = _5293 & _7745;
    assign _7754 = _7746 ? _11940 : _7752;
    assign _7756 = _805 ? _4718 : _7754;
    assign _458 = _7756;
    always @(posedge _791) begin
        if (_789)
            _4126 <= _4718;
        else
            _4126 <= _458;
    end
    assign _7763 = _5304 == _2519;
    assign _7760 = ~ _3920;
    assign _7761 = _3135 & _7760;
    assign _7764 = _7761 & _7763;
    assign _7765 = _7764 ? _4693 : _4123;
    assign _7758 = _5296 == _2519;
    assign _7759 = _5293 & _7758;
    assign _7767 = _7759 ? _11940 : _7765;
    assign _7769 = _805 ? _4718 : _7767;
    assign _459 = _7769;
    always @(posedge _791) begin
        if (_789)
            _4123 <= _4718;
        else
            _4123 <= _459;
    end
    assign _7776 = _5304 == _2528;
    assign _7773 = ~ _3920;
    assign _7774 = _3135 & _7773;
    assign _7777 = _7774 & _7776;
    assign _7778 = _7777 ? _4693 : _4120;
    assign _7771 = _5296 == _2528;
    assign _7772 = _5293 & _7771;
    assign _7780 = _7772 ? _11940 : _7778;
    assign _7782 = _805 ? _4718 : _7780;
    assign _460 = _7782;
    always @(posedge _791) begin
        if (_789)
            _4120 <= _4718;
        else
            _4120 <= _460;
    end
    assign _7789 = _5304 == _2537;
    assign _7786 = ~ _3920;
    assign _7787 = _3135 & _7786;
    assign _7790 = _7787 & _7789;
    assign _7791 = _7790 ? _4693 : _4117;
    assign _7784 = _5296 == _2537;
    assign _7785 = _5293 & _7784;
    assign _7793 = _7785 ? _11940 : _7791;
    assign _7795 = _805 ? _4718 : _7793;
    assign _461 = _7795;
    always @(posedge _791) begin
        if (_789)
            _4117 <= _4718;
        else
            _4117 <= _461;
    end
    assign _7802 = _5304 == _2546;
    assign _7799 = ~ _3920;
    assign _7800 = _3135 & _7799;
    assign _7803 = _7800 & _7802;
    assign _7804 = _7803 ? _4693 : _4114;
    assign _7797 = _5296 == _2546;
    assign _7798 = _5293 & _7797;
    assign _7806 = _7798 ? _11940 : _7804;
    assign _7808 = _805 ? _4718 : _7806;
    assign _462 = _7808;
    always @(posedge _791) begin
        if (_789)
            _4114 <= _4718;
        else
            _4114 <= _462;
    end
    assign _7815 = _5304 == _2555;
    assign _7812 = ~ _3920;
    assign _7813 = _3135 & _7812;
    assign _7816 = _7813 & _7815;
    assign _7817 = _7816 ? _4693 : _4111;
    assign _7810 = _5296 == _2555;
    assign _7811 = _5293 & _7810;
    assign _7819 = _7811 ? _11940 : _7817;
    assign _7821 = _805 ? _4718 : _7819;
    assign _463 = _7821;
    always @(posedge _791) begin
        if (_789)
            _4111 <= _4718;
        else
            _4111 <= _463;
    end
    assign _7828 = _5304 == _2564;
    assign _7825 = ~ _3920;
    assign _7826 = _3135 & _7825;
    assign _7829 = _7826 & _7828;
    assign _7830 = _7829 ? _4693 : _4108;
    assign _7823 = _5296 == _2564;
    assign _7824 = _5293 & _7823;
    assign _7832 = _7824 ? _11940 : _7830;
    assign _7834 = _805 ? _4718 : _7832;
    assign _464 = _7834;
    always @(posedge _791) begin
        if (_789)
            _4108 <= _4718;
        else
            _4108 <= _464;
    end
    assign _7841 = _5304 == _2573;
    assign _7838 = ~ _3920;
    assign _7839 = _3135 & _7838;
    assign _7842 = _7839 & _7841;
    assign _7843 = _7842 ? _4693 : _4105;
    assign _7836 = _5296 == _2573;
    assign _7837 = _5293 & _7836;
    assign _7845 = _7837 ? _11940 : _7843;
    assign _7847 = _805 ? _4718 : _7845;
    assign _465 = _7847;
    always @(posedge _791) begin
        if (_789)
            _4105 <= _4718;
        else
            _4105 <= _465;
    end
    assign _7854 = _5304 == _2582;
    assign _7851 = ~ _3920;
    assign _7852 = _3135 & _7851;
    assign _7855 = _7852 & _7854;
    assign _7856 = _7855 ? _4693 : _4102;
    assign _7849 = _5296 == _2582;
    assign _7850 = _5293 & _7849;
    assign _7858 = _7850 ? _11940 : _7856;
    assign _7860 = _805 ? _4718 : _7858;
    assign _466 = _7860;
    always @(posedge _791) begin
        if (_789)
            _4102 <= _4718;
        else
            _4102 <= _466;
    end
    assign _7867 = _5304 == _2591;
    assign _7864 = ~ _3920;
    assign _7865 = _3135 & _7864;
    assign _7868 = _7865 & _7867;
    assign _7869 = _7868 ? _4693 : _4099;
    assign _7862 = _5296 == _2591;
    assign _7863 = _5293 & _7862;
    assign _7871 = _7863 ? _11940 : _7869;
    assign _7873 = _805 ? _4718 : _7871;
    assign _467 = _7873;
    always @(posedge _791) begin
        if (_789)
            _4099 <= _4718;
        else
            _4099 <= _467;
    end
    assign _7880 = _5304 == _2600;
    assign _7877 = ~ _3920;
    assign _7878 = _3135 & _7877;
    assign _7881 = _7878 & _7880;
    assign _7882 = _7881 ? _4693 : _4096;
    assign _7875 = _5296 == _2600;
    assign _7876 = _5293 & _7875;
    assign _7884 = _7876 ? _11940 : _7882;
    assign _7886 = _805 ? _4718 : _7884;
    assign _468 = _7886;
    always @(posedge _791) begin
        if (_789)
            _4096 <= _4718;
        else
            _4096 <= _468;
    end
    assign _7893 = _5304 == _2609;
    assign _7890 = ~ _3920;
    assign _7891 = _3135 & _7890;
    assign _7894 = _7891 & _7893;
    assign _7895 = _7894 ? _4693 : _4093;
    assign _7888 = _5296 == _2609;
    assign _7889 = _5293 & _7888;
    assign _7897 = _7889 ? _11940 : _7895;
    assign _7899 = _805 ? _4718 : _7897;
    assign _469 = _7899;
    always @(posedge _791) begin
        if (_789)
            _4093 <= _4718;
        else
            _4093 <= _469;
    end
    assign _7906 = _5304 == _2618;
    assign _7903 = ~ _3920;
    assign _7904 = _3135 & _7903;
    assign _7907 = _7904 & _7906;
    assign _7908 = _7907 ? _4693 : _4090;
    assign _7901 = _5296 == _2618;
    assign _7902 = _5293 & _7901;
    assign _7910 = _7902 ? _11940 : _7908;
    assign _7912 = _805 ? _4718 : _7910;
    assign _470 = _7912;
    always @(posedge _791) begin
        if (_789)
            _4090 <= _4718;
        else
            _4090 <= _470;
    end
    assign _7919 = _5304 == _2627;
    assign _7916 = ~ _3920;
    assign _7917 = _3135 & _7916;
    assign _7920 = _7917 & _7919;
    assign _7921 = _7920 ? _4693 : _4087;
    assign _7914 = _5296 == _2627;
    assign _7915 = _5293 & _7914;
    assign _7923 = _7915 ? _11940 : _7921;
    assign _7925 = _805 ? _4718 : _7923;
    assign _471 = _7925;
    always @(posedge _791) begin
        if (_789)
            _4087 <= _4718;
        else
            _4087 <= _471;
    end
    assign _7932 = _5304 == _2636;
    assign _7929 = ~ _3920;
    assign _7930 = _3135 & _7929;
    assign _7933 = _7930 & _7932;
    assign _7934 = _7933 ? _4693 : _4084;
    assign _7927 = _5296 == _2636;
    assign _7928 = _5293 & _7927;
    assign _7936 = _7928 ? _11940 : _7934;
    assign _7938 = _805 ? _4718 : _7936;
    assign _472 = _7938;
    always @(posedge _791) begin
        if (_789)
            _4084 <= _4718;
        else
            _4084 <= _472;
    end
    assign _7945 = _5304 == _2645;
    assign _7942 = ~ _3920;
    assign _7943 = _3135 & _7942;
    assign _7946 = _7943 & _7945;
    assign _7947 = _7946 ? _4693 : _4081;
    assign _7940 = _5296 == _2645;
    assign _7941 = _5293 & _7940;
    assign _7949 = _7941 ? _11940 : _7947;
    assign _7951 = _805 ? _4718 : _7949;
    assign _473 = _7951;
    always @(posedge _791) begin
        if (_789)
            _4081 <= _4718;
        else
            _4081 <= _473;
    end
    assign _7958 = _5304 == _2654;
    assign _7955 = ~ _3920;
    assign _7956 = _3135 & _7955;
    assign _7959 = _7956 & _7958;
    assign _7960 = _7959 ? _4693 : _4078;
    assign _7953 = _5296 == _2654;
    assign _7954 = _5293 & _7953;
    assign _7962 = _7954 ? _11940 : _7960;
    assign _7964 = _805 ? _4718 : _7962;
    assign _474 = _7964;
    always @(posedge _791) begin
        if (_789)
            _4078 <= _4718;
        else
            _4078 <= _474;
    end
    assign _7971 = _5304 == _2663;
    assign _7968 = ~ _3920;
    assign _7969 = _3135 & _7968;
    assign _7972 = _7969 & _7971;
    assign _7973 = _7972 ? _4693 : _4075;
    assign _7966 = _5296 == _2663;
    assign _7967 = _5293 & _7966;
    assign _7975 = _7967 ? _11940 : _7973;
    assign _7977 = _805 ? _4718 : _7975;
    assign _475 = _7977;
    always @(posedge _791) begin
        if (_789)
            _4075 <= _4718;
        else
            _4075 <= _475;
    end
    assign _7984 = _5304 == _2672;
    assign _7981 = ~ _3920;
    assign _7982 = _3135 & _7981;
    assign _7985 = _7982 & _7984;
    assign _7986 = _7985 ? _4693 : _4072;
    assign _7979 = _5296 == _2672;
    assign _7980 = _5293 & _7979;
    assign _7988 = _7980 ? _11940 : _7986;
    assign _7990 = _805 ? _4718 : _7988;
    assign _476 = _7990;
    always @(posedge _791) begin
        if (_789)
            _4072 <= _4718;
        else
            _4072 <= _476;
    end
    assign _7997 = _5304 == _2681;
    assign _7994 = ~ _3920;
    assign _7995 = _3135 & _7994;
    assign _7998 = _7995 & _7997;
    assign _7999 = _7998 ? _4693 : _4069;
    assign _7992 = _5296 == _2681;
    assign _7993 = _5293 & _7992;
    assign _8001 = _7993 ? _11940 : _7999;
    assign _8003 = _805 ? _4718 : _8001;
    assign _477 = _8003;
    always @(posedge _791) begin
        if (_789)
            _4069 <= _4718;
        else
            _4069 <= _477;
    end
    assign _8010 = _5304 == _2690;
    assign _8007 = ~ _3920;
    assign _8008 = _3135 & _8007;
    assign _8011 = _8008 & _8010;
    assign _8012 = _8011 ? _4693 : _4066;
    assign _8005 = _5296 == _2690;
    assign _8006 = _5293 & _8005;
    assign _8014 = _8006 ? _11940 : _8012;
    assign _8016 = _805 ? _4718 : _8014;
    assign _478 = _8016;
    always @(posedge _791) begin
        if (_789)
            _4066 <= _4718;
        else
            _4066 <= _478;
    end
    assign _8023 = _5304 == _2699;
    assign _8020 = ~ _3920;
    assign _8021 = _3135 & _8020;
    assign _8024 = _8021 & _8023;
    assign _8025 = _8024 ? _4693 : _4063;
    assign _8018 = _5296 == _2699;
    assign _8019 = _5293 & _8018;
    assign _8027 = _8019 ? _11940 : _8025;
    assign _8029 = _805 ? _4718 : _8027;
    assign _479 = _8029;
    always @(posedge _791) begin
        if (_789)
            _4063 <= _4718;
        else
            _4063 <= _479;
    end
    assign _8036 = _5304 == _2708;
    assign _8033 = ~ _3920;
    assign _8034 = _3135 & _8033;
    assign _8037 = _8034 & _8036;
    assign _8038 = _8037 ? _4693 : _4060;
    assign _8031 = _5296 == _2708;
    assign _8032 = _5293 & _8031;
    assign _8040 = _8032 ? _11940 : _8038;
    assign _8042 = _805 ? _4718 : _8040;
    assign _480 = _8042;
    always @(posedge _791) begin
        if (_789)
            _4060 <= _4718;
        else
            _4060 <= _480;
    end
    assign _8049 = _5304 == _2717;
    assign _8046 = ~ _3920;
    assign _8047 = _3135 & _8046;
    assign _8050 = _8047 & _8049;
    assign _8051 = _8050 ? _4693 : _4057;
    assign _8044 = _5296 == _2717;
    assign _8045 = _5293 & _8044;
    assign _8053 = _8045 ? _11940 : _8051;
    assign _8055 = _805 ? _4718 : _8053;
    assign _481 = _8055;
    always @(posedge _791) begin
        if (_789)
            _4057 <= _4718;
        else
            _4057 <= _481;
    end
    assign _8062 = _5304 == _2726;
    assign _8059 = ~ _3920;
    assign _8060 = _3135 & _8059;
    assign _8063 = _8060 & _8062;
    assign _8064 = _8063 ? _4693 : _4054;
    assign _8057 = _5296 == _2726;
    assign _8058 = _5293 & _8057;
    assign _8066 = _8058 ? _11940 : _8064;
    assign _8068 = _805 ? _4718 : _8066;
    assign _482 = _8068;
    always @(posedge _791) begin
        if (_789)
            _4054 <= _4718;
        else
            _4054 <= _482;
    end
    assign _8075 = _5304 == _2735;
    assign _8072 = ~ _3920;
    assign _8073 = _3135 & _8072;
    assign _8076 = _8073 & _8075;
    assign _8077 = _8076 ? _4693 : _4051;
    assign _8070 = _5296 == _2735;
    assign _8071 = _5293 & _8070;
    assign _8079 = _8071 ? _11940 : _8077;
    assign _8081 = _805 ? _4718 : _8079;
    assign _483 = _8081;
    always @(posedge _791) begin
        if (_789)
            _4051 <= _4718;
        else
            _4051 <= _483;
    end
    assign _8088 = _5304 == _2744;
    assign _8085 = ~ _3920;
    assign _8086 = _3135 & _8085;
    assign _8089 = _8086 & _8088;
    assign _8090 = _8089 ? _4693 : _4048;
    assign _8083 = _5296 == _2744;
    assign _8084 = _5293 & _8083;
    assign _8092 = _8084 ? _11940 : _8090;
    assign _8094 = _805 ? _4718 : _8092;
    assign _484 = _8094;
    always @(posedge _791) begin
        if (_789)
            _4048 <= _4718;
        else
            _4048 <= _484;
    end
    assign _8101 = _5304 == _2753;
    assign _8098 = ~ _3920;
    assign _8099 = _3135 & _8098;
    assign _8102 = _8099 & _8101;
    assign _8103 = _8102 ? _4693 : _4045;
    assign _8096 = _5296 == _2753;
    assign _8097 = _5293 & _8096;
    assign _8105 = _8097 ? _11940 : _8103;
    assign _8107 = _805 ? _4718 : _8105;
    assign _485 = _8107;
    always @(posedge _791) begin
        if (_789)
            _4045 <= _4718;
        else
            _4045 <= _485;
    end
    assign _8114 = _5304 == _2762;
    assign _8111 = ~ _3920;
    assign _8112 = _3135 & _8111;
    assign _8115 = _8112 & _8114;
    assign _8116 = _8115 ? _4693 : _4042;
    assign _8109 = _5296 == _2762;
    assign _8110 = _5293 & _8109;
    assign _8118 = _8110 ? _11940 : _8116;
    assign _8120 = _805 ? _4718 : _8118;
    assign _486 = _8120;
    always @(posedge _791) begin
        if (_789)
            _4042 <= _4718;
        else
            _4042 <= _486;
    end
    assign _8127 = _5304 == _2771;
    assign _8124 = ~ _3920;
    assign _8125 = _3135 & _8124;
    assign _8128 = _8125 & _8127;
    assign _8129 = _8128 ? _4693 : _4039;
    assign _8122 = _5296 == _2771;
    assign _8123 = _5293 & _8122;
    assign _8131 = _8123 ? _11940 : _8129;
    assign _8133 = _805 ? _4718 : _8131;
    assign _487 = _8133;
    always @(posedge _791) begin
        if (_789)
            _4039 <= _4718;
        else
            _4039 <= _487;
    end
    assign _8140 = _5304 == _2780;
    assign _8137 = ~ _3920;
    assign _8138 = _3135 & _8137;
    assign _8141 = _8138 & _8140;
    assign _8142 = _8141 ? _4693 : _4036;
    assign _8135 = _5296 == _2780;
    assign _8136 = _5293 & _8135;
    assign _8144 = _8136 ? _11940 : _8142;
    assign _8146 = _805 ? _4718 : _8144;
    assign _488 = _8146;
    always @(posedge _791) begin
        if (_789)
            _4036 <= _4718;
        else
            _4036 <= _488;
    end
    assign _8153 = _5304 == _2789;
    assign _8150 = ~ _3920;
    assign _8151 = _3135 & _8150;
    assign _8154 = _8151 & _8153;
    assign _8155 = _8154 ? _4693 : _4033;
    assign _8148 = _5296 == _2789;
    assign _8149 = _5293 & _8148;
    assign _8157 = _8149 ? _11940 : _8155;
    assign _8159 = _805 ? _4718 : _8157;
    assign _489 = _8159;
    always @(posedge _791) begin
        if (_789)
            _4033 <= _4718;
        else
            _4033 <= _489;
    end
    assign _8166 = _5304 == _2798;
    assign _8163 = ~ _3920;
    assign _8164 = _3135 & _8163;
    assign _8167 = _8164 & _8166;
    assign _8168 = _8167 ? _4693 : _4030;
    assign _8161 = _5296 == _2798;
    assign _8162 = _5293 & _8161;
    assign _8170 = _8162 ? _11940 : _8168;
    assign _8172 = _805 ? _4718 : _8170;
    assign _490 = _8172;
    always @(posedge _791) begin
        if (_789)
            _4030 <= _4718;
        else
            _4030 <= _490;
    end
    assign _8179 = _5304 == _2807;
    assign _8176 = ~ _3920;
    assign _8177 = _3135 & _8176;
    assign _8180 = _8177 & _8179;
    assign _8181 = _8180 ? _4693 : _4027;
    assign _8174 = _5296 == _2807;
    assign _8175 = _5293 & _8174;
    assign _8183 = _8175 ? _11940 : _8181;
    assign _8185 = _805 ? _4718 : _8183;
    assign _491 = _8185;
    always @(posedge _791) begin
        if (_789)
            _4027 <= _4718;
        else
            _4027 <= _491;
    end
    assign _8192 = _5304 == _2816;
    assign _8189 = ~ _3920;
    assign _8190 = _3135 & _8189;
    assign _8193 = _8190 & _8192;
    assign _8194 = _8193 ? _4693 : _4024;
    assign _8187 = _5296 == _2816;
    assign _8188 = _5293 & _8187;
    assign _8196 = _8188 ? _11940 : _8194;
    assign _8198 = _805 ? _4718 : _8196;
    assign _492 = _8198;
    always @(posedge _791) begin
        if (_789)
            _4024 <= _4718;
        else
            _4024 <= _492;
    end
    assign _8205 = _5304 == _2825;
    assign _8202 = ~ _3920;
    assign _8203 = _3135 & _8202;
    assign _8206 = _8203 & _8205;
    assign _8207 = _8206 ? _4693 : _4021;
    assign _8200 = _5296 == _2825;
    assign _8201 = _5293 & _8200;
    assign _8209 = _8201 ? _11940 : _8207;
    assign _8211 = _805 ? _4718 : _8209;
    assign _493 = _8211;
    always @(posedge _791) begin
        if (_789)
            _4021 <= _4718;
        else
            _4021 <= _493;
    end
    assign _8218 = _5304 == _2834;
    assign _8215 = ~ _3920;
    assign _8216 = _3135 & _8215;
    assign _8219 = _8216 & _8218;
    assign _8220 = _8219 ? _4693 : _4018;
    assign _8213 = _5296 == _2834;
    assign _8214 = _5293 & _8213;
    assign _8222 = _8214 ? _11940 : _8220;
    assign _8224 = _805 ? _4718 : _8222;
    assign _494 = _8224;
    always @(posedge _791) begin
        if (_789)
            _4018 <= _4718;
        else
            _4018 <= _494;
    end
    assign _8231 = _5304 == _2843;
    assign _8228 = ~ _3920;
    assign _8229 = _3135 & _8228;
    assign _8232 = _8229 & _8231;
    assign _8233 = _8232 ? _4693 : _4015;
    assign _8226 = _5296 == _2843;
    assign _8227 = _5293 & _8226;
    assign _8235 = _8227 ? _11940 : _8233;
    assign _8237 = _805 ? _4718 : _8235;
    assign _495 = _8237;
    always @(posedge _791) begin
        if (_789)
            _4015 <= _4718;
        else
            _4015 <= _495;
    end
    assign _8244 = _5304 == _2852;
    assign _8241 = ~ _3920;
    assign _8242 = _3135 & _8241;
    assign _8245 = _8242 & _8244;
    assign _8246 = _8245 ? _4693 : _4012;
    assign _8239 = _5296 == _2852;
    assign _8240 = _5293 & _8239;
    assign _8248 = _8240 ? _11940 : _8246;
    assign _8250 = _805 ? _4718 : _8248;
    assign _496 = _8250;
    always @(posedge _791) begin
        if (_789)
            _4012 <= _4718;
        else
            _4012 <= _496;
    end
    assign _8257 = _5304 == _2861;
    assign _8254 = ~ _3920;
    assign _8255 = _3135 & _8254;
    assign _8258 = _8255 & _8257;
    assign _8259 = _8258 ? _4693 : _4009;
    assign _8252 = _5296 == _2861;
    assign _8253 = _5293 & _8252;
    assign _8261 = _8253 ? _11940 : _8259;
    assign _8263 = _805 ? _4718 : _8261;
    assign _497 = _8263;
    always @(posedge _791) begin
        if (_789)
            _4009 <= _4718;
        else
            _4009 <= _497;
    end
    assign _8270 = _5304 == _2870;
    assign _8267 = ~ _3920;
    assign _8268 = _3135 & _8267;
    assign _8271 = _8268 & _8270;
    assign _8272 = _8271 ? _4693 : _4006;
    assign _8265 = _5296 == _2870;
    assign _8266 = _5293 & _8265;
    assign _8274 = _8266 ? _11940 : _8272;
    assign _8276 = _805 ? _4718 : _8274;
    assign _498 = _8276;
    always @(posedge _791) begin
        if (_789)
            _4006 <= _4718;
        else
            _4006 <= _498;
    end
    assign _8283 = _5304 == _2879;
    assign _8280 = ~ _3920;
    assign _8281 = _3135 & _8280;
    assign _8284 = _8281 & _8283;
    assign _8285 = _8284 ? _4693 : _4003;
    assign _8278 = _5296 == _2879;
    assign _8279 = _5293 & _8278;
    assign _8287 = _8279 ? _11940 : _8285;
    assign _8289 = _805 ? _4718 : _8287;
    assign _499 = _8289;
    always @(posedge _791) begin
        if (_789)
            _4003 <= _4718;
        else
            _4003 <= _499;
    end
    assign _8296 = _5304 == _2888;
    assign _8293 = ~ _3920;
    assign _8294 = _3135 & _8293;
    assign _8297 = _8294 & _8296;
    assign _8298 = _8297 ? _4693 : _4000;
    assign _8291 = _5296 == _2888;
    assign _8292 = _5293 & _8291;
    assign _8300 = _8292 ? _11940 : _8298;
    assign _8302 = _805 ? _4718 : _8300;
    assign _500 = _8302;
    always @(posedge _791) begin
        if (_789)
            _4000 <= _4718;
        else
            _4000 <= _500;
    end
    assign _8309 = _5304 == _2897;
    assign _8306 = ~ _3920;
    assign _8307 = _3135 & _8306;
    assign _8310 = _8307 & _8309;
    assign _8311 = _8310 ? _4693 : _3997;
    assign _8304 = _5296 == _2897;
    assign _8305 = _5293 & _8304;
    assign _8313 = _8305 ? _11940 : _8311;
    assign _8315 = _805 ? _4718 : _8313;
    assign _501 = _8315;
    always @(posedge _791) begin
        if (_789)
            _3997 <= _4718;
        else
            _3997 <= _501;
    end
    assign _8322 = _5304 == _2906;
    assign _8319 = ~ _3920;
    assign _8320 = _3135 & _8319;
    assign _8323 = _8320 & _8322;
    assign _8324 = _8323 ? _4693 : _3994;
    assign _8317 = _5296 == _2906;
    assign _8318 = _5293 & _8317;
    assign _8326 = _8318 ? _11940 : _8324;
    assign _8328 = _805 ? _4718 : _8326;
    assign _502 = _8328;
    always @(posedge _791) begin
        if (_789)
            _3994 <= _4718;
        else
            _3994 <= _502;
    end
    assign _8335 = _5304 == _2915;
    assign _8332 = ~ _3920;
    assign _8333 = _3135 & _8332;
    assign _8336 = _8333 & _8335;
    assign _8337 = _8336 ? _4693 : _3991;
    assign _8330 = _5296 == _2915;
    assign _8331 = _5293 & _8330;
    assign _8339 = _8331 ? _11940 : _8337;
    assign _8341 = _805 ? _4718 : _8339;
    assign _503 = _8341;
    always @(posedge _791) begin
        if (_789)
            _3991 <= _4718;
        else
            _3991 <= _503;
    end
    assign _8348 = _5304 == _2924;
    assign _8345 = ~ _3920;
    assign _8346 = _3135 & _8345;
    assign _8349 = _8346 & _8348;
    assign _8350 = _8349 ? _4693 : _3988;
    assign _8343 = _5296 == _2924;
    assign _8344 = _5293 & _8343;
    assign _8352 = _8344 ? _11940 : _8350;
    assign _8354 = _805 ? _4718 : _8352;
    assign _504 = _8354;
    always @(posedge _791) begin
        if (_789)
            _3988 <= _4718;
        else
            _3988 <= _504;
    end
    assign _8361 = _5304 == _2933;
    assign _8358 = ~ _3920;
    assign _8359 = _3135 & _8358;
    assign _8362 = _8359 & _8361;
    assign _8363 = _8362 ? _4693 : _3985;
    assign _8356 = _5296 == _2933;
    assign _8357 = _5293 & _8356;
    assign _8365 = _8357 ? _11940 : _8363;
    assign _8367 = _805 ? _4718 : _8365;
    assign _505 = _8367;
    always @(posedge _791) begin
        if (_789)
            _3985 <= _4718;
        else
            _3985 <= _505;
    end
    assign _8374 = _5304 == _2942;
    assign _8371 = ~ _3920;
    assign _8372 = _3135 & _8371;
    assign _8375 = _8372 & _8374;
    assign _8376 = _8375 ? _4693 : _3982;
    assign _8369 = _5296 == _2942;
    assign _8370 = _5293 & _8369;
    assign _8378 = _8370 ? _11940 : _8376;
    assign _8380 = _805 ? _4718 : _8378;
    assign _506 = _8380;
    always @(posedge _791) begin
        if (_789)
            _3982 <= _4718;
        else
            _3982 <= _506;
    end
    assign _8387 = _5304 == _2951;
    assign _8384 = ~ _3920;
    assign _8385 = _3135 & _8384;
    assign _8388 = _8385 & _8387;
    assign _8389 = _8388 ? _4693 : _3979;
    assign _8382 = _5296 == _2951;
    assign _8383 = _5293 & _8382;
    assign _8391 = _8383 ? _11940 : _8389;
    assign _8393 = _805 ? _4718 : _8391;
    assign _507 = _8393;
    always @(posedge _791) begin
        if (_789)
            _3979 <= _4718;
        else
            _3979 <= _507;
    end
    assign _8400 = _5304 == _2960;
    assign _8397 = ~ _3920;
    assign _8398 = _3135 & _8397;
    assign _8401 = _8398 & _8400;
    assign _8402 = _8401 ? _4693 : _3976;
    assign _8395 = _5296 == _2960;
    assign _8396 = _5293 & _8395;
    assign _8404 = _8396 ? _11940 : _8402;
    assign _8406 = _805 ? _4718 : _8404;
    assign _508 = _8406;
    always @(posedge _791) begin
        if (_789)
            _3976 <= _4718;
        else
            _3976 <= _508;
    end
    assign _8413 = _5304 == _2969;
    assign _8410 = ~ _3920;
    assign _8411 = _3135 & _8410;
    assign _8414 = _8411 & _8413;
    assign _8415 = _8414 ? _4693 : _3973;
    assign _8408 = _5296 == _2969;
    assign _8409 = _5293 & _8408;
    assign _8417 = _8409 ? _11940 : _8415;
    assign _8419 = _805 ? _4718 : _8417;
    assign _509 = _8419;
    always @(posedge _791) begin
        if (_789)
            _3973 <= _4718;
        else
            _3973 <= _509;
    end
    assign _8426 = _5304 == _2978;
    assign _8423 = ~ _3920;
    assign _8424 = _3135 & _8423;
    assign _8427 = _8424 & _8426;
    assign _8428 = _8427 ? _4693 : _3970;
    assign _8421 = _5296 == _2978;
    assign _8422 = _5293 & _8421;
    assign _8430 = _8422 ? _11940 : _8428;
    assign _8432 = _805 ? _4718 : _8430;
    assign _510 = _8432;
    always @(posedge _791) begin
        if (_789)
            _3970 <= _4718;
        else
            _3970 <= _510;
    end
    assign _8439 = _5304 == _2987;
    assign _8436 = ~ _3920;
    assign _8437 = _3135 & _8436;
    assign _8440 = _8437 & _8439;
    assign _8441 = _8440 ? _4693 : _3967;
    assign _8434 = _5296 == _2987;
    assign _8435 = _5293 & _8434;
    assign _8443 = _8435 ? _11940 : _8441;
    assign _8445 = _805 ? _4718 : _8443;
    assign _511 = _8445;
    always @(posedge _791) begin
        if (_789)
            _3967 <= _4718;
        else
            _3967 <= _511;
    end
    assign _8452 = _5304 == _2996;
    assign _8449 = ~ _3920;
    assign _8450 = _3135 & _8449;
    assign _8453 = _8450 & _8452;
    assign _8454 = _8453 ? _4693 : _3964;
    assign _8447 = _5296 == _2996;
    assign _8448 = _5293 & _8447;
    assign _8456 = _8448 ? _11940 : _8454;
    assign _8458 = _805 ? _4718 : _8456;
    assign _512 = _8458;
    always @(posedge _791) begin
        if (_789)
            _3964 <= _4718;
        else
            _3964 <= _512;
    end
    assign _8465 = _5304 == _3005;
    assign _8462 = ~ _3920;
    assign _8463 = _3135 & _8462;
    assign _8466 = _8463 & _8465;
    assign _8467 = _8466 ? _4693 : _3961;
    assign _8460 = _5296 == _3005;
    assign _8461 = _5293 & _8460;
    assign _8469 = _8461 ? _11940 : _8467;
    assign _8471 = _805 ? _4718 : _8469;
    assign _513 = _8471;
    always @(posedge _791) begin
        if (_789)
            _3961 <= _4718;
        else
            _3961 <= _513;
    end
    assign _8478 = _5304 == _3014;
    assign _8475 = ~ _3920;
    assign _8476 = _3135 & _8475;
    assign _8479 = _8476 & _8478;
    assign _8480 = _8479 ? _4693 : _3958;
    assign _8473 = _5296 == _3014;
    assign _8474 = _5293 & _8473;
    assign _8482 = _8474 ? _11940 : _8480;
    assign _8484 = _805 ? _4718 : _8482;
    assign _514 = _8484;
    always @(posedge _791) begin
        if (_789)
            _3958 <= _4718;
        else
            _3958 <= _514;
    end
    assign _8491 = _5304 == _3023;
    assign _8488 = ~ _3920;
    assign _8489 = _3135 & _8488;
    assign _8492 = _8489 & _8491;
    assign _8493 = _8492 ? _4693 : _3955;
    assign _8486 = _5296 == _3023;
    assign _8487 = _5293 & _8486;
    assign _8495 = _8487 ? _11940 : _8493;
    assign _8497 = _805 ? _4718 : _8495;
    assign _515 = _8497;
    always @(posedge _791) begin
        if (_789)
            _3955 <= _4718;
        else
            _3955 <= _515;
    end
    assign _8504 = _5304 == _3032;
    assign _8501 = ~ _3920;
    assign _8502 = _3135 & _8501;
    assign _8505 = _8502 & _8504;
    assign _8506 = _8505 ? _4693 : _3952;
    assign _8499 = _5296 == _3032;
    assign _8500 = _5293 & _8499;
    assign _8508 = _8500 ? _11940 : _8506;
    assign _8510 = _805 ? _4718 : _8508;
    assign _516 = _8510;
    always @(posedge _791) begin
        if (_789)
            _3952 <= _4718;
        else
            _3952 <= _516;
    end
    assign _8517 = _5304 == _3041;
    assign _8514 = ~ _3920;
    assign _8515 = _3135 & _8514;
    assign _8518 = _8515 & _8517;
    assign _8519 = _8518 ? _4693 : _3949;
    assign _8512 = _5296 == _3041;
    assign _8513 = _5293 & _8512;
    assign _8521 = _8513 ? _11940 : _8519;
    assign _8523 = _805 ? _4718 : _8521;
    assign _517 = _8523;
    always @(posedge _791) begin
        if (_789)
            _3949 <= _4718;
        else
            _3949 <= _517;
    end
    assign _8530 = _5304 == _3050;
    assign _8527 = ~ _3920;
    assign _8528 = _3135 & _8527;
    assign _8531 = _8528 & _8530;
    assign _8532 = _8531 ? _4693 : _3946;
    assign _8525 = _5296 == _3050;
    assign _8526 = _5293 & _8525;
    assign _8534 = _8526 ? _11940 : _8532;
    assign _8536 = _805 ? _4718 : _8534;
    assign _518 = _8536;
    always @(posedge _791) begin
        if (_789)
            _3946 <= _4718;
        else
            _3946 <= _518;
    end
    assign _8543 = _5304 == _3059;
    assign _8540 = ~ _3920;
    assign _8541 = _3135 & _8540;
    assign _8544 = _8541 & _8543;
    assign _8545 = _8544 ? _4693 : _3943;
    assign _8538 = _5296 == _3059;
    assign _8539 = _5293 & _8538;
    assign _8547 = _8539 ? _11940 : _8545;
    assign _8549 = _805 ? _4718 : _8547;
    assign _519 = _8549;
    always @(posedge _791) begin
        if (_789)
            _3943 <= _4718;
        else
            _3943 <= _519;
    end
    assign _8556 = _5304 == _3068;
    assign _8553 = ~ _3920;
    assign _8554 = _3135 & _8553;
    assign _8557 = _8554 & _8556;
    assign _8558 = _8557 ? _4693 : _3940;
    assign _8551 = _5296 == _3068;
    assign _8552 = _5293 & _8551;
    assign _8560 = _8552 ? _11940 : _8558;
    assign _8562 = _805 ? _4718 : _8560;
    assign _520 = _8562;
    always @(posedge _791) begin
        if (_789)
            _3940 <= _4718;
        else
            _3940 <= _520;
    end
    assign _8569 = _5304 == _3077;
    assign _8566 = ~ _3920;
    assign _8567 = _3135 & _8566;
    assign _8570 = _8567 & _8569;
    assign _8571 = _8570 ? _4693 : _3937;
    assign _8564 = _5296 == _3077;
    assign _8565 = _5293 & _8564;
    assign _8573 = _8565 ? _11940 : _8571;
    assign _8575 = _805 ? _4718 : _8573;
    assign _521 = _8575;
    always @(posedge _791) begin
        if (_789)
            _3937 <= _4718;
        else
            _3937 <= _521;
    end
    assign _8582 = _5304 == _3086;
    assign _8579 = ~ _3920;
    assign _8580 = _3135 & _8579;
    assign _8583 = _8580 & _8582;
    assign _8584 = _8583 ? _4693 : _3934;
    assign _8577 = _5296 == _3086;
    assign _8578 = _5293 & _8577;
    assign _8586 = _8578 ? _11940 : _8584;
    assign _8588 = _805 ? _4718 : _8586;
    assign _522 = _8588;
    always @(posedge _791) begin
        if (_789)
            _3934 <= _4718;
        else
            _3934 <= _522;
    end
    assign _8595 = _5304 == _3095;
    assign _8592 = ~ _3920;
    assign _8593 = _3135 & _8592;
    assign _8596 = _8593 & _8595;
    assign _8597 = _8596 ? _4693 : _3931;
    assign _8590 = _5296 == _3095;
    assign _8591 = _5293 & _8590;
    assign _8599 = _8591 ? _11940 : _8597;
    assign _8601 = _805 ? _4718 : _8599;
    assign _523 = _8601;
    always @(posedge _791) begin
        if (_789)
            _3931 <= _4718;
        else
            _3931 <= _523;
    end
    assign _8608 = _5304 == _3104;
    assign _8605 = ~ _3920;
    assign _8606 = _3135 & _8605;
    assign _8609 = _8606 & _8608;
    assign _8610 = _8609 ? _4693 : _3928;
    assign _8603 = _5296 == _3104;
    assign _8604 = _5293 & _8603;
    assign _8612 = _8604 ? _11940 : _8610;
    assign _8614 = _805 ? _4718 : _8612;
    assign _524 = _8614;
    always @(posedge _791) begin
        if (_789)
            _3928 <= _4718;
        else
            _3928 <= _524;
    end
    always @* begin
        case (_3919)
        0:
            _4692 <= _3925;
        1:
            _4692 <= _3928;
        2:
            _4692 <= _3931;
        3:
            _4692 <= _3934;
        4:
            _4692 <= _3937;
        5:
            _4692 <= _3940;
        6:
            _4692 <= _3943;
        7:
            _4692 <= _3946;
        8:
            _4692 <= _3949;
        9:
            _4692 <= _3952;
        10:
            _4692 <= _3955;
        11:
            _4692 <= _3958;
        12:
            _4692 <= _3961;
        13:
            _4692 <= _3964;
        14:
            _4692 <= _3967;
        15:
            _4692 <= _3970;
        16:
            _4692 <= _3973;
        17:
            _4692 <= _3976;
        18:
            _4692 <= _3979;
        19:
            _4692 <= _3982;
        20:
            _4692 <= _3985;
        21:
            _4692 <= _3988;
        22:
            _4692 <= _3991;
        23:
            _4692 <= _3994;
        24:
            _4692 <= _3997;
        25:
            _4692 <= _4000;
        26:
            _4692 <= _4003;
        27:
            _4692 <= _4006;
        28:
            _4692 <= _4009;
        29:
            _4692 <= _4012;
        30:
            _4692 <= _4015;
        31:
            _4692 <= _4018;
        32:
            _4692 <= _4021;
        33:
            _4692 <= _4024;
        34:
            _4692 <= _4027;
        35:
            _4692 <= _4030;
        36:
            _4692 <= _4033;
        37:
            _4692 <= _4036;
        38:
            _4692 <= _4039;
        39:
            _4692 <= _4042;
        40:
            _4692 <= _4045;
        41:
            _4692 <= _4048;
        42:
            _4692 <= _4051;
        43:
            _4692 <= _4054;
        44:
            _4692 <= _4057;
        45:
            _4692 <= _4060;
        46:
            _4692 <= _4063;
        47:
            _4692 <= _4066;
        48:
            _4692 <= _4069;
        49:
            _4692 <= _4072;
        50:
            _4692 <= _4075;
        51:
            _4692 <= _4078;
        52:
            _4692 <= _4081;
        53:
            _4692 <= _4084;
        54:
            _4692 <= _4087;
        55:
            _4692 <= _4090;
        56:
            _4692 <= _4093;
        57:
            _4692 <= _4096;
        58:
            _4692 <= _4099;
        59:
            _4692 <= _4102;
        60:
            _4692 <= _4105;
        61:
            _4692 <= _4108;
        62:
            _4692 <= _4111;
        63:
            _4692 <= _4114;
        64:
            _4692 <= _4117;
        65:
            _4692 <= _4120;
        66:
            _4692 <= _4123;
        67:
            _4692 <= _4126;
        68:
            _4692 <= _4129;
        69:
            _4692 <= _4132;
        70:
            _4692 <= _4135;
        71:
            _4692 <= _4138;
        72:
            _4692 <= _4141;
        73:
            _4692 <= _4144;
        74:
            _4692 <= _4147;
        75:
            _4692 <= _4150;
        76:
            _4692 <= _4153;
        77:
            _4692 <= _4156;
        78:
            _4692 <= _4159;
        79:
            _4692 <= _4162;
        80:
            _4692 <= _4165;
        81:
            _4692 <= _4168;
        82:
            _4692 <= _4171;
        83:
            _4692 <= _4174;
        84:
            _4692 <= _4177;
        85:
            _4692 <= _4180;
        86:
            _4692 <= _4183;
        87:
            _4692 <= _4186;
        88:
            _4692 <= _4189;
        89:
            _4692 <= _4192;
        90:
            _4692 <= _4195;
        91:
            _4692 <= _4198;
        92:
            _4692 <= _4201;
        93:
            _4692 <= _4204;
        94:
            _4692 <= _4207;
        95:
            _4692 <= _4210;
        96:
            _4692 <= _4213;
        97:
            _4692 <= _4216;
        98:
            _4692 <= _4219;
        99:
            _4692 <= _4222;
        100:
            _4692 <= _4225;
        101:
            _4692 <= _4228;
        102:
            _4692 <= _4231;
        103:
            _4692 <= _4234;
        104:
            _4692 <= _4237;
        105:
            _4692 <= _4240;
        106:
            _4692 <= _4243;
        107:
            _4692 <= _4246;
        108:
            _4692 <= _4249;
        109:
            _4692 <= _4252;
        110:
            _4692 <= _4255;
        111:
            _4692 <= _4258;
        112:
            _4692 <= _4261;
        113:
            _4692 <= _4264;
        114:
            _4692 <= _4267;
        115:
            _4692 <= _4270;
        116:
            _4692 <= _4273;
        117:
            _4692 <= _4276;
        118:
            _4692 <= _4279;
        119:
            _4692 <= _4282;
        120:
            _4692 <= _4285;
        121:
            _4692 <= _4288;
        122:
            _4692 <= _4291;
        123:
            _4692 <= _4294;
        124:
            _4692 <= _4297;
        125:
            _4692 <= _4300;
        126:
            _4692 <= _4303;
        127:
            _4692 <= _4306;
        128:
            _4692 <= _4309;
        129:
            _4692 <= _4312;
        130:
            _4692 <= _4315;
        131:
            _4692 <= _4318;
        132:
            _4692 <= _4321;
        133:
            _4692 <= _4324;
        134:
            _4692 <= _4327;
        135:
            _4692 <= _4330;
        136:
            _4692 <= _4333;
        137:
            _4692 <= _4336;
        138:
            _4692 <= _4339;
        139:
            _4692 <= _4342;
        140:
            _4692 <= _4345;
        141:
            _4692 <= _4348;
        142:
            _4692 <= _4351;
        143:
            _4692 <= _4354;
        144:
            _4692 <= _4357;
        145:
            _4692 <= _4360;
        146:
            _4692 <= _4363;
        147:
            _4692 <= _4366;
        148:
            _4692 <= _4369;
        149:
            _4692 <= _4372;
        150:
            _4692 <= _4375;
        151:
            _4692 <= _4378;
        152:
            _4692 <= _4381;
        153:
            _4692 <= _4384;
        154:
            _4692 <= _4387;
        155:
            _4692 <= _4390;
        156:
            _4692 <= _4393;
        157:
            _4692 <= _4396;
        158:
            _4692 <= _4399;
        159:
            _4692 <= _4402;
        160:
            _4692 <= _4405;
        161:
            _4692 <= _4408;
        162:
            _4692 <= _4411;
        163:
            _4692 <= _4414;
        164:
            _4692 <= _4417;
        165:
            _4692 <= _4420;
        166:
            _4692 <= _4423;
        167:
            _4692 <= _4426;
        168:
            _4692 <= _4429;
        169:
            _4692 <= _4432;
        170:
            _4692 <= _4435;
        171:
            _4692 <= _4438;
        172:
            _4692 <= _4441;
        173:
            _4692 <= _4444;
        174:
            _4692 <= _4447;
        175:
            _4692 <= _4450;
        176:
            _4692 <= _4453;
        177:
            _4692 <= _4456;
        178:
            _4692 <= _4459;
        179:
            _4692 <= _4462;
        180:
            _4692 <= _4465;
        181:
            _4692 <= _4468;
        182:
            _4692 <= _4471;
        183:
            _4692 <= _4474;
        184:
            _4692 <= _4477;
        185:
            _4692 <= _4480;
        186:
            _4692 <= _4483;
        187:
            _4692 <= _4486;
        188:
            _4692 <= _4489;
        189:
            _4692 <= _4492;
        190:
            _4692 <= _4495;
        191:
            _4692 <= _4498;
        192:
            _4692 <= _4501;
        193:
            _4692 <= _4504;
        194:
            _4692 <= _4507;
        195:
            _4692 <= _4510;
        196:
            _4692 <= _4513;
        197:
            _4692 <= _4516;
        198:
            _4692 <= _4519;
        199:
            _4692 <= _4522;
        200:
            _4692 <= _4525;
        201:
            _4692 <= _4528;
        202:
            _4692 <= _4531;
        203:
            _4692 <= _4534;
        204:
            _4692 <= _4537;
        205:
            _4692 <= _4540;
        206:
            _4692 <= _4543;
        207:
            _4692 <= _4546;
        208:
            _4692 <= _4549;
        209:
            _4692 <= _4552;
        210:
            _4692 <= _4555;
        211:
            _4692 <= _4558;
        212:
            _4692 <= _4561;
        213:
            _4692 <= _4564;
        214:
            _4692 <= _4567;
        215:
            _4692 <= _4570;
        216:
            _4692 <= _4573;
        217:
            _4692 <= _4576;
        218:
            _4692 <= _4579;
        219:
            _4692 <= _4582;
        220:
            _4692 <= _4585;
        221:
            _4692 <= _4588;
        222:
            _4692 <= _4591;
        223:
            _4692 <= _4594;
        224:
            _4692 <= _4597;
        225:
            _4692 <= _4600;
        226:
            _4692 <= _4603;
        227:
            _4692 <= _4606;
        228:
            _4692 <= _4609;
        229:
            _4692 <= _4612;
        230:
            _4692 <= _4615;
        231:
            _4692 <= _4618;
        232:
            _4692 <= _4621;
        233:
            _4692 <= _4624;
        234:
            _4692 <= _4627;
        235:
            _4692 <= _4630;
        236:
            _4692 <= _4633;
        237:
            _4692 <= _4636;
        238:
            _4692 <= _4639;
        239:
            _4692 <= _4642;
        240:
            _4692 <= _4645;
        241:
            _4692 <= _4648;
        242:
            _4692 <= _4651;
        243:
            _4692 <= _4654;
        244:
            _4692 <= _4657;
        245:
            _4692 <= _4660;
        246:
            _4692 <= _4663;
        247:
            _4692 <= _4666;
        248:
            _4692 <= _4669;
        249:
            _4692 <= _4672;
        250:
            _4692 <= _4675;
        251:
            _4692 <= _4678;
        252:
            _4692 <= _4681;
        253:
            _4692 <= _4684;
        254:
            _4692 <= _4687;
        default:
            _4692 <= _4690;
        endcase
    end
    assign _4693 = _4691 + _4692;
    assign _8622 = _8620 == _818;
    assign _8618 = ~ _3920;
    assign _8619 = _3135 & _8618;
    assign _8623 = _8619 & _8622;
    assign _8624 = _8623 ? _5304 : _3903;
    assign _8616 = _5296 == _818;
    assign _8617 = _5293 & _8616;
    assign _8626 = _8617 ? _818 : _8624;
    assign _8628 = _805 ? _3118 : _8626;
    assign _525 = _8628;
    always @(posedge _791) begin
        if (_789)
            _3903 <= _3118;
        else
            _3903 <= _525;
    end
    assign _8635 = _8620 == _827;
    assign _8632 = ~ _3920;
    assign _8633 = _3135 & _8632;
    assign _8636 = _8633 & _8635;
    assign _8637 = _8636 ? _5304 : _3900;
    assign _8630 = _5296 == _827;
    assign _8631 = _5293 & _8630;
    assign _8639 = _8631 ? _827 : _8637;
    assign _8641 = _805 ? _3118 : _8639;
    assign _526 = _8641;
    always @(posedge _791) begin
        if (_789)
            _3900 <= _3118;
        else
            _3900 <= _526;
    end
    assign _8648 = _8620 == _836;
    assign _8645 = ~ _3920;
    assign _8646 = _3135 & _8645;
    assign _8649 = _8646 & _8648;
    assign _8650 = _8649 ? _5304 : _3897;
    assign _8643 = _5296 == _836;
    assign _8644 = _5293 & _8643;
    assign _8652 = _8644 ? _836 : _8650;
    assign _8654 = _805 ? _3118 : _8652;
    assign _527 = _8654;
    always @(posedge _791) begin
        if (_789)
            _3897 <= _3118;
        else
            _3897 <= _527;
    end
    assign _8661 = _8620 == _845;
    assign _8658 = ~ _3920;
    assign _8659 = _3135 & _8658;
    assign _8662 = _8659 & _8661;
    assign _8663 = _8662 ? _5304 : _3894;
    assign _8656 = _5296 == _845;
    assign _8657 = _5293 & _8656;
    assign _8665 = _8657 ? _845 : _8663;
    assign _8667 = _805 ? _3118 : _8665;
    assign _528 = _8667;
    always @(posedge _791) begin
        if (_789)
            _3894 <= _3118;
        else
            _3894 <= _528;
    end
    assign _8674 = _8620 == _854;
    assign _8671 = ~ _3920;
    assign _8672 = _3135 & _8671;
    assign _8675 = _8672 & _8674;
    assign _8676 = _8675 ? _5304 : _3891;
    assign _8669 = _5296 == _854;
    assign _8670 = _5293 & _8669;
    assign _8678 = _8670 ? _854 : _8676;
    assign _8680 = _805 ? _3118 : _8678;
    assign _529 = _8680;
    always @(posedge _791) begin
        if (_789)
            _3891 <= _3118;
        else
            _3891 <= _529;
    end
    assign _8687 = _8620 == _863;
    assign _8684 = ~ _3920;
    assign _8685 = _3135 & _8684;
    assign _8688 = _8685 & _8687;
    assign _8689 = _8688 ? _5304 : _3888;
    assign _8682 = _5296 == _863;
    assign _8683 = _5293 & _8682;
    assign _8691 = _8683 ? _863 : _8689;
    assign _8693 = _805 ? _3118 : _8691;
    assign _530 = _8693;
    always @(posedge _791) begin
        if (_789)
            _3888 <= _3118;
        else
            _3888 <= _530;
    end
    assign _8700 = _8620 == _872;
    assign _8697 = ~ _3920;
    assign _8698 = _3135 & _8697;
    assign _8701 = _8698 & _8700;
    assign _8702 = _8701 ? _5304 : _3885;
    assign _8695 = _5296 == _872;
    assign _8696 = _5293 & _8695;
    assign _8704 = _8696 ? _872 : _8702;
    assign _8706 = _805 ? _3118 : _8704;
    assign _531 = _8706;
    always @(posedge _791) begin
        if (_789)
            _3885 <= _3118;
        else
            _3885 <= _531;
    end
    assign _8713 = _8620 == _881;
    assign _8710 = ~ _3920;
    assign _8711 = _3135 & _8710;
    assign _8714 = _8711 & _8713;
    assign _8715 = _8714 ? _5304 : _3882;
    assign _8708 = _5296 == _881;
    assign _8709 = _5293 & _8708;
    assign _8717 = _8709 ? _881 : _8715;
    assign _8719 = _805 ? _3118 : _8717;
    assign _532 = _8719;
    always @(posedge _791) begin
        if (_789)
            _3882 <= _3118;
        else
            _3882 <= _532;
    end
    assign _8726 = _8620 == _890;
    assign _8723 = ~ _3920;
    assign _8724 = _3135 & _8723;
    assign _8727 = _8724 & _8726;
    assign _8728 = _8727 ? _5304 : _3879;
    assign _8721 = _5296 == _890;
    assign _8722 = _5293 & _8721;
    assign _8730 = _8722 ? _890 : _8728;
    assign _8732 = _805 ? _3118 : _8730;
    assign _533 = _8732;
    always @(posedge _791) begin
        if (_789)
            _3879 <= _3118;
        else
            _3879 <= _533;
    end
    assign _8739 = _8620 == _899;
    assign _8736 = ~ _3920;
    assign _8737 = _3135 & _8736;
    assign _8740 = _8737 & _8739;
    assign _8741 = _8740 ? _5304 : _3876;
    assign _8734 = _5296 == _899;
    assign _8735 = _5293 & _8734;
    assign _8743 = _8735 ? _899 : _8741;
    assign _8745 = _805 ? _3118 : _8743;
    assign _534 = _8745;
    always @(posedge _791) begin
        if (_789)
            _3876 <= _3118;
        else
            _3876 <= _534;
    end
    assign _8752 = _8620 == _908;
    assign _8749 = ~ _3920;
    assign _8750 = _3135 & _8749;
    assign _8753 = _8750 & _8752;
    assign _8754 = _8753 ? _5304 : _3873;
    assign _8747 = _5296 == _908;
    assign _8748 = _5293 & _8747;
    assign _8756 = _8748 ? _908 : _8754;
    assign _8758 = _805 ? _3118 : _8756;
    assign _535 = _8758;
    always @(posedge _791) begin
        if (_789)
            _3873 <= _3118;
        else
            _3873 <= _535;
    end
    assign _8765 = _8620 == _917;
    assign _8762 = ~ _3920;
    assign _8763 = _3135 & _8762;
    assign _8766 = _8763 & _8765;
    assign _8767 = _8766 ? _5304 : _3870;
    assign _8760 = _5296 == _917;
    assign _8761 = _5293 & _8760;
    assign _8769 = _8761 ? _917 : _8767;
    assign _8771 = _805 ? _3118 : _8769;
    assign _536 = _8771;
    always @(posedge _791) begin
        if (_789)
            _3870 <= _3118;
        else
            _3870 <= _536;
    end
    assign _8778 = _8620 == _926;
    assign _8775 = ~ _3920;
    assign _8776 = _3135 & _8775;
    assign _8779 = _8776 & _8778;
    assign _8780 = _8779 ? _5304 : _3867;
    assign _8773 = _5296 == _926;
    assign _8774 = _5293 & _8773;
    assign _8782 = _8774 ? _926 : _8780;
    assign _8784 = _805 ? _3118 : _8782;
    assign _537 = _8784;
    always @(posedge _791) begin
        if (_789)
            _3867 <= _3118;
        else
            _3867 <= _537;
    end
    assign _8791 = _8620 == _935;
    assign _8788 = ~ _3920;
    assign _8789 = _3135 & _8788;
    assign _8792 = _8789 & _8791;
    assign _8793 = _8792 ? _5304 : _3864;
    assign _8786 = _5296 == _935;
    assign _8787 = _5293 & _8786;
    assign _8795 = _8787 ? _935 : _8793;
    assign _8797 = _805 ? _3118 : _8795;
    assign _538 = _8797;
    always @(posedge _791) begin
        if (_789)
            _3864 <= _3118;
        else
            _3864 <= _538;
    end
    assign _8804 = _8620 == _944;
    assign _8801 = ~ _3920;
    assign _8802 = _3135 & _8801;
    assign _8805 = _8802 & _8804;
    assign _8806 = _8805 ? _5304 : _3861;
    assign _8799 = _5296 == _944;
    assign _8800 = _5293 & _8799;
    assign _8808 = _8800 ? _944 : _8806;
    assign _8810 = _805 ? _3118 : _8808;
    assign _539 = _8810;
    always @(posedge _791) begin
        if (_789)
            _3861 <= _3118;
        else
            _3861 <= _539;
    end
    assign _8817 = _8620 == _953;
    assign _8814 = ~ _3920;
    assign _8815 = _3135 & _8814;
    assign _8818 = _8815 & _8817;
    assign _8819 = _8818 ? _5304 : _3858;
    assign _8812 = _5296 == _953;
    assign _8813 = _5293 & _8812;
    assign _8821 = _8813 ? _953 : _8819;
    assign _8823 = _805 ? _3118 : _8821;
    assign _540 = _8823;
    always @(posedge _791) begin
        if (_789)
            _3858 <= _3118;
        else
            _3858 <= _540;
    end
    assign _8830 = _8620 == _962;
    assign _8827 = ~ _3920;
    assign _8828 = _3135 & _8827;
    assign _8831 = _8828 & _8830;
    assign _8832 = _8831 ? _5304 : _3855;
    assign _8825 = _5296 == _962;
    assign _8826 = _5293 & _8825;
    assign _8834 = _8826 ? _962 : _8832;
    assign _8836 = _805 ? _3118 : _8834;
    assign _541 = _8836;
    always @(posedge _791) begin
        if (_789)
            _3855 <= _3118;
        else
            _3855 <= _541;
    end
    assign _8843 = _8620 == _971;
    assign _8840 = ~ _3920;
    assign _8841 = _3135 & _8840;
    assign _8844 = _8841 & _8843;
    assign _8845 = _8844 ? _5304 : _3852;
    assign _8838 = _5296 == _971;
    assign _8839 = _5293 & _8838;
    assign _8847 = _8839 ? _971 : _8845;
    assign _8849 = _805 ? _3118 : _8847;
    assign _542 = _8849;
    always @(posedge _791) begin
        if (_789)
            _3852 <= _3118;
        else
            _3852 <= _542;
    end
    assign _8856 = _8620 == _980;
    assign _8853 = ~ _3920;
    assign _8854 = _3135 & _8853;
    assign _8857 = _8854 & _8856;
    assign _8858 = _8857 ? _5304 : _3849;
    assign _8851 = _5296 == _980;
    assign _8852 = _5293 & _8851;
    assign _8860 = _8852 ? _980 : _8858;
    assign _8862 = _805 ? _3118 : _8860;
    assign _543 = _8862;
    always @(posedge _791) begin
        if (_789)
            _3849 <= _3118;
        else
            _3849 <= _543;
    end
    assign _8869 = _8620 == _989;
    assign _8866 = ~ _3920;
    assign _8867 = _3135 & _8866;
    assign _8870 = _8867 & _8869;
    assign _8871 = _8870 ? _5304 : _3846;
    assign _8864 = _5296 == _989;
    assign _8865 = _5293 & _8864;
    assign _8873 = _8865 ? _989 : _8871;
    assign _8875 = _805 ? _3118 : _8873;
    assign _544 = _8875;
    always @(posedge _791) begin
        if (_789)
            _3846 <= _3118;
        else
            _3846 <= _544;
    end
    assign _8882 = _8620 == _998;
    assign _8879 = ~ _3920;
    assign _8880 = _3135 & _8879;
    assign _8883 = _8880 & _8882;
    assign _8884 = _8883 ? _5304 : _3843;
    assign _8877 = _5296 == _998;
    assign _8878 = _5293 & _8877;
    assign _8886 = _8878 ? _998 : _8884;
    assign _8888 = _805 ? _3118 : _8886;
    assign _545 = _8888;
    always @(posedge _791) begin
        if (_789)
            _3843 <= _3118;
        else
            _3843 <= _545;
    end
    assign _8895 = _8620 == _1007;
    assign _8892 = ~ _3920;
    assign _8893 = _3135 & _8892;
    assign _8896 = _8893 & _8895;
    assign _8897 = _8896 ? _5304 : _3840;
    assign _8890 = _5296 == _1007;
    assign _8891 = _5293 & _8890;
    assign _8899 = _8891 ? _1007 : _8897;
    assign _8901 = _805 ? _3118 : _8899;
    assign _546 = _8901;
    always @(posedge _791) begin
        if (_789)
            _3840 <= _3118;
        else
            _3840 <= _546;
    end
    assign _8908 = _8620 == _1016;
    assign _8905 = ~ _3920;
    assign _8906 = _3135 & _8905;
    assign _8909 = _8906 & _8908;
    assign _8910 = _8909 ? _5304 : _3837;
    assign _8903 = _5296 == _1016;
    assign _8904 = _5293 & _8903;
    assign _8912 = _8904 ? _1016 : _8910;
    assign _8914 = _805 ? _3118 : _8912;
    assign _547 = _8914;
    always @(posedge _791) begin
        if (_789)
            _3837 <= _3118;
        else
            _3837 <= _547;
    end
    assign _8921 = _8620 == _1025;
    assign _8918 = ~ _3920;
    assign _8919 = _3135 & _8918;
    assign _8922 = _8919 & _8921;
    assign _8923 = _8922 ? _5304 : _3834;
    assign _8916 = _5296 == _1025;
    assign _8917 = _5293 & _8916;
    assign _8925 = _8917 ? _1025 : _8923;
    assign _8927 = _805 ? _3118 : _8925;
    assign _548 = _8927;
    always @(posedge _791) begin
        if (_789)
            _3834 <= _3118;
        else
            _3834 <= _548;
    end
    assign _8934 = _8620 == _1034;
    assign _8931 = ~ _3920;
    assign _8932 = _3135 & _8931;
    assign _8935 = _8932 & _8934;
    assign _8936 = _8935 ? _5304 : _3831;
    assign _8929 = _5296 == _1034;
    assign _8930 = _5293 & _8929;
    assign _8938 = _8930 ? _1034 : _8936;
    assign _8940 = _805 ? _3118 : _8938;
    assign _549 = _8940;
    always @(posedge _791) begin
        if (_789)
            _3831 <= _3118;
        else
            _3831 <= _549;
    end
    assign _8947 = _8620 == _1043;
    assign _8944 = ~ _3920;
    assign _8945 = _3135 & _8944;
    assign _8948 = _8945 & _8947;
    assign _8949 = _8948 ? _5304 : _3828;
    assign _8942 = _5296 == _1043;
    assign _8943 = _5293 & _8942;
    assign _8951 = _8943 ? _1043 : _8949;
    assign _8953 = _805 ? _3118 : _8951;
    assign _550 = _8953;
    always @(posedge _791) begin
        if (_789)
            _3828 <= _3118;
        else
            _3828 <= _550;
    end
    assign _8960 = _8620 == _1052;
    assign _8957 = ~ _3920;
    assign _8958 = _3135 & _8957;
    assign _8961 = _8958 & _8960;
    assign _8962 = _8961 ? _5304 : _3825;
    assign _8955 = _5296 == _1052;
    assign _8956 = _5293 & _8955;
    assign _8964 = _8956 ? _1052 : _8962;
    assign _8966 = _805 ? _3118 : _8964;
    assign _551 = _8966;
    always @(posedge _791) begin
        if (_789)
            _3825 <= _3118;
        else
            _3825 <= _551;
    end
    assign _8973 = _8620 == _1061;
    assign _8970 = ~ _3920;
    assign _8971 = _3135 & _8970;
    assign _8974 = _8971 & _8973;
    assign _8975 = _8974 ? _5304 : _3822;
    assign _8968 = _5296 == _1061;
    assign _8969 = _5293 & _8968;
    assign _8977 = _8969 ? _1061 : _8975;
    assign _8979 = _805 ? _3118 : _8977;
    assign _552 = _8979;
    always @(posedge _791) begin
        if (_789)
            _3822 <= _3118;
        else
            _3822 <= _552;
    end
    assign _8986 = _8620 == _1070;
    assign _8983 = ~ _3920;
    assign _8984 = _3135 & _8983;
    assign _8987 = _8984 & _8986;
    assign _8988 = _8987 ? _5304 : _3819;
    assign _8981 = _5296 == _1070;
    assign _8982 = _5293 & _8981;
    assign _8990 = _8982 ? _1070 : _8988;
    assign _8992 = _805 ? _3118 : _8990;
    assign _553 = _8992;
    always @(posedge _791) begin
        if (_789)
            _3819 <= _3118;
        else
            _3819 <= _553;
    end
    assign _8999 = _8620 == _1079;
    assign _8996 = ~ _3920;
    assign _8997 = _3135 & _8996;
    assign _9000 = _8997 & _8999;
    assign _9001 = _9000 ? _5304 : _3816;
    assign _8994 = _5296 == _1079;
    assign _8995 = _5293 & _8994;
    assign _9003 = _8995 ? _1079 : _9001;
    assign _9005 = _805 ? _3118 : _9003;
    assign _554 = _9005;
    always @(posedge _791) begin
        if (_789)
            _3816 <= _3118;
        else
            _3816 <= _554;
    end
    assign _9012 = _8620 == _1088;
    assign _9009 = ~ _3920;
    assign _9010 = _3135 & _9009;
    assign _9013 = _9010 & _9012;
    assign _9014 = _9013 ? _5304 : _3813;
    assign _9007 = _5296 == _1088;
    assign _9008 = _5293 & _9007;
    assign _9016 = _9008 ? _1088 : _9014;
    assign _9018 = _805 ? _3118 : _9016;
    assign _555 = _9018;
    always @(posedge _791) begin
        if (_789)
            _3813 <= _3118;
        else
            _3813 <= _555;
    end
    assign _9025 = _8620 == _1097;
    assign _9022 = ~ _3920;
    assign _9023 = _3135 & _9022;
    assign _9026 = _9023 & _9025;
    assign _9027 = _9026 ? _5304 : _3810;
    assign _9020 = _5296 == _1097;
    assign _9021 = _5293 & _9020;
    assign _9029 = _9021 ? _1097 : _9027;
    assign _9031 = _805 ? _3118 : _9029;
    assign _556 = _9031;
    always @(posedge _791) begin
        if (_789)
            _3810 <= _3118;
        else
            _3810 <= _556;
    end
    assign _9038 = _8620 == _1106;
    assign _9035 = ~ _3920;
    assign _9036 = _3135 & _9035;
    assign _9039 = _9036 & _9038;
    assign _9040 = _9039 ? _5304 : _3807;
    assign _9033 = _5296 == _1106;
    assign _9034 = _5293 & _9033;
    assign _9042 = _9034 ? _1106 : _9040;
    assign _9044 = _805 ? _3118 : _9042;
    assign _557 = _9044;
    always @(posedge _791) begin
        if (_789)
            _3807 <= _3118;
        else
            _3807 <= _557;
    end
    assign _9051 = _8620 == _1115;
    assign _9048 = ~ _3920;
    assign _9049 = _3135 & _9048;
    assign _9052 = _9049 & _9051;
    assign _9053 = _9052 ? _5304 : _3804;
    assign _9046 = _5296 == _1115;
    assign _9047 = _5293 & _9046;
    assign _9055 = _9047 ? _1115 : _9053;
    assign _9057 = _805 ? _3118 : _9055;
    assign _558 = _9057;
    always @(posedge _791) begin
        if (_789)
            _3804 <= _3118;
        else
            _3804 <= _558;
    end
    assign _9064 = _8620 == _1124;
    assign _9061 = ~ _3920;
    assign _9062 = _3135 & _9061;
    assign _9065 = _9062 & _9064;
    assign _9066 = _9065 ? _5304 : _3801;
    assign _9059 = _5296 == _1124;
    assign _9060 = _5293 & _9059;
    assign _9068 = _9060 ? _1124 : _9066;
    assign _9070 = _805 ? _3118 : _9068;
    assign _559 = _9070;
    always @(posedge _791) begin
        if (_789)
            _3801 <= _3118;
        else
            _3801 <= _559;
    end
    assign _9077 = _8620 == _1133;
    assign _9074 = ~ _3920;
    assign _9075 = _3135 & _9074;
    assign _9078 = _9075 & _9077;
    assign _9079 = _9078 ? _5304 : _3798;
    assign _9072 = _5296 == _1133;
    assign _9073 = _5293 & _9072;
    assign _9081 = _9073 ? _1133 : _9079;
    assign _9083 = _805 ? _3118 : _9081;
    assign _560 = _9083;
    always @(posedge _791) begin
        if (_789)
            _3798 <= _3118;
        else
            _3798 <= _560;
    end
    assign _9090 = _8620 == _1142;
    assign _9087 = ~ _3920;
    assign _9088 = _3135 & _9087;
    assign _9091 = _9088 & _9090;
    assign _9092 = _9091 ? _5304 : _3795;
    assign _9085 = _5296 == _1142;
    assign _9086 = _5293 & _9085;
    assign _9094 = _9086 ? _1142 : _9092;
    assign _9096 = _805 ? _3118 : _9094;
    assign _561 = _9096;
    always @(posedge _791) begin
        if (_789)
            _3795 <= _3118;
        else
            _3795 <= _561;
    end
    assign _9103 = _8620 == _1151;
    assign _9100 = ~ _3920;
    assign _9101 = _3135 & _9100;
    assign _9104 = _9101 & _9103;
    assign _9105 = _9104 ? _5304 : _3792;
    assign _9098 = _5296 == _1151;
    assign _9099 = _5293 & _9098;
    assign _9107 = _9099 ? _1151 : _9105;
    assign _9109 = _805 ? _3118 : _9107;
    assign _562 = _9109;
    always @(posedge _791) begin
        if (_789)
            _3792 <= _3118;
        else
            _3792 <= _562;
    end
    assign _9116 = _8620 == _1160;
    assign _9113 = ~ _3920;
    assign _9114 = _3135 & _9113;
    assign _9117 = _9114 & _9116;
    assign _9118 = _9117 ? _5304 : _3789;
    assign _9111 = _5296 == _1160;
    assign _9112 = _5293 & _9111;
    assign _9120 = _9112 ? _1160 : _9118;
    assign _9122 = _805 ? _3118 : _9120;
    assign _563 = _9122;
    always @(posedge _791) begin
        if (_789)
            _3789 <= _3118;
        else
            _3789 <= _563;
    end
    assign _9129 = _8620 == _1169;
    assign _9126 = ~ _3920;
    assign _9127 = _3135 & _9126;
    assign _9130 = _9127 & _9129;
    assign _9131 = _9130 ? _5304 : _3786;
    assign _9124 = _5296 == _1169;
    assign _9125 = _5293 & _9124;
    assign _9133 = _9125 ? _1169 : _9131;
    assign _9135 = _805 ? _3118 : _9133;
    assign _564 = _9135;
    always @(posedge _791) begin
        if (_789)
            _3786 <= _3118;
        else
            _3786 <= _564;
    end
    assign _9142 = _8620 == _1178;
    assign _9139 = ~ _3920;
    assign _9140 = _3135 & _9139;
    assign _9143 = _9140 & _9142;
    assign _9144 = _9143 ? _5304 : _3783;
    assign _9137 = _5296 == _1178;
    assign _9138 = _5293 & _9137;
    assign _9146 = _9138 ? _1178 : _9144;
    assign _9148 = _805 ? _3118 : _9146;
    assign _565 = _9148;
    always @(posedge _791) begin
        if (_789)
            _3783 <= _3118;
        else
            _3783 <= _565;
    end
    assign _9155 = _8620 == _1187;
    assign _9152 = ~ _3920;
    assign _9153 = _3135 & _9152;
    assign _9156 = _9153 & _9155;
    assign _9157 = _9156 ? _5304 : _3780;
    assign _9150 = _5296 == _1187;
    assign _9151 = _5293 & _9150;
    assign _9159 = _9151 ? _1187 : _9157;
    assign _9161 = _805 ? _3118 : _9159;
    assign _566 = _9161;
    always @(posedge _791) begin
        if (_789)
            _3780 <= _3118;
        else
            _3780 <= _566;
    end
    assign _9168 = _8620 == _1196;
    assign _9165 = ~ _3920;
    assign _9166 = _3135 & _9165;
    assign _9169 = _9166 & _9168;
    assign _9170 = _9169 ? _5304 : _3777;
    assign _9163 = _5296 == _1196;
    assign _9164 = _5293 & _9163;
    assign _9172 = _9164 ? _1196 : _9170;
    assign _9174 = _805 ? _3118 : _9172;
    assign _567 = _9174;
    always @(posedge _791) begin
        if (_789)
            _3777 <= _3118;
        else
            _3777 <= _567;
    end
    assign _9181 = _8620 == _1205;
    assign _9178 = ~ _3920;
    assign _9179 = _3135 & _9178;
    assign _9182 = _9179 & _9181;
    assign _9183 = _9182 ? _5304 : _3774;
    assign _9176 = _5296 == _1205;
    assign _9177 = _5293 & _9176;
    assign _9185 = _9177 ? _1205 : _9183;
    assign _9187 = _805 ? _3118 : _9185;
    assign _568 = _9187;
    always @(posedge _791) begin
        if (_789)
            _3774 <= _3118;
        else
            _3774 <= _568;
    end
    assign _9194 = _8620 == _1214;
    assign _9191 = ~ _3920;
    assign _9192 = _3135 & _9191;
    assign _9195 = _9192 & _9194;
    assign _9196 = _9195 ? _5304 : _3771;
    assign _9189 = _5296 == _1214;
    assign _9190 = _5293 & _9189;
    assign _9198 = _9190 ? _1214 : _9196;
    assign _9200 = _805 ? _3118 : _9198;
    assign _569 = _9200;
    always @(posedge _791) begin
        if (_789)
            _3771 <= _3118;
        else
            _3771 <= _569;
    end
    assign _9207 = _8620 == _1223;
    assign _9204 = ~ _3920;
    assign _9205 = _3135 & _9204;
    assign _9208 = _9205 & _9207;
    assign _9209 = _9208 ? _5304 : _3768;
    assign _9202 = _5296 == _1223;
    assign _9203 = _5293 & _9202;
    assign _9211 = _9203 ? _1223 : _9209;
    assign _9213 = _805 ? _3118 : _9211;
    assign _570 = _9213;
    always @(posedge _791) begin
        if (_789)
            _3768 <= _3118;
        else
            _3768 <= _570;
    end
    assign _9220 = _8620 == _1232;
    assign _9217 = ~ _3920;
    assign _9218 = _3135 & _9217;
    assign _9221 = _9218 & _9220;
    assign _9222 = _9221 ? _5304 : _3765;
    assign _9215 = _5296 == _1232;
    assign _9216 = _5293 & _9215;
    assign _9224 = _9216 ? _1232 : _9222;
    assign _9226 = _805 ? _3118 : _9224;
    assign _571 = _9226;
    always @(posedge _791) begin
        if (_789)
            _3765 <= _3118;
        else
            _3765 <= _571;
    end
    assign _9233 = _8620 == _1241;
    assign _9230 = ~ _3920;
    assign _9231 = _3135 & _9230;
    assign _9234 = _9231 & _9233;
    assign _9235 = _9234 ? _5304 : _3762;
    assign _9228 = _5296 == _1241;
    assign _9229 = _5293 & _9228;
    assign _9237 = _9229 ? _1241 : _9235;
    assign _9239 = _805 ? _3118 : _9237;
    assign _572 = _9239;
    always @(posedge _791) begin
        if (_789)
            _3762 <= _3118;
        else
            _3762 <= _572;
    end
    assign _9246 = _8620 == _1250;
    assign _9243 = ~ _3920;
    assign _9244 = _3135 & _9243;
    assign _9247 = _9244 & _9246;
    assign _9248 = _9247 ? _5304 : _3759;
    assign _9241 = _5296 == _1250;
    assign _9242 = _5293 & _9241;
    assign _9250 = _9242 ? _1250 : _9248;
    assign _9252 = _805 ? _3118 : _9250;
    assign _573 = _9252;
    always @(posedge _791) begin
        if (_789)
            _3759 <= _3118;
        else
            _3759 <= _573;
    end
    assign _9259 = _8620 == _1259;
    assign _9256 = ~ _3920;
    assign _9257 = _3135 & _9256;
    assign _9260 = _9257 & _9259;
    assign _9261 = _9260 ? _5304 : _3756;
    assign _9254 = _5296 == _1259;
    assign _9255 = _5293 & _9254;
    assign _9263 = _9255 ? _1259 : _9261;
    assign _9265 = _805 ? _3118 : _9263;
    assign _574 = _9265;
    always @(posedge _791) begin
        if (_789)
            _3756 <= _3118;
        else
            _3756 <= _574;
    end
    assign _9272 = _8620 == _1268;
    assign _9269 = ~ _3920;
    assign _9270 = _3135 & _9269;
    assign _9273 = _9270 & _9272;
    assign _9274 = _9273 ? _5304 : _3753;
    assign _9267 = _5296 == _1268;
    assign _9268 = _5293 & _9267;
    assign _9276 = _9268 ? _1268 : _9274;
    assign _9278 = _805 ? _3118 : _9276;
    assign _575 = _9278;
    always @(posedge _791) begin
        if (_789)
            _3753 <= _3118;
        else
            _3753 <= _575;
    end
    assign _9285 = _8620 == _1277;
    assign _9282 = ~ _3920;
    assign _9283 = _3135 & _9282;
    assign _9286 = _9283 & _9285;
    assign _9287 = _9286 ? _5304 : _3750;
    assign _9280 = _5296 == _1277;
    assign _9281 = _5293 & _9280;
    assign _9289 = _9281 ? _1277 : _9287;
    assign _9291 = _805 ? _3118 : _9289;
    assign _576 = _9291;
    always @(posedge _791) begin
        if (_789)
            _3750 <= _3118;
        else
            _3750 <= _576;
    end
    assign _9298 = _8620 == _1286;
    assign _9295 = ~ _3920;
    assign _9296 = _3135 & _9295;
    assign _9299 = _9296 & _9298;
    assign _9300 = _9299 ? _5304 : _3747;
    assign _9293 = _5296 == _1286;
    assign _9294 = _5293 & _9293;
    assign _9302 = _9294 ? _1286 : _9300;
    assign _9304 = _805 ? _3118 : _9302;
    assign _577 = _9304;
    always @(posedge _791) begin
        if (_789)
            _3747 <= _3118;
        else
            _3747 <= _577;
    end
    assign _9311 = _8620 == _1295;
    assign _9308 = ~ _3920;
    assign _9309 = _3135 & _9308;
    assign _9312 = _9309 & _9311;
    assign _9313 = _9312 ? _5304 : _3744;
    assign _9306 = _5296 == _1295;
    assign _9307 = _5293 & _9306;
    assign _9315 = _9307 ? _1295 : _9313;
    assign _9317 = _805 ? _3118 : _9315;
    assign _578 = _9317;
    always @(posedge _791) begin
        if (_789)
            _3744 <= _3118;
        else
            _3744 <= _578;
    end
    assign _9324 = _8620 == _1304;
    assign _9321 = ~ _3920;
    assign _9322 = _3135 & _9321;
    assign _9325 = _9322 & _9324;
    assign _9326 = _9325 ? _5304 : _3741;
    assign _9319 = _5296 == _1304;
    assign _9320 = _5293 & _9319;
    assign _9328 = _9320 ? _1304 : _9326;
    assign _9330 = _805 ? _3118 : _9328;
    assign _579 = _9330;
    always @(posedge _791) begin
        if (_789)
            _3741 <= _3118;
        else
            _3741 <= _579;
    end
    assign _9337 = _8620 == _1313;
    assign _9334 = ~ _3920;
    assign _9335 = _3135 & _9334;
    assign _9338 = _9335 & _9337;
    assign _9339 = _9338 ? _5304 : _3738;
    assign _9332 = _5296 == _1313;
    assign _9333 = _5293 & _9332;
    assign _9341 = _9333 ? _1313 : _9339;
    assign _9343 = _805 ? _3118 : _9341;
    assign _580 = _9343;
    always @(posedge _791) begin
        if (_789)
            _3738 <= _3118;
        else
            _3738 <= _580;
    end
    assign _9350 = _8620 == _1322;
    assign _9347 = ~ _3920;
    assign _9348 = _3135 & _9347;
    assign _9351 = _9348 & _9350;
    assign _9352 = _9351 ? _5304 : _3735;
    assign _9345 = _5296 == _1322;
    assign _9346 = _5293 & _9345;
    assign _9354 = _9346 ? _1322 : _9352;
    assign _9356 = _805 ? _3118 : _9354;
    assign _581 = _9356;
    always @(posedge _791) begin
        if (_789)
            _3735 <= _3118;
        else
            _3735 <= _581;
    end
    assign _9363 = _8620 == _1331;
    assign _9360 = ~ _3920;
    assign _9361 = _3135 & _9360;
    assign _9364 = _9361 & _9363;
    assign _9365 = _9364 ? _5304 : _3732;
    assign _9358 = _5296 == _1331;
    assign _9359 = _5293 & _9358;
    assign _9367 = _9359 ? _1331 : _9365;
    assign _9369 = _805 ? _3118 : _9367;
    assign _582 = _9369;
    always @(posedge _791) begin
        if (_789)
            _3732 <= _3118;
        else
            _3732 <= _582;
    end
    assign _9376 = _8620 == _1340;
    assign _9373 = ~ _3920;
    assign _9374 = _3135 & _9373;
    assign _9377 = _9374 & _9376;
    assign _9378 = _9377 ? _5304 : _3729;
    assign _9371 = _5296 == _1340;
    assign _9372 = _5293 & _9371;
    assign _9380 = _9372 ? _1340 : _9378;
    assign _9382 = _805 ? _3118 : _9380;
    assign _583 = _9382;
    always @(posedge _791) begin
        if (_789)
            _3729 <= _3118;
        else
            _3729 <= _583;
    end
    assign _9389 = _8620 == _1349;
    assign _9386 = ~ _3920;
    assign _9387 = _3135 & _9386;
    assign _9390 = _9387 & _9389;
    assign _9391 = _9390 ? _5304 : _3726;
    assign _9384 = _5296 == _1349;
    assign _9385 = _5293 & _9384;
    assign _9393 = _9385 ? _1349 : _9391;
    assign _9395 = _805 ? _3118 : _9393;
    assign _584 = _9395;
    always @(posedge _791) begin
        if (_789)
            _3726 <= _3118;
        else
            _3726 <= _584;
    end
    assign _9402 = _8620 == _1358;
    assign _9399 = ~ _3920;
    assign _9400 = _3135 & _9399;
    assign _9403 = _9400 & _9402;
    assign _9404 = _9403 ? _5304 : _3723;
    assign _9397 = _5296 == _1358;
    assign _9398 = _5293 & _9397;
    assign _9406 = _9398 ? _1358 : _9404;
    assign _9408 = _805 ? _3118 : _9406;
    assign _585 = _9408;
    always @(posedge _791) begin
        if (_789)
            _3723 <= _3118;
        else
            _3723 <= _585;
    end
    assign _9415 = _8620 == _1367;
    assign _9412 = ~ _3920;
    assign _9413 = _3135 & _9412;
    assign _9416 = _9413 & _9415;
    assign _9417 = _9416 ? _5304 : _3720;
    assign _9410 = _5296 == _1367;
    assign _9411 = _5293 & _9410;
    assign _9419 = _9411 ? _1367 : _9417;
    assign _9421 = _805 ? _3118 : _9419;
    assign _586 = _9421;
    always @(posedge _791) begin
        if (_789)
            _3720 <= _3118;
        else
            _3720 <= _586;
    end
    assign _9428 = _8620 == _1376;
    assign _9425 = ~ _3920;
    assign _9426 = _3135 & _9425;
    assign _9429 = _9426 & _9428;
    assign _9430 = _9429 ? _5304 : _3717;
    assign _9423 = _5296 == _1376;
    assign _9424 = _5293 & _9423;
    assign _9432 = _9424 ? _1376 : _9430;
    assign _9434 = _805 ? _3118 : _9432;
    assign _587 = _9434;
    always @(posedge _791) begin
        if (_789)
            _3717 <= _3118;
        else
            _3717 <= _587;
    end
    assign _9441 = _8620 == _1385;
    assign _9438 = ~ _3920;
    assign _9439 = _3135 & _9438;
    assign _9442 = _9439 & _9441;
    assign _9443 = _9442 ? _5304 : _3714;
    assign _9436 = _5296 == _1385;
    assign _9437 = _5293 & _9436;
    assign _9445 = _9437 ? _1385 : _9443;
    assign _9447 = _805 ? _3118 : _9445;
    assign _588 = _9447;
    always @(posedge _791) begin
        if (_789)
            _3714 <= _3118;
        else
            _3714 <= _588;
    end
    assign _9454 = _8620 == _1394;
    assign _9451 = ~ _3920;
    assign _9452 = _3135 & _9451;
    assign _9455 = _9452 & _9454;
    assign _9456 = _9455 ? _5304 : _3711;
    assign _9449 = _5296 == _1394;
    assign _9450 = _5293 & _9449;
    assign _9458 = _9450 ? _1394 : _9456;
    assign _9460 = _805 ? _3118 : _9458;
    assign _589 = _9460;
    always @(posedge _791) begin
        if (_789)
            _3711 <= _3118;
        else
            _3711 <= _589;
    end
    assign _9467 = _8620 == _1403;
    assign _9464 = ~ _3920;
    assign _9465 = _3135 & _9464;
    assign _9468 = _9465 & _9467;
    assign _9469 = _9468 ? _5304 : _3708;
    assign _9462 = _5296 == _1403;
    assign _9463 = _5293 & _9462;
    assign _9471 = _9463 ? _1403 : _9469;
    assign _9473 = _805 ? _3118 : _9471;
    assign _590 = _9473;
    always @(posedge _791) begin
        if (_789)
            _3708 <= _3118;
        else
            _3708 <= _590;
    end
    assign _9480 = _8620 == _1412;
    assign _9477 = ~ _3920;
    assign _9478 = _3135 & _9477;
    assign _9481 = _9478 & _9480;
    assign _9482 = _9481 ? _5304 : _3705;
    assign _9475 = _5296 == _1412;
    assign _9476 = _5293 & _9475;
    assign _9484 = _9476 ? _1412 : _9482;
    assign _9486 = _805 ? _3118 : _9484;
    assign _591 = _9486;
    always @(posedge _791) begin
        if (_789)
            _3705 <= _3118;
        else
            _3705 <= _591;
    end
    assign _9493 = _8620 == _1421;
    assign _9490 = ~ _3920;
    assign _9491 = _3135 & _9490;
    assign _9494 = _9491 & _9493;
    assign _9495 = _9494 ? _5304 : _3702;
    assign _9488 = _5296 == _1421;
    assign _9489 = _5293 & _9488;
    assign _9497 = _9489 ? _1421 : _9495;
    assign _9499 = _805 ? _3118 : _9497;
    assign _592 = _9499;
    always @(posedge _791) begin
        if (_789)
            _3702 <= _3118;
        else
            _3702 <= _592;
    end
    assign _9506 = _8620 == _1430;
    assign _9503 = ~ _3920;
    assign _9504 = _3135 & _9503;
    assign _9507 = _9504 & _9506;
    assign _9508 = _9507 ? _5304 : _3699;
    assign _9501 = _5296 == _1430;
    assign _9502 = _5293 & _9501;
    assign _9510 = _9502 ? _1430 : _9508;
    assign _9512 = _805 ? _3118 : _9510;
    assign _593 = _9512;
    always @(posedge _791) begin
        if (_789)
            _3699 <= _3118;
        else
            _3699 <= _593;
    end
    assign _9519 = _8620 == _1439;
    assign _9516 = ~ _3920;
    assign _9517 = _3135 & _9516;
    assign _9520 = _9517 & _9519;
    assign _9521 = _9520 ? _5304 : _3696;
    assign _9514 = _5296 == _1439;
    assign _9515 = _5293 & _9514;
    assign _9523 = _9515 ? _1439 : _9521;
    assign _9525 = _805 ? _3118 : _9523;
    assign _594 = _9525;
    always @(posedge _791) begin
        if (_789)
            _3696 <= _3118;
        else
            _3696 <= _594;
    end
    assign _9532 = _8620 == _1448;
    assign _9529 = ~ _3920;
    assign _9530 = _3135 & _9529;
    assign _9533 = _9530 & _9532;
    assign _9534 = _9533 ? _5304 : _3693;
    assign _9527 = _5296 == _1448;
    assign _9528 = _5293 & _9527;
    assign _9536 = _9528 ? _1448 : _9534;
    assign _9538 = _805 ? _3118 : _9536;
    assign _595 = _9538;
    always @(posedge _791) begin
        if (_789)
            _3693 <= _3118;
        else
            _3693 <= _595;
    end
    assign _9545 = _8620 == _1457;
    assign _9542 = ~ _3920;
    assign _9543 = _3135 & _9542;
    assign _9546 = _9543 & _9545;
    assign _9547 = _9546 ? _5304 : _3690;
    assign _9540 = _5296 == _1457;
    assign _9541 = _5293 & _9540;
    assign _9549 = _9541 ? _1457 : _9547;
    assign _9551 = _805 ? _3118 : _9549;
    assign _596 = _9551;
    always @(posedge _791) begin
        if (_789)
            _3690 <= _3118;
        else
            _3690 <= _596;
    end
    assign _9558 = _8620 == _1466;
    assign _9555 = ~ _3920;
    assign _9556 = _3135 & _9555;
    assign _9559 = _9556 & _9558;
    assign _9560 = _9559 ? _5304 : _3687;
    assign _9553 = _5296 == _1466;
    assign _9554 = _5293 & _9553;
    assign _9562 = _9554 ? _1466 : _9560;
    assign _9564 = _805 ? _3118 : _9562;
    assign _597 = _9564;
    always @(posedge _791) begin
        if (_789)
            _3687 <= _3118;
        else
            _3687 <= _597;
    end
    assign _9571 = _8620 == _1475;
    assign _9568 = ~ _3920;
    assign _9569 = _3135 & _9568;
    assign _9572 = _9569 & _9571;
    assign _9573 = _9572 ? _5304 : _3684;
    assign _9566 = _5296 == _1475;
    assign _9567 = _5293 & _9566;
    assign _9575 = _9567 ? _1475 : _9573;
    assign _9577 = _805 ? _3118 : _9575;
    assign _598 = _9577;
    always @(posedge _791) begin
        if (_789)
            _3684 <= _3118;
        else
            _3684 <= _598;
    end
    assign _9584 = _8620 == _1484;
    assign _9581 = ~ _3920;
    assign _9582 = _3135 & _9581;
    assign _9585 = _9582 & _9584;
    assign _9586 = _9585 ? _5304 : _3681;
    assign _9579 = _5296 == _1484;
    assign _9580 = _5293 & _9579;
    assign _9588 = _9580 ? _1484 : _9586;
    assign _9590 = _805 ? _3118 : _9588;
    assign _599 = _9590;
    always @(posedge _791) begin
        if (_789)
            _3681 <= _3118;
        else
            _3681 <= _599;
    end
    assign _9597 = _8620 == _1493;
    assign _9594 = ~ _3920;
    assign _9595 = _3135 & _9594;
    assign _9598 = _9595 & _9597;
    assign _9599 = _9598 ? _5304 : _3678;
    assign _9592 = _5296 == _1493;
    assign _9593 = _5293 & _9592;
    assign _9601 = _9593 ? _1493 : _9599;
    assign _9603 = _805 ? _3118 : _9601;
    assign _600 = _9603;
    always @(posedge _791) begin
        if (_789)
            _3678 <= _3118;
        else
            _3678 <= _600;
    end
    assign _9610 = _8620 == _1502;
    assign _9607 = ~ _3920;
    assign _9608 = _3135 & _9607;
    assign _9611 = _9608 & _9610;
    assign _9612 = _9611 ? _5304 : _3675;
    assign _9605 = _5296 == _1502;
    assign _9606 = _5293 & _9605;
    assign _9614 = _9606 ? _1502 : _9612;
    assign _9616 = _805 ? _3118 : _9614;
    assign _601 = _9616;
    always @(posedge _791) begin
        if (_789)
            _3675 <= _3118;
        else
            _3675 <= _601;
    end
    assign _9623 = _8620 == _1511;
    assign _9620 = ~ _3920;
    assign _9621 = _3135 & _9620;
    assign _9624 = _9621 & _9623;
    assign _9625 = _9624 ? _5304 : _3672;
    assign _9618 = _5296 == _1511;
    assign _9619 = _5293 & _9618;
    assign _9627 = _9619 ? _1511 : _9625;
    assign _9629 = _805 ? _3118 : _9627;
    assign _602 = _9629;
    always @(posedge _791) begin
        if (_789)
            _3672 <= _3118;
        else
            _3672 <= _602;
    end
    assign _9636 = _8620 == _1520;
    assign _9633 = ~ _3920;
    assign _9634 = _3135 & _9633;
    assign _9637 = _9634 & _9636;
    assign _9638 = _9637 ? _5304 : _3669;
    assign _9631 = _5296 == _1520;
    assign _9632 = _5293 & _9631;
    assign _9640 = _9632 ? _1520 : _9638;
    assign _9642 = _805 ? _3118 : _9640;
    assign _603 = _9642;
    always @(posedge _791) begin
        if (_789)
            _3669 <= _3118;
        else
            _3669 <= _603;
    end
    assign _9649 = _8620 == _1529;
    assign _9646 = ~ _3920;
    assign _9647 = _3135 & _9646;
    assign _9650 = _9647 & _9649;
    assign _9651 = _9650 ? _5304 : _3666;
    assign _9644 = _5296 == _1529;
    assign _9645 = _5293 & _9644;
    assign _9653 = _9645 ? _1529 : _9651;
    assign _9655 = _805 ? _3118 : _9653;
    assign _604 = _9655;
    always @(posedge _791) begin
        if (_789)
            _3666 <= _3118;
        else
            _3666 <= _604;
    end
    assign _9662 = _8620 == _1538;
    assign _9659 = ~ _3920;
    assign _9660 = _3135 & _9659;
    assign _9663 = _9660 & _9662;
    assign _9664 = _9663 ? _5304 : _3663;
    assign _9657 = _5296 == _1538;
    assign _9658 = _5293 & _9657;
    assign _9666 = _9658 ? _1538 : _9664;
    assign _9668 = _805 ? _3118 : _9666;
    assign _605 = _9668;
    always @(posedge _791) begin
        if (_789)
            _3663 <= _3118;
        else
            _3663 <= _605;
    end
    assign _9675 = _8620 == _1547;
    assign _9672 = ~ _3920;
    assign _9673 = _3135 & _9672;
    assign _9676 = _9673 & _9675;
    assign _9677 = _9676 ? _5304 : _3660;
    assign _9670 = _5296 == _1547;
    assign _9671 = _5293 & _9670;
    assign _9679 = _9671 ? _1547 : _9677;
    assign _9681 = _805 ? _3118 : _9679;
    assign _606 = _9681;
    always @(posedge _791) begin
        if (_789)
            _3660 <= _3118;
        else
            _3660 <= _606;
    end
    assign _9688 = _8620 == _1556;
    assign _9685 = ~ _3920;
    assign _9686 = _3135 & _9685;
    assign _9689 = _9686 & _9688;
    assign _9690 = _9689 ? _5304 : _3657;
    assign _9683 = _5296 == _1556;
    assign _9684 = _5293 & _9683;
    assign _9692 = _9684 ? _1556 : _9690;
    assign _9694 = _805 ? _3118 : _9692;
    assign _607 = _9694;
    always @(posedge _791) begin
        if (_789)
            _3657 <= _3118;
        else
            _3657 <= _607;
    end
    assign _9701 = _8620 == _1565;
    assign _9698 = ~ _3920;
    assign _9699 = _3135 & _9698;
    assign _9702 = _9699 & _9701;
    assign _9703 = _9702 ? _5304 : _3654;
    assign _9696 = _5296 == _1565;
    assign _9697 = _5293 & _9696;
    assign _9705 = _9697 ? _1565 : _9703;
    assign _9707 = _805 ? _3118 : _9705;
    assign _608 = _9707;
    always @(posedge _791) begin
        if (_789)
            _3654 <= _3118;
        else
            _3654 <= _608;
    end
    assign _9714 = _8620 == _1574;
    assign _9711 = ~ _3920;
    assign _9712 = _3135 & _9711;
    assign _9715 = _9712 & _9714;
    assign _9716 = _9715 ? _5304 : _3651;
    assign _9709 = _5296 == _1574;
    assign _9710 = _5293 & _9709;
    assign _9718 = _9710 ? _1574 : _9716;
    assign _9720 = _805 ? _3118 : _9718;
    assign _609 = _9720;
    always @(posedge _791) begin
        if (_789)
            _3651 <= _3118;
        else
            _3651 <= _609;
    end
    assign _9727 = _8620 == _1583;
    assign _9724 = ~ _3920;
    assign _9725 = _3135 & _9724;
    assign _9728 = _9725 & _9727;
    assign _9729 = _9728 ? _5304 : _3648;
    assign _9722 = _5296 == _1583;
    assign _9723 = _5293 & _9722;
    assign _9731 = _9723 ? _1583 : _9729;
    assign _9733 = _805 ? _3118 : _9731;
    assign _610 = _9733;
    always @(posedge _791) begin
        if (_789)
            _3648 <= _3118;
        else
            _3648 <= _610;
    end
    assign _9740 = _8620 == _1592;
    assign _9737 = ~ _3920;
    assign _9738 = _3135 & _9737;
    assign _9741 = _9738 & _9740;
    assign _9742 = _9741 ? _5304 : _3645;
    assign _9735 = _5296 == _1592;
    assign _9736 = _5293 & _9735;
    assign _9744 = _9736 ? _1592 : _9742;
    assign _9746 = _805 ? _3118 : _9744;
    assign _611 = _9746;
    always @(posedge _791) begin
        if (_789)
            _3645 <= _3118;
        else
            _3645 <= _611;
    end
    assign _9753 = _8620 == _1601;
    assign _9750 = ~ _3920;
    assign _9751 = _3135 & _9750;
    assign _9754 = _9751 & _9753;
    assign _9755 = _9754 ? _5304 : _3642;
    assign _9748 = _5296 == _1601;
    assign _9749 = _5293 & _9748;
    assign _9757 = _9749 ? _1601 : _9755;
    assign _9759 = _805 ? _3118 : _9757;
    assign _612 = _9759;
    always @(posedge _791) begin
        if (_789)
            _3642 <= _3118;
        else
            _3642 <= _612;
    end
    assign _9766 = _8620 == _1610;
    assign _9763 = ~ _3920;
    assign _9764 = _3135 & _9763;
    assign _9767 = _9764 & _9766;
    assign _9768 = _9767 ? _5304 : _3639;
    assign _9761 = _5296 == _1610;
    assign _9762 = _5293 & _9761;
    assign _9770 = _9762 ? _1610 : _9768;
    assign _9772 = _805 ? _3118 : _9770;
    assign _613 = _9772;
    always @(posedge _791) begin
        if (_789)
            _3639 <= _3118;
        else
            _3639 <= _613;
    end
    assign _9779 = _8620 == _1619;
    assign _9776 = ~ _3920;
    assign _9777 = _3135 & _9776;
    assign _9780 = _9777 & _9779;
    assign _9781 = _9780 ? _5304 : _3636;
    assign _9774 = _5296 == _1619;
    assign _9775 = _5293 & _9774;
    assign _9783 = _9775 ? _1619 : _9781;
    assign _9785 = _805 ? _3118 : _9783;
    assign _614 = _9785;
    always @(posedge _791) begin
        if (_789)
            _3636 <= _3118;
        else
            _3636 <= _614;
    end
    assign _9792 = _8620 == _1628;
    assign _9789 = ~ _3920;
    assign _9790 = _3135 & _9789;
    assign _9793 = _9790 & _9792;
    assign _9794 = _9793 ? _5304 : _3633;
    assign _9787 = _5296 == _1628;
    assign _9788 = _5293 & _9787;
    assign _9796 = _9788 ? _1628 : _9794;
    assign _9798 = _805 ? _3118 : _9796;
    assign _615 = _9798;
    always @(posedge _791) begin
        if (_789)
            _3633 <= _3118;
        else
            _3633 <= _615;
    end
    assign _9805 = _8620 == _1637;
    assign _9802 = ~ _3920;
    assign _9803 = _3135 & _9802;
    assign _9806 = _9803 & _9805;
    assign _9807 = _9806 ? _5304 : _3630;
    assign _9800 = _5296 == _1637;
    assign _9801 = _5293 & _9800;
    assign _9809 = _9801 ? _1637 : _9807;
    assign _9811 = _805 ? _3118 : _9809;
    assign _616 = _9811;
    always @(posedge _791) begin
        if (_789)
            _3630 <= _3118;
        else
            _3630 <= _616;
    end
    assign _9818 = _8620 == _1646;
    assign _9815 = ~ _3920;
    assign _9816 = _3135 & _9815;
    assign _9819 = _9816 & _9818;
    assign _9820 = _9819 ? _5304 : _3627;
    assign _9813 = _5296 == _1646;
    assign _9814 = _5293 & _9813;
    assign _9822 = _9814 ? _1646 : _9820;
    assign _9824 = _805 ? _3118 : _9822;
    assign _617 = _9824;
    always @(posedge _791) begin
        if (_789)
            _3627 <= _3118;
        else
            _3627 <= _617;
    end
    assign _9831 = _8620 == _1655;
    assign _9828 = ~ _3920;
    assign _9829 = _3135 & _9828;
    assign _9832 = _9829 & _9831;
    assign _9833 = _9832 ? _5304 : _3624;
    assign _9826 = _5296 == _1655;
    assign _9827 = _5293 & _9826;
    assign _9835 = _9827 ? _1655 : _9833;
    assign _9837 = _805 ? _3118 : _9835;
    assign _618 = _9837;
    always @(posedge _791) begin
        if (_789)
            _3624 <= _3118;
        else
            _3624 <= _618;
    end
    assign _9844 = _8620 == _1664;
    assign _9841 = ~ _3920;
    assign _9842 = _3135 & _9841;
    assign _9845 = _9842 & _9844;
    assign _9846 = _9845 ? _5304 : _3621;
    assign _9839 = _5296 == _1664;
    assign _9840 = _5293 & _9839;
    assign _9848 = _9840 ? _1664 : _9846;
    assign _9850 = _805 ? _3118 : _9848;
    assign _619 = _9850;
    always @(posedge _791) begin
        if (_789)
            _3621 <= _3118;
        else
            _3621 <= _619;
    end
    assign _9857 = _8620 == _1673;
    assign _9854 = ~ _3920;
    assign _9855 = _3135 & _9854;
    assign _9858 = _9855 & _9857;
    assign _9859 = _9858 ? _5304 : _3618;
    assign _9852 = _5296 == _1673;
    assign _9853 = _5293 & _9852;
    assign _9861 = _9853 ? _1673 : _9859;
    assign _9863 = _805 ? _3118 : _9861;
    assign _620 = _9863;
    always @(posedge _791) begin
        if (_789)
            _3618 <= _3118;
        else
            _3618 <= _620;
    end
    assign _9870 = _8620 == _1682;
    assign _9867 = ~ _3920;
    assign _9868 = _3135 & _9867;
    assign _9871 = _9868 & _9870;
    assign _9872 = _9871 ? _5304 : _3615;
    assign _9865 = _5296 == _1682;
    assign _9866 = _5293 & _9865;
    assign _9874 = _9866 ? _1682 : _9872;
    assign _9876 = _805 ? _3118 : _9874;
    assign _621 = _9876;
    always @(posedge _791) begin
        if (_789)
            _3615 <= _3118;
        else
            _3615 <= _621;
    end
    assign _9883 = _8620 == _1691;
    assign _9880 = ~ _3920;
    assign _9881 = _3135 & _9880;
    assign _9884 = _9881 & _9883;
    assign _9885 = _9884 ? _5304 : _3612;
    assign _9878 = _5296 == _1691;
    assign _9879 = _5293 & _9878;
    assign _9887 = _9879 ? _1691 : _9885;
    assign _9889 = _805 ? _3118 : _9887;
    assign _622 = _9889;
    always @(posedge _791) begin
        if (_789)
            _3612 <= _3118;
        else
            _3612 <= _622;
    end
    assign _9896 = _8620 == _1700;
    assign _9893 = ~ _3920;
    assign _9894 = _3135 & _9893;
    assign _9897 = _9894 & _9896;
    assign _9898 = _9897 ? _5304 : _3609;
    assign _9891 = _5296 == _1700;
    assign _9892 = _5293 & _9891;
    assign _9900 = _9892 ? _1700 : _9898;
    assign _9902 = _805 ? _3118 : _9900;
    assign _623 = _9902;
    always @(posedge _791) begin
        if (_789)
            _3609 <= _3118;
        else
            _3609 <= _623;
    end
    assign _9909 = _8620 == _1709;
    assign _9906 = ~ _3920;
    assign _9907 = _3135 & _9906;
    assign _9910 = _9907 & _9909;
    assign _9911 = _9910 ? _5304 : _3606;
    assign _9904 = _5296 == _1709;
    assign _9905 = _5293 & _9904;
    assign _9913 = _9905 ? _1709 : _9911;
    assign _9915 = _805 ? _3118 : _9913;
    assign _624 = _9915;
    always @(posedge _791) begin
        if (_789)
            _3606 <= _3118;
        else
            _3606 <= _624;
    end
    assign _9922 = _8620 == _1718;
    assign _9919 = ~ _3920;
    assign _9920 = _3135 & _9919;
    assign _9923 = _9920 & _9922;
    assign _9924 = _9923 ? _5304 : _3603;
    assign _9917 = _5296 == _1718;
    assign _9918 = _5293 & _9917;
    assign _9926 = _9918 ? _1718 : _9924;
    assign _9928 = _805 ? _3118 : _9926;
    assign _625 = _9928;
    always @(posedge _791) begin
        if (_789)
            _3603 <= _3118;
        else
            _3603 <= _625;
    end
    assign _9935 = _8620 == _1727;
    assign _9932 = ~ _3920;
    assign _9933 = _3135 & _9932;
    assign _9936 = _9933 & _9935;
    assign _9937 = _9936 ? _5304 : _3600;
    assign _9930 = _5296 == _1727;
    assign _9931 = _5293 & _9930;
    assign _9939 = _9931 ? _1727 : _9937;
    assign _9941 = _805 ? _3118 : _9939;
    assign _626 = _9941;
    always @(posedge _791) begin
        if (_789)
            _3600 <= _3118;
        else
            _3600 <= _626;
    end
    assign _9948 = _8620 == _1736;
    assign _9945 = ~ _3920;
    assign _9946 = _3135 & _9945;
    assign _9949 = _9946 & _9948;
    assign _9950 = _9949 ? _5304 : _3597;
    assign _9943 = _5296 == _1736;
    assign _9944 = _5293 & _9943;
    assign _9952 = _9944 ? _1736 : _9950;
    assign _9954 = _805 ? _3118 : _9952;
    assign _627 = _9954;
    always @(posedge _791) begin
        if (_789)
            _3597 <= _3118;
        else
            _3597 <= _627;
    end
    assign _9961 = _8620 == _1745;
    assign _9958 = ~ _3920;
    assign _9959 = _3135 & _9958;
    assign _9962 = _9959 & _9961;
    assign _9963 = _9962 ? _5304 : _3594;
    assign _9956 = _5296 == _1745;
    assign _9957 = _5293 & _9956;
    assign _9965 = _9957 ? _1745 : _9963;
    assign _9967 = _805 ? _3118 : _9965;
    assign _628 = _9967;
    always @(posedge _791) begin
        if (_789)
            _3594 <= _3118;
        else
            _3594 <= _628;
    end
    assign _9974 = _8620 == _1754;
    assign _9971 = ~ _3920;
    assign _9972 = _3135 & _9971;
    assign _9975 = _9972 & _9974;
    assign _9976 = _9975 ? _5304 : _3591;
    assign _9969 = _5296 == _1754;
    assign _9970 = _5293 & _9969;
    assign _9978 = _9970 ? _1754 : _9976;
    assign _9980 = _805 ? _3118 : _9978;
    assign _629 = _9980;
    always @(posedge _791) begin
        if (_789)
            _3591 <= _3118;
        else
            _3591 <= _629;
    end
    assign _9987 = _8620 == _1763;
    assign _9984 = ~ _3920;
    assign _9985 = _3135 & _9984;
    assign _9988 = _9985 & _9987;
    assign _9989 = _9988 ? _5304 : _3588;
    assign _9982 = _5296 == _1763;
    assign _9983 = _5293 & _9982;
    assign _9991 = _9983 ? _1763 : _9989;
    assign _9993 = _805 ? _3118 : _9991;
    assign _630 = _9993;
    always @(posedge _791) begin
        if (_789)
            _3588 <= _3118;
        else
            _3588 <= _630;
    end
    assign _10000 = _8620 == _1772;
    assign _9997 = ~ _3920;
    assign _9998 = _3135 & _9997;
    assign _10001 = _9998 & _10000;
    assign _10002 = _10001 ? _5304 : _3585;
    assign _9995 = _5296 == _1772;
    assign _9996 = _5293 & _9995;
    assign _10004 = _9996 ? _1772 : _10002;
    assign _10006 = _805 ? _3118 : _10004;
    assign _631 = _10006;
    always @(posedge _791) begin
        if (_789)
            _3585 <= _3118;
        else
            _3585 <= _631;
    end
    assign _10013 = _8620 == _1781;
    assign _10010 = ~ _3920;
    assign _10011 = _3135 & _10010;
    assign _10014 = _10011 & _10013;
    assign _10015 = _10014 ? _5304 : _3582;
    assign _10008 = _5296 == _1781;
    assign _10009 = _5293 & _10008;
    assign _10017 = _10009 ? _1781 : _10015;
    assign _10019 = _805 ? _3118 : _10017;
    assign _632 = _10019;
    always @(posedge _791) begin
        if (_789)
            _3582 <= _3118;
        else
            _3582 <= _632;
    end
    assign _10026 = _8620 == _1790;
    assign _10023 = ~ _3920;
    assign _10024 = _3135 & _10023;
    assign _10027 = _10024 & _10026;
    assign _10028 = _10027 ? _5304 : _3579;
    assign _10021 = _5296 == _1790;
    assign _10022 = _5293 & _10021;
    assign _10030 = _10022 ? _1790 : _10028;
    assign _10032 = _805 ? _3118 : _10030;
    assign _633 = _10032;
    always @(posedge _791) begin
        if (_789)
            _3579 <= _3118;
        else
            _3579 <= _633;
    end
    assign _10039 = _8620 == _1799;
    assign _10036 = ~ _3920;
    assign _10037 = _3135 & _10036;
    assign _10040 = _10037 & _10039;
    assign _10041 = _10040 ? _5304 : _3576;
    assign _10034 = _5296 == _1799;
    assign _10035 = _5293 & _10034;
    assign _10043 = _10035 ? _1799 : _10041;
    assign _10045 = _805 ? _3118 : _10043;
    assign _634 = _10045;
    always @(posedge _791) begin
        if (_789)
            _3576 <= _3118;
        else
            _3576 <= _634;
    end
    assign _10052 = _8620 == _1808;
    assign _10049 = ~ _3920;
    assign _10050 = _3135 & _10049;
    assign _10053 = _10050 & _10052;
    assign _10054 = _10053 ? _5304 : _3573;
    assign _10047 = _5296 == _1808;
    assign _10048 = _5293 & _10047;
    assign _10056 = _10048 ? _1808 : _10054;
    assign _10058 = _805 ? _3118 : _10056;
    assign _635 = _10058;
    always @(posedge _791) begin
        if (_789)
            _3573 <= _3118;
        else
            _3573 <= _635;
    end
    assign _10065 = _8620 == _1817;
    assign _10062 = ~ _3920;
    assign _10063 = _3135 & _10062;
    assign _10066 = _10063 & _10065;
    assign _10067 = _10066 ? _5304 : _3570;
    assign _10060 = _5296 == _1817;
    assign _10061 = _5293 & _10060;
    assign _10069 = _10061 ? _1817 : _10067;
    assign _10071 = _805 ? _3118 : _10069;
    assign _636 = _10071;
    always @(posedge _791) begin
        if (_789)
            _3570 <= _3118;
        else
            _3570 <= _636;
    end
    assign _10078 = _8620 == _1826;
    assign _10075 = ~ _3920;
    assign _10076 = _3135 & _10075;
    assign _10079 = _10076 & _10078;
    assign _10080 = _10079 ? _5304 : _3567;
    assign _10073 = _5296 == _1826;
    assign _10074 = _5293 & _10073;
    assign _10082 = _10074 ? _1826 : _10080;
    assign _10084 = _805 ? _3118 : _10082;
    assign _637 = _10084;
    always @(posedge _791) begin
        if (_789)
            _3567 <= _3118;
        else
            _3567 <= _637;
    end
    assign _10091 = _8620 == _1835;
    assign _10088 = ~ _3920;
    assign _10089 = _3135 & _10088;
    assign _10092 = _10089 & _10091;
    assign _10093 = _10092 ? _5304 : _3564;
    assign _10086 = _5296 == _1835;
    assign _10087 = _5293 & _10086;
    assign _10095 = _10087 ? _1835 : _10093;
    assign _10097 = _805 ? _3118 : _10095;
    assign _638 = _10097;
    always @(posedge _791) begin
        if (_789)
            _3564 <= _3118;
        else
            _3564 <= _638;
    end
    assign _10104 = _8620 == _1844;
    assign _10101 = ~ _3920;
    assign _10102 = _3135 & _10101;
    assign _10105 = _10102 & _10104;
    assign _10106 = _10105 ? _5304 : _3561;
    assign _10099 = _5296 == _1844;
    assign _10100 = _5293 & _10099;
    assign _10108 = _10100 ? _1844 : _10106;
    assign _10110 = _805 ? _3118 : _10108;
    assign _639 = _10110;
    always @(posedge _791) begin
        if (_789)
            _3561 <= _3118;
        else
            _3561 <= _639;
    end
    assign _10117 = _8620 == _1853;
    assign _10114 = ~ _3920;
    assign _10115 = _3135 & _10114;
    assign _10118 = _10115 & _10117;
    assign _10119 = _10118 ? _5304 : _3558;
    assign _10112 = _5296 == _1853;
    assign _10113 = _5293 & _10112;
    assign _10121 = _10113 ? _1853 : _10119;
    assign _10123 = _805 ? _3118 : _10121;
    assign _640 = _10123;
    always @(posedge _791) begin
        if (_789)
            _3558 <= _3118;
        else
            _3558 <= _640;
    end
    assign _10130 = _8620 == _1862;
    assign _10127 = ~ _3920;
    assign _10128 = _3135 & _10127;
    assign _10131 = _10128 & _10130;
    assign _10132 = _10131 ? _5304 : _3555;
    assign _10125 = _5296 == _1862;
    assign _10126 = _5293 & _10125;
    assign _10134 = _10126 ? _1862 : _10132;
    assign _10136 = _805 ? _3118 : _10134;
    assign _641 = _10136;
    always @(posedge _791) begin
        if (_789)
            _3555 <= _3118;
        else
            _3555 <= _641;
    end
    assign _10143 = _8620 == _1871;
    assign _10140 = ~ _3920;
    assign _10141 = _3135 & _10140;
    assign _10144 = _10141 & _10143;
    assign _10145 = _10144 ? _5304 : _3552;
    assign _10138 = _5296 == _1871;
    assign _10139 = _5293 & _10138;
    assign _10147 = _10139 ? _1871 : _10145;
    assign _10149 = _805 ? _3118 : _10147;
    assign _642 = _10149;
    always @(posedge _791) begin
        if (_789)
            _3552 <= _3118;
        else
            _3552 <= _642;
    end
    assign _10156 = _8620 == _1880;
    assign _10153 = ~ _3920;
    assign _10154 = _3135 & _10153;
    assign _10157 = _10154 & _10156;
    assign _10158 = _10157 ? _5304 : _3549;
    assign _10151 = _5296 == _1880;
    assign _10152 = _5293 & _10151;
    assign _10160 = _10152 ? _1880 : _10158;
    assign _10162 = _805 ? _3118 : _10160;
    assign _643 = _10162;
    always @(posedge _791) begin
        if (_789)
            _3549 <= _3118;
        else
            _3549 <= _643;
    end
    assign _10169 = _8620 == _1889;
    assign _10166 = ~ _3920;
    assign _10167 = _3135 & _10166;
    assign _10170 = _10167 & _10169;
    assign _10171 = _10170 ? _5304 : _3546;
    assign _10164 = _5296 == _1889;
    assign _10165 = _5293 & _10164;
    assign _10173 = _10165 ? _1889 : _10171;
    assign _10175 = _805 ? _3118 : _10173;
    assign _644 = _10175;
    always @(posedge _791) begin
        if (_789)
            _3546 <= _3118;
        else
            _3546 <= _644;
    end
    assign _10182 = _8620 == _1898;
    assign _10179 = ~ _3920;
    assign _10180 = _3135 & _10179;
    assign _10183 = _10180 & _10182;
    assign _10184 = _10183 ? _5304 : _3543;
    assign _10177 = _5296 == _1898;
    assign _10178 = _5293 & _10177;
    assign _10186 = _10178 ? _1898 : _10184;
    assign _10188 = _805 ? _3118 : _10186;
    assign _645 = _10188;
    always @(posedge _791) begin
        if (_789)
            _3543 <= _3118;
        else
            _3543 <= _645;
    end
    assign _10195 = _8620 == _1907;
    assign _10192 = ~ _3920;
    assign _10193 = _3135 & _10192;
    assign _10196 = _10193 & _10195;
    assign _10197 = _10196 ? _5304 : _3540;
    assign _10190 = _5296 == _1907;
    assign _10191 = _5293 & _10190;
    assign _10199 = _10191 ? _1907 : _10197;
    assign _10201 = _805 ? _3118 : _10199;
    assign _646 = _10201;
    always @(posedge _791) begin
        if (_789)
            _3540 <= _3118;
        else
            _3540 <= _646;
    end
    assign _10208 = _8620 == _1916;
    assign _10205 = ~ _3920;
    assign _10206 = _3135 & _10205;
    assign _10209 = _10206 & _10208;
    assign _10210 = _10209 ? _5304 : _3537;
    assign _10203 = _5296 == _1916;
    assign _10204 = _5293 & _10203;
    assign _10212 = _10204 ? _1916 : _10210;
    assign _10214 = _805 ? _3118 : _10212;
    assign _647 = _10214;
    always @(posedge _791) begin
        if (_789)
            _3537 <= _3118;
        else
            _3537 <= _647;
    end
    assign _10221 = _8620 == _1925;
    assign _10218 = ~ _3920;
    assign _10219 = _3135 & _10218;
    assign _10222 = _10219 & _10221;
    assign _10223 = _10222 ? _5304 : _3534;
    assign _10216 = _5296 == _1925;
    assign _10217 = _5293 & _10216;
    assign _10225 = _10217 ? _1925 : _10223;
    assign _10227 = _805 ? _3118 : _10225;
    assign _648 = _10227;
    always @(posedge _791) begin
        if (_789)
            _3534 <= _3118;
        else
            _3534 <= _648;
    end
    assign _10234 = _8620 == _1934;
    assign _10231 = ~ _3920;
    assign _10232 = _3135 & _10231;
    assign _10235 = _10232 & _10234;
    assign _10236 = _10235 ? _5304 : _3531;
    assign _10229 = _5296 == _1934;
    assign _10230 = _5293 & _10229;
    assign _10238 = _10230 ? _1934 : _10236;
    assign _10240 = _805 ? _3118 : _10238;
    assign _649 = _10240;
    always @(posedge _791) begin
        if (_789)
            _3531 <= _3118;
        else
            _3531 <= _649;
    end
    assign _10247 = _8620 == _1943;
    assign _10244 = ~ _3920;
    assign _10245 = _3135 & _10244;
    assign _10248 = _10245 & _10247;
    assign _10249 = _10248 ? _5304 : _3528;
    assign _10242 = _5296 == _1943;
    assign _10243 = _5293 & _10242;
    assign _10251 = _10243 ? _1943 : _10249;
    assign _10253 = _805 ? _3118 : _10251;
    assign _650 = _10253;
    always @(posedge _791) begin
        if (_789)
            _3528 <= _3118;
        else
            _3528 <= _650;
    end
    assign _10260 = _8620 == _1952;
    assign _10257 = ~ _3920;
    assign _10258 = _3135 & _10257;
    assign _10261 = _10258 & _10260;
    assign _10262 = _10261 ? _5304 : _3525;
    assign _10255 = _5296 == _1952;
    assign _10256 = _5293 & _10255;
    assign _10264 = _10256 ? _1952 : _10262;
    assign _10266 = _805 ? _3118 : _10264;
    assign _651 = _10266;
    always @(posedge _791) begin
        if (_789)
            _3525 <= _3118;
        else
            _3525 <= _651;
    end
    assign _10273 = _8620 == _1961;
    assign _10270 = ~ _3920;
    assign _10271 = _3135 & _10270;
    assign _10274 = _10271 & _10273;
    assign _10275 = _10274 ? _5304 : _3522;
    assign _10268 = _5296 == _1961;
    assign _10269 = _5293 & _10268;
    assign _10277 = _10269 ? _1961 : _10275;
    assign _10279 = _805 ? _3118 : _10277;
    assign _652 = _10279;
    always @(posedge _791) begin
        if (_789)
            _3522 <= _3118;
        else
            _3522 <= _652;
    end
    assign _10286 = _8620 == _1970;
    assign _10283 = ~ _3920;
    assign _10284 = _3135 & _10283;
    assign _10287 = _10284 & _10286;
    assign _10288 = _10287 ? _5304 : _3519;
    assign _10281 = _5296 == _1970;
    assign _10282 = _5293 & _10281;
    assign _10290 = _10282 ? _1970 : _10288;
    assign _10292 = _805 ? _3118 : _10290;
    assign _653 = _10292;
    always @(posedge _791) begin
        if (_789)
            _3519 <= _3118;
        else
            _3519 <= _653;
    end
    assign _10299 = _8620 == _1979;
    assign _10296 = ~ _3920;
    assign _10297 = _3135 & _10296;
    assign _10300 = _10297 & _10299;
    assign _10301 = _10300 ? _5304 : _3516;
    assign _10294 = _5296 == _1979;
    assign _10295 = _5293 & _10294;
    assign _10303 = _10295 ? _1979 : _10301;
    assign _10305 = _805 ? _3118 : _10303;
    assign _654 = _10305;
    always @(posedge _791) begin
        if (_789)
            _3516 <= _3118;
        else
            _3516 <= _654;
    end
    assign _10312 = _8620 == _1988;
    assign _10309 = ~ _3920;
    assign _10310 = _3135 & _10309;
    assign _10313 = _10310 & _10312;
    assign _10314 = _10313 ? _5304 : _3513;
    assign _10307 = _5296 == _1988;
    assign _10308 = _5293 & _10307;
    assign _10316 = _10308 ? _1988 : _10314;
    assign _10318 = _805 ? _3118 : _10316;
    assign _655 = _10318;
    always @(posedge _791) begin
        if (_789)
            _3513 <= _3118;
        else
            _3513 <= _655;
    end
    assign _10325 = _8620 == _1997;
    assign _10322 = ~ _3920;
    assign _10323 = _3135 & _10322;
    assign _10326 = _10323 & _10325;
    assign _10327 = _10326 ? _5304 : _3510;
    assign _10320 = _5296 == _1997;
    assign _10321 = _5293 & _10320;
    assign _10329 = _10321 ? _1997 : _10327;
    assign _10331 = _805 ? _3118 : _10329;
    assign _656 = _10331;
    always @(posedge _791) begin
        if (_789)
            _3510 <= _3118;
        else
            _3510 <= _656;
    end
    assign _10338 = _8620 == _2006;
    assign _10335 = ~ _3920;
    assign _10336 = _3135 & _10335;
    assign _10339 = _10336 & _10338;
    assign _10340 = _10339 ? _5304 : _3507;
    assign _10333 = _5296 == _2006;
    assign _10334 = _5293 & _10333;
    assign _10342 = _10334 ? _2006 : _10340;
    assign _10344 = _805 ? _3118 : _10342;
    assign _657 = _10344;
    always @(posedge _791) begin
        if (_789)
            _3507 <= _3118;
        else
            _3507 <= _657;
    end
    assign _10351 = _8620 == _2015;
    assign _10348 = ~ _3920;
    assign _10349 = _3135 & _10348;
    assign _10352 = _10349 & _10351;
    assign _10353 = _10352 ? _5304 : _3504;
    assign _10346 = _5296 == _2015;
    assign _10347 = _5293 & _10346;
    assign _10355 = _10347 ? _2015 : _10353;
    assign _10357 = _805 ? _3118 : _10355;
    assign _658 = _10357;
    always @(posedge _791) begin
        if (_789)
            _3504 <= _3118;
        else
            _3504 <= _658;
    end
    assign _10364 = _8620 == _2024;
    assign _10361 = ~ _3920;
    assign _10362 = _3135 & _10361;
    assign _10365 = _10362 & _10364;
    assign _10366 = _10365 ? _5304 : _3501;
    assign _10359 = _5296 == _2024;
    assign _10360 = _5293 & _10359;
    assign _10368 = _10360 ? _2024 : _10366;
    assign _10370 = _805 ? _3118 : _10368;
    assign _659 = _10370;
    always @(posedge _791) begin
        if (_789)
            _3501 <= _3118;
        else
            _3501 <= _659;
    end
    assign _10377 = _8620 == _2033;
    assign _10374 = ~ _3920;
    assign _10375 = _3135 & _10374;
    assign _10378 = _10375 & _10377;
    assign _10379 = _10378 ? _5304 : _3498;
    assign _10372 = _5296 == _2033;
    assign _10373 = _5293 & _10372;
    assign _10381 = _10373 ? _2033 : _10379;
    assign _10383 = _805 ? _3118 : _10381;
    assign _660 = _10383;
    always @(posedge _791) begin
        if (_789)
            _3498 <= _3118;
        else
            _3498 <= _660;
    end
    assign _10390 = _8620 == _2042;
    assign _10387 = ~ _3920;
    assign _10388 = _3135 & _10387;
    assign _10391 = _10388 & _10390;
    assign _10392 = _10391 ? _5304 : _3495;
    assign _10385 = _5296 == _2042;
    assign _10386 = _5293 & _10385;
    assign _10394 = _10386 ? _2042 : _10392;
    assign _10396 = _805 ? _3118 : _10394;
    assign _661 = _10396;
    always @(posedge _791) begin
        if (_789)
            _3495 <= _3118;
        else
            _3495 <= _661;
    end
    assign _10403 = _8620 == _2051;
    assign _10400 = ~ _3920;
    assign _10401 = _3135 & _10400;
    assign _10404 = _10401 & _10403;
    assign _10405 = _10404 ? _5304 : _3492;
    assign _10398 = _5296 == _2051;
    assign _10399 = _5293 & _10398;
    assign _10407 = _10399 ? _2051 : _10405;
    assign _10409 = _805 ? _3118 : _10407;
    assign _662 = _10409;
    always @(posedge _791) begin
        if (_789)
            _3492 <= _3118;
        else
            _3492 <= _662;
    end
    assign _10416 = _8620 == _2060;
    assign _10413 = ~ _3920;
    assign _10414 = _3135 & _10413;
    assign _10417 = _10414 & _10416;
    assign _10418 = _10417 ? _5304 : _3489;
    assign _10411 = _5296 == _2060;
    assign _10412 = _5293 & _10411;
    assign _10420 = _10412 ? _2060 : _10418;
    assign _10422 = _805 ? _3118 : _10420;
    assign _663 = _10422;
    always @(posedge _791) begin
        if (_789)
            _3489 <= _3118;
        else
            _3489 <= _663;
    end
    assign _10429 = _8620 == _2069;
    assign _10426 = ~ _3920;
    assign _10427 = _3135 & _10426;
    assign _10430 = _10427 & _10429;
    assign _10431 = _10430 ? _5304 : _3486;
    assign _10424 = _5296 == _2069;
    assign _10425 = _5293 & _10424;
    assign _10433 = _10425 ? _2069 : _10431;
    assign _10435 = _805 ? _3118 : _10433;
    assign _664 = _10435;
    always @(posedge _791) begin
        if (_789)
            _3486 <= _3118;
        else
            _3486 <= _664;
    end
    assign _10442 = _8620 == _2078;
    assign _10439 = ~ _3920;
    assign _10440 = _3135 & _10439;
    assign _10443 = _10440 & _10442;
    assign _10444 = _10443 ? _5304 : _3483;
    assign _10437 = _5296 == _2078;
    assign _10438 = _5293 & _10437;
    assign _10446 = _10438 ? _2078 : _10444;
    assign _10448 = _805 ? _3118 : _10446;
    assign _665 = _10448;
    always @(posedge _791) begin
        if (_789)
            _3483 <= _3118;
        else
            _3483 <= _665;
    end
    assign _10455 = _8620 == _2087;
    assign _10452 = ~ _3920;
    assign _10453 = _3135 & _10452;
    assign _10456 = _10453 & _10455;
    assign _10457 = _10456 ? _5304 : _3480;
    assign _10450 = _5296 == _2087;
    assign _10451 = _5293 & _10450;
    assign _10459 = _10451 ? _2087 : _10457;
    assign _10461 = _805 ? _3118 : _10459;
    assign _666 = _10461;
    always @(posedge _791) begin
        if (_789)
            _3480 <= _3118;
        else
            _3480 <= _666;
    end
    assign _10468 = _8620 == _2096;
    assign _10465 = ~ _3920;
    assign _10466 = _3135 & _10465;
    assign _10469 = _10466 & _10468;
    assign _10470 = _10469 ? _5304 : _3477;
    assign _10463 = _5296 == _2096;
    assign _10464 = _5293 & _10463;
    assign _10472 = _10464 ? _2096 : _10470;
    assign _10474 = _805 ? _3118 : _10472;
    assign _667 = _10474;
    always @(posedge _791) begin
        if (_789)
            _3477 <= _3118;
        else
            _3477 <= _667;
    end
    assign _10481 = _8620 == _2105;
    assign _10478 = ~ _3920;
    assign _10479 = _3135 & _10478;
    assign _10482 = _10479 & _10481;
    assign _10483 = _10482 ? _5304 : _3474;
    assign _10476 = _5296 == _2105;
    assign _10477 = _5293 & _10476;
    assign _10485 = _10477 ? _2105 : _10483;
    assign _10487 = _805 ? _3118 : _10485;
    assign _668 = _10487;
    always @(posedge _791) begin
        if (_789)
            _3474 <= _3118;
        else
            _3474 <= _668;
    end
    assign _10494 = _8620 == _2114;
    assign _10491 = ~ _3920;
    assign _10492 = _3135 & _10491;
    assign _10495 = _10492 & _10494;
    assign _10496 = _10495 ? _5304 : _3471;
    assign _10489 = _5296 == _2114;
    assign _10490 = _5293 & _10489;
    assign _10498 = _10490 ? _2114 : _10496;
    assign _10500 = _805 ? _3118 : _10498;
    assign _669 = _10500;
    always @(posedge _791) begin
        if (_789)
            _3471 <= _3118;
        else
            _3471 <= _669;
    end
    assign _10507 = _8620 == _2123;
    assign _10504 = ~ _3920;
    assign _10505 = _3135 & _10504;
    assign _10508 = _10505 & _10507;
    assign _10509 = _10508 ? _5304 : _3468;
    assign _10502 = _5296 == _2123;
    assign _10503 = _5293 & _10502;
    assign _10511 = _10503 ? _2123 : _10509;
    assign _10513 = _805 ? _3118 : _10511;
    assign _670 = _10513;
    always @(posedge _791) begin
        if (_789)
            _3468 <= _3118;
        else
            _3468 <= _670;
    end
    assign _10520 = _8620 == _2132;
    assign _10517 = ~ _3920;
    assign _10518 = _3135 & _10517;
    assign _10521 = _10518 & _10520;
    assign _10522 = _10521 ? _5304 : _3465;
    assign _10515 = _5296 == _2132;
    assign _10516 = _5293 & _10515;
    assign _10524 = _10516 ? _2132 : _10522;
    assign _10526 = _805 ? _3118 : _10524;
    assign _671 = _10526;
    always @(posedge _791) begin
        if (_789)
            _3465 <= _3118;
        else
            _3465 <= _671;
    end
    assign _10533 = _8620 == _2141;
    assign _10530 = ~ _3920;
    assign _10531 = _3135 & _10530;
    assign _10534 = _10531 & _10533;
    assign _10535 = _10534 ? _5304 : _3462;
    assign _10528 = _5296 == _2141;
    assign _10529 = _5293 & _10528;
    assign _10537 = _10529 ? _2141 : _10535;
    assign _10539 = _805 ? _3118 : _10537;
    assign _672 = _10539;
    always @(posedge _791) begin
        if (_789)
            _3462 <= _3118;
        else
            _3462 <= _672;
    end
    assign _10546 = _8620 == _2150;
    assign _10543 = ~ _3920;
    assign _10544 = _3135 & _10543;
    assign _10547 = _10544 & _10546;
    assign _10548 = _10547 ? _5304 : _3459;
    assign _10541 = _5296 == _2150;
    assign _10542 = _5293 & _10541;
    assign _10550 = _10542 ? _2150 : _10548;
    assign _10552 = _805 ? _3118 : _10550;
    assign _673 = _10552;
    always @(posedge _791) begin
        if (_789)
            _3459 <= _3118;
        else
            _3459 <= _673;
    end
    assign _10559 = _8620 == _2159;
    assign _10556 = ~ _3920;
    assign _10557 = _3135 & _10556;
    assign _10560 = _10557 & _10559;
    assign _10561 = _10560 ? _5304 : _3456;
    assign _10554 = _5296 == _2159;
    assign _10555 = _5293 & _10554;
    assign _10563 = _10555 ? _2159 : _10561;
    assign _10565 = _805 ? _3118 : _10563;
    assign _674 = _10565;
    always @(posedge _791) begin
        if (_789)
            _3456 <= _3118;
        else
            _3456 <= _674;
    end
    assign _10572 = _8620 == _2168;
    assign _10569 = ~ _3920;
    assign _10570 = _3135 & _10569;
    assign _10573 = _10570 & _10572;
    assign _10574 = _10573 ? _5304 : _3453;
    assign _10567 = _5296 == _2168;
    assign _10568 = _5293 & _10567;
    assign _10576 = _10568 ? _2168 : _10574;
    assign _10578 = _805 ? _3118 : _10576;
    assign _675 = _10578;
    always @(posedge _791) begin
        if (_789)
            _3453 <= _3118;
        else
            _3453 <= _675;
    end
    assign _10585 = _8620 == _2177;
    assign _10582 = ~ _3920;
    assign _10583 = _3135 & _10582;
    assign _10586 = _10583 & _10585;
    assign _10587 = _10586 ? _5304 : _3450;
    assign _10580 = _5296 == _2177;
    assign _10581 = _5293 & _10580;
    assign _10589 = _10581 ? _2177 : _10587;
    assign _10591 = _805 ? _3118 : _10589;
    assign _676 = _10591;
    always @(posedge _791) begin
        if (_789)
            _3450 <= _3118;
        else
            _3450 <= _676;
    end
    assign _10598 = _8620 == _2186;
    assign _10595 = ~ _3920;
    assign _10596 = _3135 & _10595;
    assign _10599 = _10596 & _10598;
    assign _10600 = _10599 ? _5304 : _3447;
    assign _10593 = _5296 == _2186;
    assign _10594 = _5293 & _10593;
    assign _10602 = _10594 ? _2186 : _10600;
    assign _10604 = _805 ? _3118 : _10602;
    assign _677 = _10604;
    always @(posedge _791) begin
        if (_789)
            _3447 <= _3118;
        else
            _3447 <= _677;
    end
    assign _10611 = _8620 == _2195;
    assign _10608 = ~ _3920;
    assign _10609 = _3135 & _10608;
    assign _10612 = _10609 & _10611;
    assign _10613 = _10612 ? _5304 : _3444;
    assign _10606 = _5296 == _2195;
    assign _10607 = _5293 & _10606;
    assign _10615 = _10607 ? _2195 : _10613;
    assign _10617 = _805 ? _3118 : _10615;
    assign _678 = _10617;
    always @(posedge _791) begin
        if (_789)
            _3444 <= _3118;
        else
            _3444 <= _678;
    end
    assign _10624 = _8620 == _2204;
    assign _10621 = ~ _3920;
    assign _10622 = _3135 & _10621;
    assign _10625 = _10622 & _10624;
    assign _10626 = _10625 ? _5304 : _3441;
    assign _10619 = _5296 == _2204;
    assign _10620 = _5293 & _10619;
    assign _10628 = _10620 ? _2204 : _10626;
    assign _10630 = _805 ? _3118 : _10628;
    assign _679 = _10630;
    always @(posedge _791) begin
        if (_789)
            _3441 <= _3118;
        else
            _3441 <= _679;
    end
    assign _10637 = _8620 == _2213;
    assign _10634 = ~ _3920;
    assign _10635 = _3135 & _10634;
    assign _10638 = _10635 & _10637;
    assign _10639 = _10638 ? _5304 : _3438;
    assign _10632 = _5296 == _2213;
    assign _10633 = _5293 & _10632;
    assign _10641 = _10633 ? _2213 : _10639;
    assign _10643 = _805 ? _3118 : _10641;
    assign _680 = _10643;
    always @(posedge _791) begin
        if (_789)
            _3438 <= _3118;
        else
            _3438 <= _680;
    end
    assign _10650 = _8620 == _2222;
    assign _10647 = ~ _3920;
    assign _10648 = _3135 & _10647;
    assign _10651 = _10648 & _10650;
    assign _10652 = _10651 ? _5304 : _3435;
    assign _10645 = _5296 == _2222;
    assign _10646 = _5293 & _10645;
    assign _10654 = _10646 ? _2222 : _10652;
    assign _10656 = _805 ? _3118 : _10654;
    assign _681 = _10656;
    always @(posedge _791) begin
        if (_789)
            _3435 <= _3118;
        else
            _3435 <= _681;
    end
    assign _10663 = _8620 == _2231;
    assign _10660 = ~ _3920;
    assign _10661 = _3135 & _10660;
    assign _10664 = _10661 & _10663;
    assign _10665 = _10664 ? _5304 : _3432;
    assign _10658 = _5296 == _2231;
    assign _10659 = _5293 & _10658;
    assign _10667 = _10659 ? _2231 : _10665;
    assign _10669 = _805 ? _3118 : _10667;
    assign _682 = _10669;
    always @(posedge _791) begin
        if (_789)
            _3432 <= _3118;
        else
            _3432 <= _682;
    end
    assign _10676 = _8620 == _2240;
    assign _10673 = ~ _3920;
    assign _10674 = _3135 & _10673;
    assign _10677 = _10674 & _10676;
    assign _10678 = _10677 ? _5304 : _3429;
    assign _10671 = _5296 == _2240;
    assign _10672 = _5293 & _10671;
    assign _10680 = _10672 ? _2240 : _10678;
    assign _10682 = _805 ? _3118 : _10680;
    assign _683 = _10682;
    always @(posedge _791) begin
        if (_789)
            _3429 <= _3118;
        else
            _3429 <= _683;
    end
    assign _10689 = _8620 == _2249;
    assign _10686 = ~ _3920;
    assign _10687 = _3135 & _10686;
    assign _10690 = _10687 & _10689;
    assign _10691 = _10690 ? _5304 : _3426;
    assign _10684 = _5296 == _2249;
    assign _10685 = _5293 & _10684;
    assign _10693 = _10685 ? _2249 : _10691;
    assign _10695 = _805 ? _3118 : _10693;
    assign _684 = _10695;
    always @(posedge _791) begin
        if (_789)
            _3426 <= _3118;
        else
            _3426 <= _684;
    end
    assign _10702 = _8620 == _2258;
    assign _10699 = ~ _3920;
    assign _10700 = _3135 & _10699;
    assign _10703 = _10700 & _10702;
    assign _10704 = _10703 ? _5304 : _3423;
    assign _10697 = _5296 == _2258;
    assign _10698 = _5293 & _10697;
    assign _10706 = _10698 ? _2258 : _10704;
    assign _10708 = _805 ? _3118 : _10706;
    assign _685 = _10708;
    always @(posedge _791) begin
        if (_789)
            _3423 <= _3118;
        else
            _3423 <= _685;
    end
    assign _10715 = _8620 == _2267;
    assign _10712 = ~ _3920;
    assign _10713 = _3135 & _10712;
    assign _10716 = _10713 & _10715;
    assign _10717 = _10716 ? _5304 : _3420;
    assign _10710 = _5296 == _2267;
    assign _10711 = _5293 & _10710;
    assign _10719 = _10711 ? _2267 : _10717;
    assign _10721 = _805 ? _3118 : _10719;
    assign _686 = _10721;
    always @(posedge _791) begin
        if (_789)
            _3420 <= _3118;
        else
            _3420 <= _686;
    end
    assign _10728 = _8620 == _2276;
    assign _10725 = ~ _3920;
    assign _10726 = _3135 & _10725;
    assign _10729 = _10726 & _10728;
    assign _10730 = _10729 ? _5304 : _3417;
    assign _10723 = _5296 == _2276;
    assign _10724 = _5293 & _10723;
    assign _10732 = _10724 ? _2276 : _10730;
    assign _10734 = _805 ? _3118 : _10732;
    assign _687 = _10734;
    always @(posedge _791) begin
        if (_789)
            _3417 <= _3118;
        else
            _3417 <= _687;
    end
    assign _10741 = _8620 == _2285;
    assign _10738 = ~ _3920;
    assign _10739 = _3135 & _10738;
    assign _10742 = _10739 & _10741;
    assign _10743 = _10742 ? _5304 : _3414;
    assign _10736 = _5296 == _2285;
    assign _10737 = _5293 & _10736;
    assign _10745 = _10737 ? _2285 : _10743;
    assign _10747 = _805 ? _3118 : _10745;
    assign _688 = _10747;
    always @(posedge _791) begin
        if (_789)
            _3414 <= _3118;
        else
            _3414 <= _688;
    end
    assign _10754 = _8620 == _2294;
    assign _10751 = ~ _3920;
    assign _10752 = _3135 & _10751;
    assign _10755 = _10752 & _10754;
    assign _10756 = _10755 ? _5304 : _3411;
    assign _10749 = _5296 == _2294;
    assign _10750 = _5293 & _10749;
    assign _10758 = _10750 ? _2294 : _10756;
    assign _10760 = _805 ? _3118 : _10758;
    assign _689 = _10760;
    always @(posedge _791) begin
        if (_789)
            _3411 <= _3118;
        else
            _3411 <= _689;
    end
    assign _10767 = _8620 == _2303;
    assign _10764 = ~ _3920;
    assign _10765 = _3135 & _10764;
    assign _10768 = _10765 & _10767;
    assign _10769 = _10768 ? _5304 : _3408;
    assign _10762 = _5296 == _2303;
    assign _10763 = _5293 & _10762;
    assign _10771 = _10763 ? _2303 : _10769;
    assign _10773 = _805 ? _3118 : _10771;
    assign _690 = _10773;
    always @(posedge _791) begin
        if (_789)
            _3408 <= _3118;
        else
            _3408 <= _690;
    end
    assign _10780 = _8620 == _2312;
    assign _10777 = ~ _3920;
    assign _10778 = _3135 & _10777;
    assign _10781 = _10778 & _10780;
    assign _10782 = _10781 ? _5304 : _3405;
    assign _10775 = _5296 == _2312;
    assign _10776 = _5293 & _10775;
    assign _10784 = _10776 ? _2312 : _10782;
    assign _10786 = _805 ? _3118 : _10784;
    assign _691 = _10786;
    always @(posedge _791) begin
        if (_789)
            _3405 <= _3118;
        else
            _3405 <= _691;
    end
    assign _10793 = _8620 == _2321;
    assign _10790 = ~ _3920;
    assign _10791 = _3135 & _10790;
    assign _10794 = _10791 & _10793;
    assign _10795 = _10794 ? _5304 : _3402;
    assign _10788 = _5296 == _2321;
    assign _10789 = _5293 & _10788;
    assign _10797 = _10789 ? _2321 : _10795;
    assign _10799 = _805 ? _3118 : _10797;
    assign _692 = _10799;
    always @(posedge _791) begin
        if (_789)
            _3402 <= _3118;
        else
            _3402 <= _692;
    end
    assign _10806 = _8620 == _2330;
    assign _10803 = ~ _3920;
    assign _10804 = _3135 & _10803;
    assign _10807 = _10804 & _10806;
    assign _10808 = _10807 ? _5304 : _3399;
    assign _10801 = _5296 == _2330;
    assign _10802 = _5293 & _10801;
    assign _10810 = _10802 ? _2330 : _10808;
    assign _10812 = _805 ? _3118 : _10810;
    assign _693 = _10812;
    always @(posedge _791) begin
        if (_789)
            _3399 <= _3118;
        else
            _3399 <= _693;
    end
    assign _10819 = _8620 == _2339;
    assign _10816 = ~ _3920;
    assign _10817 = _3135 & _10816;
    assign _10820 = _10817 & _10819;
    assign _10821 = _10820 ? _5304 : _3396;
    assign _10814 = _5296 == _2339;
    assign _10815 = _5293 & _10814;
    assign _10823 = _10815 ? _2339 : _10821;
    assign _10825 = _805 ? _3118 : _10823;
    assign _694 = _10825;
    always @(posedge _791) begin
        if (_789)
            _3396 <= _3118;
        else
            _3396 <= _694;
    end
    assign _10832 = _8620 == _2348;
    assign _10829 = ~ _3920;
    assign _10830 = _3135 & _10829;
    assign _10833 = _10830 & _10832;
    assign _10834 = _10833 ? _5304 : _3393;
    assign _10827 = _5296 == _2348;
    assign _10828 = _5293 & _10827;
    assign _10836 = _10828 ? _2348 : _10834;
    assign _10838 = _805 ? _3118 : _10836;
    assign _695 = _10838;
    always @(posedge _791) begin
        if (_789)
            _3393 <= _3118;
        else
            _3393 <= _695;
    end
    assign _10845 = _8620 == _2357;
    assign _10842 = ~ _3920;
    assign _10843 = _3135 & _10842;
    assign _10846 = _10843 & _10845;
    assign _10847 = _10846 ? _5304 : _3390;
    assign _10840 = _5296 == _2357;
    assign _10841 = _5293 & _10840;
    assign _10849 = _10841 ? _2357 : _10847;
    assign _10851 = _805 ? _3118 : _10849;
    assign _696 = _10851;
    always @(posedge _791) begin
        if (_789)
            _3390 <= _3118;
        else
            _3390 <= _696;
    end
    assign _10858 = _8620 == _2366;
    assign _10855 = ~ _3920;
    assign _10856 = _3135 & _10855;
    assign _10859 = _10856 & _10858;
    assign _10860 = _10859 ? _5304 : _3387;
    assign _10853 = _5296 == _2366;
    assign _10854 = _5293 & _10853;
    assign _10862 = _10854 ? _2366 : _10860;
    assign _10864 = _805 ? _3118 : _10862;
    assign _697 = _10864;
    always @(posedge _791) begin
        if (_789)
            _3387 <= _3118;
        else
            _3387 <= _697;
    end
    assign _10871 = _8620 == _2375;
    assign _10868 = ~ _3920;
    assign _10869 = _3135 & _10868;
    assign _10872 = _10869 & _10871;
    assign _10873 = _10872 ? _5304 : _3384;
    assign _10866 = _5296 == _2375;
    assign _10867 = _5293 & _10866;
    assign _10875 = _10867 ? _2375 : _10873;
    assign _10877 = _805 ? _3118 : _10875;
    assign _698 = _10877;
    always @(posedge _791) begin
        if (_789)
            _3384 <= _3118;
        else
            _3384 <= _698;
    end
    assign _10884 = _8620 == _2384;
    assign _10881 = ~ _3920;
    assign _10882 = _3135 & _10881;
    assign _10885 = _10882 & _10884;
    assign _10886 = _10885 ? _5304 : _3381;
    assign _10879 = _5296 == _2384;
    assign _10880 = _5293 & _10879;
    assign _10888 = _10880 ? _2384 : _10886;
    assign _10890 = _805 ? _3118 : _10888;
    assign _699 = _10890;
    always @(posedge _791) begin
        if (_789)
            _3381 <= _3118;
        else
            _3381 <= _699;
    end
    assign _10897 = _8620 == _2393;
    assign _10894 = ~ _3920;
    assign _10895 = _3135 & _10894;
    assign _10898 = _10895 & _10897;
    assign _10899 = _10898 ? _5304 : _3378;
    assign _10892 = _5296 == _2393;
    assign _10893 = _5293 & _10892;
    assign _10901 = _10893 ? _2393 : _10899;
    assign _10903 = _805 ? _3118 : _10901;
    assign _700 = _10903;
    always @(posedge _791) begin
        if (_789)
            _3378 <= _3118;
        else
            _3378 <= _700;
    end
    assign _10910 = _8620 == _2402;
    assign _10907 = ~ _3920;
    assign _10908 = _3135 & _10907;
    assign _10911 = _10908 & _10910;
    assign _10912 = _10911 ? _5304 : _3375;
    assign _10905 = _5296 == _2402;
    assign _10906 = _5293 & _10905;
    assign _10914 = _10906 ? _2402 : _10912;
    assign _10916 = _805 ? _3118 : _10914;
    assign _701 = _10916;
    always @(posedge _791) begin
        if (_789)
            _3375 <= _3118;
        else
            _3375 <= _701;
    end
    assign _10923 = _8620 == _2411;
    assign _10920 = ~ _3920;
    assign _10921 = _3135 & _10920;
    assign _10924 = _10921 & _10923;
    assign _10925 = _10924 ? _5304 : _3372;
    assign _10918 = _5296 == _2411;
    assign _10919 = _5293 & _10918;
    assign _10927 = _10919 ? _2411 : _10925;
    assign _10929 = _805 ? _3118 : _10927;
    assign _702 = _10929;
    always @(posedge _791) begin
        if (_789)
            _3372 <= _3118;
        else
            _3372 <= _702;
    end
    assign _10936 = _8620 == _2420;
    assign _10933 = ~ _3920;
    assign _10934 = _3135 & _10933;
    assign _10937 = _10934 & _10936;
    assign _10938 = _10937 ? _5304 : _3369;
    assign _10931 = _5296 == _2420;
    assign _10932 = _5293 & _10931;
    assign _10940 = _10932 ? _2420 : _10938;
    assign _10942 = _805 ? _3118 : _10940;
    assign _703 = _10942;
    always @(posedge _791) begin
        if (_789)
            _3369 <= _3118;
        else
            _3369 <= _703;
    end
    assign _10949 = _8620 == _2429;
    assign _10946 = ~ _3920;
    assign _10947 = _3135 & _10946;
    assign _10950 = _10947 & _10949;
    assign _10951 = _10950 ? _5304 : _3366;
    assign _10944 = _5296 == _2429;
    assign _10945 = _5293 & _10944;
    assign _10953 = _10945 ? _2429 : _10951;
    assign _10955 = _805 ? _3118 : _10953;
    assign _704 = _10955;
    always @(posedge _791) begin
        if (_789)
            _3366 <= _3118;
        else
            _3366 <= _704;
    end
    assign _10962 = _8620 == _2438;
    assign _10959 = ~ _3920;
    assign _10960 = _3135 & _10959;
    assign _10963 = _10960 & _10962;
    assign _10964 = _10963 ? _5304 : _3363;
    assign _10957 = _5296 == _2438;
    assign _10958 = _5293 & _10957;
    assign _10966 = _10958 ? _2438 : _10964;
    assign _10968 = _805 ? _3118 : _10966;
    assign _705 = _10968;
    always @(posedge _791) begin
        if (_789)
            _3363 <= _3118;
        else
            _3363 <= _705;
    end
    assign _10975 = _8620 == _2447;
    assign _10972 = ~ _3920;
    assign _10973 = _3135 & _10972;
    assign _10976 = _10973 & _10975;
    assign _10977 = _10976 ? _5304 : _3360;
    assign _10970 = _5296 == _2447;
    assign _10971 = _5293 & _10970;
    assign _10979 = _10971 ? _2447 : _10977;
    assign _10981 = _805 ? _3118 : _10979;
    assign _706 = _10981;
    always @(posedge _791) begin
        if (_789)
            _3360 <= _3118;
        else
            _3360 <= _706;
    end
    assign _10988 = _8620 == _2456;
    assign _10985 = ~ _3920;
    assign _10986 = _3135 & _10985;
    assign _10989 = _10986 & _10988;
    assign _10990 = _10989 ? _5304 : _3357;
    assign _10983 = _5296 == _2456;
    assign _10984 = _5293 & _10983;
    assign _10992 = _10984 ? _2456 : _10990;
    assign _10994 = _805 ? _3118 : _10992;
    assign _707 = _10994;
    always @(posedge _791) begin
        if (_789)
            _3357 <= _3118;
        else
            _3357 <= _707;
    end
    assign _11001 = _8620 == _2465;
    assign _10998 = ~ _3920;
    assign _10999 = _3135 & _10998;
    assign _11002 = _10999 & _11001;
    assign _11003 = _11002 ? _5304 : _3354;
    assign _10996 = _5296 == _2465;
    assign _10997 = _5293 & _10996;
    assign _11005 = _10997 ? _2465 : _11003;
    assign _11007 = _805 ? _3118 : _11005;
    assign _708 = _11007;
    always @(posedge _791) begin
        if (_789)
            _3354 <= _3118;
        else
            _3354 <= _708;
    end
    assign _11014 = _8620 == _2474;
    assign _11011 = ~ _3920;
    assign _11012 = _3135 & _11011;
    assign _11015 = _11012 & _11014;
    assign _11016 = _11015 ? _5304 : _3351;
    assign _11009 = _5296 == _2474;
    assign _11010 = _5293 & _11009;
    assign _11018 = _11010 ? _2474 : _11016;
    assign _11020 = _805 ? _3118 : _11018;
    assign _709 = _11020;
    always @(posedge _791) begin
        if (_789)
            _3351 <= _3118;
        else
            _3351 <= _709;
    end
    assign _11027 = _8620 == _2483;
    assign _11024 = ~ _3920;
    assign _11025 = _3135 & _11024;
    assign _11028 = _11025 & _11027;
    assign _11029 = _11028 ? _5304 : _3348;
    assign _11022 = _5296 == _2483;
    assign _11023 = _5293 & _11022;
    assign _11031 = _11023 ? _2483 : _11029;
    assign _11033 = _805 ? _3118 : _11031;
    assign _710 = _11033;
    always @(posedge _791) begin
        if (_789)
            _3348 <= _3118;
        else
            _3348 <= _710;
    end
    assign _11040 = _8620 == _2492;
    assign _11037 = ~ _3920;
    assign _11038 = _3135 & _11037;
    assign _11041 = _11038 & _11040;
    assign _11042 = _11041 ? _5304 : _3345;
    assign _11035 = _5296 == _2492;
    assign _11036 = _5293 & _11035;
    assign _11044 = _11036 ? _2492 : _11042;
    assign _11046 = _805 ? _3118 : _11044;
    assign _711 = _11046;
    always @(posedge _791) begin
        if (_789)
            _3345 <= _3118;
        else
            _3345 <= _711;
    end
    assign _11053 = _8620 == _2501;
    assign _11050 = ~ _3920;
    assign _11051 = _3135 & _11050;
    assign _11054 = _11051 & _11053;
    assign _11055 = _11054 ? _5304 : _3342;
    assign _11048 = _5296 == _2501;
    assign _11049 = _5293 & _11048;
    assign _11057 = _11049 ? _2501 : _11055;
    assign _11059 = _805 ? _3118 : _11057;
    assign _712 = _11059;
    always @(posedge _791) begin
        if (_789)
            _3342 <= _3118;
        else
            _3342 <= _712;
    end
    assign _11066 = _8620 == _2510;
    assign _11063 = ~ _3920;
    assign _11064 = _3135 & _11063;
    assign _11067 = _11064 & _11066;
    assign _11068 = _11067 ? _5304 : _3339;
    assign _11061 = _5296 == _2510;
    assign _11062 = _5293 & _11061;
    assign _11070 = _11062 ? _2510 : _11068;
    assign _11072 = _805 ? _3118 : _11070;
    assign _713 = _11072;
    always @(posedge _791) begin
        if (_789)
            _3339 <= _3118;
        else
            _3339 <= _713;
    end
    assign _11079 = _8620 == _2519;
    assign _11076 = ~ _3920;
    assign _11077 = _3135 & _11076;
    assign _11080 = _11077 & _11079;
    assign _11081 = _11080 ? _5304 : _3336;
    assign _11074 = _5296 == _2519;
    assign _11075 = _5293 & _11074;
    assign _11083 = _11075 ? _2519 : _11081;
    assign _11085 = _805 ? _3118 : _11083;
    assign _714 = _11085;
    always @(posedge _791) begin
        if (_789)
            _3336 <= _3118;
        else
            _3336 <= _714;
    end
    assign _11092 = _8620 == _2528;
    assign _11089 = ~ _3920;
    assign _11090 = _3135 & _11089;
    assign _11093 = _11090 & _11092;
    assign _11094 = _11093 ? _5304 : _3333;
    assign _11087 = _5296 == _2528;
    assign _11088 = _5293 & _11087;
    assign _11096 = _11088 ? _2528 : _11094;
    assign _11098 = _805 ? _3118 : _11096;
    assign _715 = _11098;
    always @(posedge _791) begin
        if (_789)
            _3333 <= _3118;
        else
            _3333 <= _715;
    end
    assign _11105 = _8620 == _2537;
    assign _11102 = ~ _3920;
    assign _11103 = _3135 & _11102;
    assign _11106 = _11103 & _11105;
    assign _11107 = _11106 ? _5304 : _3330;
    assign _11100 = _5296 == _2537;
    assign _11101 = _5293 & _11100;
    assign _11109 = _11101 ? _2537 : _11107;
    assign _11111 = _805 ? _3118 : _11109;
    assign _716 = _11111;
    always @(posedge _791) begin
        if (_789)
            _3330 <= _3118;
        else
            _3330 <= _716;
    end
    assign _11118 = _8620 == _2546;
    assign _11115 = ~ _3920;
    assign _11116 = _3135 & _11115;
    assign _11119 = _11116 & _11118;
    assign _11120 = _11119 ? _5304 : _3327;
    assign _11113 = _5296 == _2546;
    assign _11114 = _5293 & _11113;
    assign _11122 = _11114 ? _2546 : _11120;
    assign _11124 = _805 ? _3118 : _11122;
    assign _717 = _11124;
    always @(posedge _791) begin
        if (_789)
            _3327 <= _3118;
        else
            _3327 <= _717;
    end
    assign _11131 = _8620 == _2555;
    assign _11128 = ~ _3920;
    assign _11129 = _3135 & _11128;
    assign _11132 = _11129 & _11131;
    assign _11133 = _11132 ? _5304 : _3324;
    assign _11126 = _5296 == _2555;
    assign _11127 = _5293 & _11126;
    assign _11135 = _11127 ? _2555 : _11133;
    assign _11137 = _805 ? _3118 : _11135;
    assign _718 = _11137;
    always @(posedge _791) begin
        if (_789)
            _3324 <= _3118;
        else
            _3324 <= _718;
    end
    assign _11144 = _8620 == _2564;
    assign _11141 = ~ _3920;
    assign _11142 = _3135 & _11141;
    assign _11145 = _11142 & _11144;
    assign _11146 = _11145 ? _5304 : _3321;
    assign _11139 = _5296 == _2564;
    assign _11140 = _5293 & _11139;
    assign _11148 = _11140 ? _2564 : _11146;
    assign _11150 = _805 ? _3118 : _11148;
    assign _719 = _11150;
    always @(posedge _791) begin
        if (_789)
            _3321 <= _3118;
        else
            _3321 <= _719;
    end
    assign _11157 = _8620 == _2573;
    assign _11154 = ~ _3920;
    assign _11155 = _3135 & _11154;
    assign _11158 = _11155 & _11157;
    assign _11159 = _11158 ? _5304 : _3318;
    assign _11152 = _5296 == _2573;
    assign _11153 = _5293 & _11152;
    assign _11161 = _11153 ? _2573 : _11159;
    assign _11163 = _805 ? _3118 : _11161;
    assign _720 = _11163;
    always @(posedge _791) begin
        if (_789)
            _3318 <= _3118;
        else
            _3318 <= _720;
    end
    assign _11170 = _8620 == _2582;
    assign _11167 = ~ _3920;
    assign _11168 = _3135 & _11167;
    assign _11171 = _11168 & _11170;
    assign _11172 = _11171 ? _5304 : _3315;
    assign _11165 = _5296 == _2582;
    assign _11166 = _5293 & _11165;
    assign _11174 = _11166 ? _2582 : _11172;
    assign _11176 = _805 ? _3118 : _11174;
    assign _721 = _11176;
    always @(posedge _791) begin
        if (_789)
            _3315 <= _3118;
        else
            _3315 <= _721;
    end
    assign _11183 = _8620 == _2591;
    assign _11180 = ~ _3920;
    assign _11181 = _3135 & _11180;
    assign _11184 = _11181 & _11183;
    assign _11185 = _11184 ? _5304 : _3312;
    assign _11178 = _5296 == _2591;
    assign _11179 = _5293 & _11178;
    assign _11187 = _11179 ? _2591 : _11185;
    assign _11189 = _805 ? _3118 : _11187;
    assign _722 = _11189;
    always @(posedge _791) begin
        if (_789)
            _3312 <= _3118;
        else
            _3312 <= _722;
    end
    assign _11196 = _8620 == _2600;
    assign _11193 = ~ _3920;
    assign _11194 = _3135 & _11193;
    assign _11197 = _11194 & _11196;
    assign _11198 = _11197 ? _5304 : _3309;
    assign _11191 = _5296 == _2600;
    assign _11192 = _5293 & _11191;
    assign _11200 = _11192 ? _2600 : _11198;
    assign _11202 = _805 ? _3118 : _11200;
    assign _723 = _11202;
    always @(posedge _791) begin
        if (_789)
            _3309 <= _3118;
        else
            _3309 <= _723;
    end
    assign _11209 = _8620 == _2609;
    assign _11206 = ~ _3920;
    assign _11207 = _3135 & _11206;
    assign _11210 = _11207 & _11209;
    assign _11211 = _11210 ? _5304 : _3306;
    assign _11204 = _5296 == _2609;
    assign _11205 = _5293 & _11204;
    assign _11213 = _11205 ? _2609 : _11211;
    assign _11215 = _805 ? _3118 : _11213;
    assign _724 = _11215;
    always @(posedge _791) begin
        if (_789)
            _3306 <= _3118;
        else
            _3306 <= _724;
    end
    assign _11222 = _8620 == _2618;
    assign _11219 = ~ _3920;
    assign _11220 = _3135 & _11219;
    assign _11223 = _11220 & _11222;
    assign _11224 = _11223 ? _5304 : _3303;
    assign _11217 = _5296 == _2618;
    assign _11218 = _5293 & _11217;
    assign _11226 = _11218 ? _2618 : _11224;
    assign _11228 = _805 ? _3118 : _11226;
    assign _725 = _11228;
    always @(posedge _791) begin
        if (_789)
            _3303 <= _3118;
        else
            _3303 <= _725;
    end
    assign _11235 = _8620 == _2627;
    assign _11232 = ~ _3920;
    assign _11233 = _3135 & _11232;
    assign _11236 = _11233 & _11235;
    assign _11237 = _11236 ? _5304 : _3300;
    assign _11230 = _5296 == _2627;
    assign _11231 = _5293 & _11230;
    assign _11239 = _11231 ? _2627 : _11237;
    assign _11241 = _805 ? _3118 : _11239;
    assign _726 = _11241;
    always @(posedge _791) begin
        if (_789)
            _3300 <= _3118;
        else
            _3300 <= _726;
    end
    assign _11248 = _8620 == _2636;
    assign _11245 = ~ _3920;
    assign _11246 = _3135 & _11245;
    assign _11249 = _11246 & _11248;
    assign _11250 = _11249 ? _5304 : _3297;
    assign _11243 = _5296 == _2636;
    assign _11244 = _5293 & _11243;
    assign _11252 = _11244 ? _2636 : _11250;
    assign _11254 = _805 ? _3118 : _11252;
    assign _727 = _11254;
    always @(posedge _791) begin
        if (_789)
            _3297 <= _3118;
        else
            _3297 <= _727;
    end
    assign _11261 = _8620 == _2645;
    assign _11258 = ~ _3920;
    assign _11259 = _3135 & _11258;
    assign _11262 = _11259 & _11261;
    assign _11263 = _11262 ? _5304 : _3294;
    assign _11256 = _5296 == _2645;
    assign _11257 = _5293 & _11256;
    assign _11265 = _11257 ? _2645 : _11263;
    assign _11267 = _805 ? _3118 : _11265;
    assign _728 = _11267;
    always @(posedge _791) begin
        if (_789)
            _3294 <= _3118;
        else
            _3294 <= _728;
    end
    assign _11274 = _8620 == _2654;
    assign _11271 = ~ _3920;
    assign _11272 = _3135 & _11271;
    assign _11275 = _11272 & _11274;
    assign _11276 = _11275 ? _5304 : _3291;
    assign _11269 = _5296 == _2654;
    assign _11270 = _5293 & _11269;
    assign _11278 = _11270 ? _2654 : _11276;
    assign _11280 = _805 ? _3118 : _11278;
    assign _729 = _11280;
    always @(posedge _791) begin
        if (_789)
            _3291 <= _3118;
        else
            _3291 <= _729;
    end
    assign _11287 = _8620 == _2663;
    assign _11284 = ~ _3920;
    assign _11285 = _3135 & _11284;
    assign _11288 = _11285 & _11287;
    assign _11289 = _11288 ? _5304 : _3288;
    assign _11282 = _5296 == _2663;
    assign _11283 = _5293 & _11282;
    assign _11291 = _11283 ? _2663 : _11289;
    assign _11293 = _805 ? _3118 : _11291;
    assign _730 = _11293;
    always @(posedge _791) begin
        if (_789)
            _3288 <= _3118;
        else
            _3288 <= _730;
    end
    assign _11300 = _8620 == _2672;
    assign _11297 = ~ _3920;
    assign _11298 = _3135 & _11297;
    assign _11301 = _11298 & _11300;
    assign _11302 = _11301 ? _5304 : _3285;
    assign _11295 = _5296 == _2672;
    assign _11296 = _5293 & _11295;
    assign _11304 = _11296 ? _2672 : _11302;
    assign _11306 = _805 ? _3118 : _11304;
    assign _731 = _11306;
    always @(posedge _791) begin
        if (_789)
            _3285 <= _3118;
        else
            _3285 <= _731;
    end
    assign _11313 = _8620 == _2681;
    assign _11310 = ~ _3920;
    assign _11311 = _3135 & _11310;
    assign _11314 = _11311 & _11313;
    assign _11315 = _11314 ? _5304 : _3282;
    assign _11308 = _5296 == _2681;
    assign _11309 = _5293 & _11308;
    assign _11317 = _11309 ? _2681 : _11315;
    assign _11319 = _805 ? _3118 : _11317;
    assign _732 = _11319;
    always @(posedge _791) begin
        if (_789)
            _3282 <= _3118;
        else
            _3282 <= _732;
    end
    assign _11326 = _8620 == _2690;
    assign _11323 = ~ _3920;
    assign _11324 = _3135 & _11323;
    assign _11327 = _11324 & _11326;
    assign _11328 = _11327 ? _5304 : _3279;
    assign _11321 = _5296 == _2690;
    assign _11322 = _5293 & _11321;
    assign _11330 = _11322 ? _2690 : _11328;
    assign _11332 = _805 ? _3118 : _11330;
    assign _733 = _11332;
    always @(posedge _791) begin
        if (_789)
            _3279 <= _3118;
        else
            _3279 <= _733;
    end
    assign _11339 = _8620 == _2699;
    assign _11336 = ~ _3920;
    assign _11337 = _3135 & _11336;
    assign _11340 = _11337 & _11339;
    assign _11341 = _11340 ? _5304 : _3276;
    assign _11334 = _5296 == _2699;
    assign _11335 = _5293 & _11334;
    assign _11343 = _11335 ? _2699 : _11341;
    assign _11345 = _805 ? _3118 : _11343;
    assign _734 = _11345;
    always @(posedge _791) begin
        if (_789)
            _3276 <= _3118;
        else
            _3276 <= _734;
    end
    assign _11352 = _8620 == _2708;
    assign _11349 = ~ _3920;
    assign _11350 = _3135 & _11349;
    assign _11353 = _11350 & _11352;
    assign _11354 = _11353 ? _5304 : _3273;
    assign _11347 = _5296 == _2708;
    assign _11348 = _5293 & _11347;
    assign _11356 = _11348 ? _2708 : _11354;
    assign _11358 = _805 ? _3118 : _11356;
    assign _735 = _11358;
    always @(posedge _791) begin
        if (_789)
            _3273 <= _3118;
        else
            _3273 <= _735;
    end
    assign _11365 = _8620 == _2717;
    assign _11362 = ~ _3920;
    assign _11363 = _3135 & _11362;
    assign _11366 = _11363 & _11365;
    assign _11367 = _11366 ? _5304 : _3270;
    assign _11360 = _5296 == _2717;
    assign _11361 = _5293 & _11360;
    assign _11369 = _11361 ? _2717 : _11367;
    assign _11371 = _805 ? _3118 : _11369;
    assign _736 = _11371;
    always @(posedge _791) begin
        if (_789)
            _3270 <= _3118;
        else
            _3270 <= _736;
    end
    assign _11378 = _8620 == _2726;
    assign _11375 = ~ _3920;
    assign _11376 = _3135 & _11375;
    assign _11379 = _11376 & _11378;
    assign _11380 = _11379 ? _5304 : _3267;
    assign _11373 = _5296 == _2726;
    assign _11374 = _5293 & _11373;
    assign _11382 = _11374 ? _2726 : _11380;
    assign _11384 = _805 ? _3118 : _11382;
    assign _737 = _11384;
    always @(posedge _791) begin
        if (_789)
            _3267 <= _3118;
        else
            _3267 <= _737;
    end
    assign _11391 = _8620 == _2735;
    assign _11388 = ~ _3920;
    assign _11389 = _3135 & _11388;
    assign _11392 = _11389 & _11391;
    assign _11393 = _11392 ? _5304 : _3264;
    assign _11386 = _5296 == _2735;
    assign _11387 = _5293 & _11386;
    assign _11395 = _11387 ? _2735 : _11393;
    assign _11397 = _805 ? _3118 : _11395;
    assign _738 = _11397;
    always @(posedge _791) begin
        if (_789)
            _3264 <= _3118;
        else
            _3264 <= _738;
    end
    assign _11404 = _8620 == _2744;
    assign _11401 = ~ _3920;
    assign _11402 = _3135 & _11401;
    assign _11405 = _11402 & _11404;
    assign _11406 = _11405 ? _5304 : _3261;
    assign _11399 = _5296 == _2744;
    assign _11400 = _5293 & _11399;
    assign _11408 = _11400 ? _2744 : _11406;
    assign _11410 = _805 ? _3118 : _11408;
    assign _739 = _11410;
    always @(posedge _791) begin
        if (_789)
            _3261 <= _3118;
        else
            _3261 <= _739;
    end
    assign _11417 = _8620 == _2753;
    assign _11414 = ~ _3920;
    assign _11415 = _3135 & _11414;
    assign _11418 = _11415 & _11417;
    assign _11419 = _11418 ? _5304 : _3258;
    assign _11412 = _5296 == _2753;
    assign _11413 = _5293 & _11412;
    assign _11421 = _11413 ? _2753 : _11419;
    assign _11423 = _805 ? _3118 : _11421;
    assign _740 = _11423;
    always @(posedge _791) begin
        if (_789)
            _3258 <= _3118;
        else
            _3258 <= _740;
    end
    assign _11430 = _8620 == _2762;
    assign _11427 = ~ _3920;
    assign _11428 = _3135 & _11427;
    assign _11431 = _11428 & _11430;
    assign _11432 = _11431 ? _5304 : _3255;
    assign _11425 = _5296 == _2762;
    assign _11426 = _5293 & _11425;
    assign _11434 = _11426 ? _2762 : _11432;
    assign _11436 = _805 ? _3118 : _11434;
    assign _741 = _11436;
    always @(posedge _791) begin
        if (_789)
            _3255 <= _3118;
        else
            _3255 <= _741;
    end
    assign _11443 = _8620 == _2771;
    assign _11440 = ~ _3920;
    assign _11441 = _3135 & _11440;
    assign _11444 = _11441 & _11443;
    assign _11445 = _11444 ? _5304 : _3252;
    assign _11438 = _5296 == _2771;
    assign _11439 = _5293 & _11438;
    assign _11447 = _11439 ? _2771 : _11445;
    assign _11449 = _805 ? _3118 : _11447;
    assign _742 = _11449;
    always @(posedge _791) begin
        if (_789)
            _3252 <= _3118;
        else
            _3252 <= _742;
    end
    assign _11456 = _8620 == _2780;
    assign _11453 = ~ _3920;
    assign _11454 = _3135 & _11453;
    assign _11457 = _11454 & _11456;
    assign _11458 = _11457 ? _5304 : _3249;
    assign _11451 = _5296 == _2780;
    assign _11452 = _5293 & _11451;
    assign _11460 = _11452 ? _2780 : _11458;
    assign _11462 = _805 ? _3118 : _11460;
    assign _743 = _11462;
    always @(posedge _791) begin
        if (_789)
            _3249 <= _3118;
        else
            _3249 <= _743;
    end
    assign _11469 = _8620 == _2789;
    assign _11466 = ~ _3920;
    assign _11467 = _3135 & _11466;
    assign _11470 = _11467 & _11469;
    assign _11471 = _11470 ? _5304 : _3246;
    assign _11464 = _5296 == _2789;
    assign _11465 = _5293 & _11464;
    assign _11473 = _11465 ? _2789 : _11471;
    assign _11475 = _805 ? _3118 : _11473;
    assign _744 = _11475;
    always @(posedge _791) begin
        if (_789)
            _3246 <= _3118;
        else
            _3246 <= _744;
    end
    assign _11482 = _8620 == _2798;
    assign _11479 = ~ _3920;
    assign _11480 = _3135 & _11479;
    assign _11483 = _11480 & _11482;
    assign _11484 = _11483 ? _5304 : _3243;
    assign _11477 = _5296 == _2798;
    assign _11478 = _5293 & _11477;
    assign _11486 = _11478 ? _2798 : _11484;
    assign _11488 = _805 ? _3118 : _11486;
    assign _745 = _11488;
    always @(posedge _791) begin
        if (_789)
            _3243 <= _3118;
        else
            _3243 <= _745;
    end
    assign _11495 = _8620 == _2807;
    assign _11492 = ~ _3920;
    assign _11493 = _3135 & _11492;
    assign _11496 = _11493 & _11495;
    assign _11497 = _11496 ? _5304 : _3240;
    assign _11490 = _5296 == _2807;
    assign _11491 = _5293 & _11490;
    assign _11499 = _11491 ? _2807 : _11497;
    assign _11501 = _805 ? _3118 : _11499;
    assign _746 = _11501;
    always @(posedge _791) begin
        if (_789)
            _3240 <= _3118;
        else
            _3240 <= _746;
    end
    assign _11508 = _8620 == _2816;
    assign _11505 = ~ _3920;
    assign _11506 = _3135 & _11505;
    assign _11509 = _11506 & _11508;
    assign _11510 = _11509 ? _5304 : _3237;
    assign _11503 = _5296 == _2816;
    assign _11504 = _5293 & _11503;
    assign _11512 = _11504 ? _2816 : _11510;
    assign _11514 = _805 ? _3118 : _11512;
    assign _747 = _11514;
    always @(posedge _791) begin
        if (_789)
            _3237 <= _3118;
        else
            _3237 <= _747;
    end
    assign _11521 = _8620 == _2825;
    assign _11518 = ~ _3920;
    assign _11519 = _3135 & _11518;
    assign _11522 = _11519 & _11521;
    assign _11523 = _11522 ? _5304 : _3234;
    assign _11516 = _5296 == _2825;
    assign _11517 = _5293 & _11516;
    assign _11525 = _11517 ? _2825 : _11523;
    assign _11527 = _805 ? _3118 : _11525;
    assign _748 = _11527;
    always @(posedge _791) begin
        if (_789)
            _3234 <= _3118;
        else
            _3234 <= _748;
    end
    assign _11534 = _8620 == _2834;
    assign _11531 = ~ _3920;
    assign _11532 = _3135 & _11531;
    assign _11535 = _11532 & _11534;
    assign _11536 = _11535 ? _5304 : _3231;
    assign _11529 = _5296 == _2834;
    assign _11530 = _5293 & _11529;
    assign _11538 = _11530 ? _2834 : _11536;
    assign _11540 = _805 ? _3118 : _11538;
    assign _749 = _11540;
    always @(posedge _791) begin
        if (_789)
            _3231 <= _3118;
        else
            _3231 <= _749;
    end
    assign _11547 = _8620 == _2843;
    assign _11544 = ~ _3920;
    assign _11545 = _3135 & _11544;
    assign _11548 = _11545 & _11547;
    assign _11549 = _11548 ? _5304 : _3228;
    assign _11542 = _5296 == _2843;
    assign _11543 = _5293 & _11542;
    assign _11551 = _11543 ? _2843 : _11549;
    assign _11553 = _805 ? _3118 : _11551;
    assign _750 = _11553;
    always @(posedge _791) begin
        if (_789)
            _3228 <= _3118;
        else
            _3228 <= _750;
    end
    assign _11560 = _8620 == _2852;
    assign _11557 = ~ _3920;
    assign _11558 = _3135 & _11557;
    assign _11561 = _11558 & _11560;
    assign _11562 = _11561 ? _5304 : _3225;
    assign _11555 = _5296 == _2852;
    assign _11556 = _5293 & _11555;
    assign _11564 = _11556 ? _2852 : _11562;
    assign _11566 = _805 ? _3118 : _11564;
    assign _751 = _11566;
    always @(posedge _791) begin
        if (_789)
            _3225 <= _3118;
        else
            _3225 <= _751;
    end
    assign _11573 = _8620 == _2861;
    assign _11570 = ~ _3920;
    assign _11571 = _3135 & _11570;
    assign _11574 = _11571 & _11573;
    assign _11575 = _11574 ? _5304 : _3222;
    assign _11568 = _5296 == _2861;
    assign _11569 = _5293 & _11568;
    assign _11577 = _11569 ? _2861 : _11575;
    assign _11579 = _805 ? _3118 : _11577;
    assign _752 = _11579;
    always @(posedge _791) begin
        if (_789)
            _3222 <= _3118;
        else
            _3222 <= _752;
    end
    assign _11586 = _8620 == _2870;
    assign _11583 = ~ _3920;
    assign _11584 = _3135 & _11583;
    assign _11587 = _11584 & _11586;
    assign _11588 = _11587 ? _5304 : _3219;
    assign _11581 = _5296 == _2870;
    assign _11582 = _5293 & _11581;
    assign _11590 = _11582 ? _2870 : _11588;
    assign _11592 = _805 ? _3118 : _11590;
    assign _753 = _11592;
    always @(posedge _791) begin
        if (_789)
            _3219 <= _3118;
        else
            _3219 <= _753;
    end
    assign _11599 = _8620 == _2879;
    assign _11596 = ~ _3920;
    assign _11597 = _3135 & _11596;
    assign _11600 = _11597 & _11599;
    assign _11601 = _11600 ? _5304 : _3216;
    assign _11594 = _5296 == _2879;
    assign _11595 = _5293 & _11594;
    assign _11603 = _11595 ? _2879 : _11601;
    assign _11605 = _805 ? _3118 : _11603;
    assign _754 = _11605;
    always @(posedge _791) begin
        if (_789)
            _3216 <= _3118;
        else
            _3216 <= _754;
    end
    assign _11612 = _8620 == _2888;
    assign _11609 = ~ _3920;
    assign _11610 = _3135 & _11609;
    assign _11613 = _11610 & _11612;
    assign _11614 = _11613 ? _5304 : _3213;
    assign _11607 = _5296 == _2888;
    assign _11608 = _5293 & _11607;
    assign _11616 = _11608 ? _2888 : _11614;
    assign _11618 = _805 ? _3118 : _11616;
    assign _755 = _11618;
    always @(posedge _791) begin
        if (_789)
            _3213 <= _3118;
        else
            _3213 <= _755;
    end
    assign _11625 = _8620 == _2897;
    assign _11622 = ~ _3920;
    assign _11623 = _3135 & _11622;
    assign _11626 = _11623 & _11625;
    assign _11627 = _11626 ? _5304 : _3210;
    assign _11620 = _5296 == _2897;
    assign _11621 = _5293 & _11620;
    assign _11629 = _11621 ? _2897 : _11627;
    assign _11631 = _805 ? _3118 : _11629;
    assign _756 = _11631;
    always @(posedge _791) begin
        if (_789)
            _3210 <= _3118;
        else
            _3210 <= _756;
    end
    assign _11638 = _8620 == _2906;
    assign _11635 = ~ _3920;
    assign _11636 = _3135 & _11635;
    assign _11639 = _11636 & _11638;
    assign _11640 = _11639 ? _5304 : _3207;
    assign _11633 = _5296 == _2906;
    assign _11634 = _5293 & _11633;
    assign _11642 = _11634 ? _2906 : _11640;
    assign _11644 = _805 ? _3118 : _11642;
    assign _757 = _11644;
    always @(posedge _791) begin
        if (_789)
            _3207 <= _3118;
        else
            _3207 <= _757;
    end
    assign _11651 = _8620 == _2915;
    assign _11648 = ~ _3920;
    assign _11649 = _3135 & _11648;
    assign _11652 = _11649 & _11651;
    assign _11653 = _11652 ? _5304 : _3204;
    assign _11646 = _5296 == _2915;
    assign _11647 = _5293 & _11646;
    assign _11655 = _11647 ? _2915 : _11653;
    assign _11657 = _805 ? _3118 : _11655;
    assign _758 = _11657;
    always @(posedge _791) begin
        if (_789)
            _3204 <= _3118;
        else
            _3204 <= _758;
    end
    assign _11664 = _8620 == _2924;
    assign _11661 = ~ _3920;
    assign _11662 = _3135 & _11661;
    assign _11665 = _11662 & _11664;
    assign _11666 = _11665 ? _5304 : _3201;
    assign _11659 = _5296 == _2924;
    assign _11660 = _5293 & _11659;
    assign _11668 = _11660 ? _2924 : _11666;
    assign _11670 = _805 ? _3118 : _11668;
    assign _759 = _11670;
    always @(posedge _791) begin
        if (_789)
            _3201 <= _3118;
        else
            _3201 <= _759;
    end
    assign _11677 = _8620 == _2933;
    assign _11674 = ~ _3920;
    assign _11675 = _3135 & _11674;
    assign _11678 = _11675 & _11677;
    assign _11679 = _11678 ? _5304 : _3198;
    assign _11672 = _5296 == _2933;
    assign _11673 = _5293 & _11672;
    assign _11681 = _11673 ? _2933 : _11679;
    assign _11683 = _805 ? _3118 : _11681;
    assign _760 = _11683;
    always @(posedge _791) begin
        if (_789)
            _3198 <= _3118;
        else
            _3198 <= _760;
    end
    assign _11690 = _8620 == _2942;
    assign _11687 = ~ _3920;
    assign _11688 = _3135 & _11687;
    assign _11691 = _11688 & _11690;
    assign _11692 = _11691 ? _5304 : _3195;
    assign _11685 = _5296 == _2942;
    assign _11686 = _5293 & _11685;
    assign _11694 = _11686 ? _2942 : _11692;
    assign _11696 = _805 ? _3118 : _11694;
    assign _761 = _11696;
    always @(posedge _791) begin
        if (_789)
            _3195 <= _3118;
        else
            _3195 <= _761;
    end
    assign _11703 = _8620 == _2951;
    assign _11700 = ~ _3920;
    assign _11701 = _3135 & _11700;
    assign _11704 = _11701 & _11703;
    assign _11705 = _11704 ? _5304 : _3192;
    assign _11698 = _5296 == _2951;
    assign _11699 = _5293 & _11698;
    assign _11707 = _11699 ? _2951 : _11705;
    assign _11709 = _805 ? _3118 : _11707;
    assign _762 = _11709;
    always @(posedge _791) begin
        if (_789)
            _3192 <= _3118;
        else
            _3192 <= _762;
    end
    assign _11716 = _8620 == _2960;
    assign _11713 = ~ _3920;
    assign _11714 = _3135 & _11713;
    assign _11717 = _11714 & _11716;
    assign _11718 = _11717 ? _5304 : _3189;
    assign _11711 = _5296 == _2960;
    assign _11712 = _5293 & _11711;
    assign _11720 = _11712 ? _2960 : _11718;
    assign _11722 = _805 ? _3118 : _11720;
    assign _763 = _11722;
    always @(posedge _791) begin
        if (_789)
            _3189 <= _3118;
        else
            _3189 <= _763;
    end
    assign _11729 = _8620 == _2969;
    assign _11726 = ~ _3920;
    assign _11727 = _3135 & _11726;
    assign _11730 = _11727 & _11729;
    assign _11731 = _11730 ? _5304 : _3186;
    assign _11724 = _5296 == _2969;
    assign _11725 = _5293 & _11724;
    assign _11733 = _11725 ? _2969 : _11731;
    assign _11735 = _805 ? _3118 : _11733;
    assign _764 = _11735;
    always @(posedge _791) begin
        if (_789)
            _3186 <= _3118;
        else
            _3186 <= _764;
    end
    assign _11742 = _8620 == _2978;
    assign _11739 = ~ _3920;
    assign _11740 = _3135 & _11739;
    assign _11743 = _11740 & _11742;
    assign _11744 = _11743 ? _5304 : _3183;
    assign _11737 = _5296 == _2978;
    assign _11738 = _5293 & _11737;
    assign _11746 = _11738 ? _2978 : _11744;
    assign _11748 = _805 ? _3118 : _11746;
    assign _765 = _11748;
    always @(posedge _791) begin
        if (_789)
            _3183 <= _3118;
        else
            _3183 <= _765;
    end
    assign _11755 = _8620 == _2987;
    assign _11752 = ~ _3920;
    assign _11753 = _3135 & _11752;
    assign _11756 = _11753 & _11755;
    assign _11757 = _11756 ? _5304 : _3180;
    assign _11750 = _5296 == _2987;
    assign _11751 = _5293 & _11750;
    assign _11759 = _11751 ? _2987 : _11757;
    assign _11761 = _805 ? _3118 : _11759;
    assign _766 = _11761;
    always @(posedge _791) begin
        if (_789)
            _3180 <= _3118;
        else
            _3180 <= _766;
    end
    assign _11768 = _8620 == _2996;
    assign _11765 = ~ _3920;
    assign _11766 = _3135 & _11765;
    assign _11769 = _11766 & _11768;
    assign _11770 = _11769 ? _5304 : _3177;
    assign _11763 = _5296 == _2996;
    assign _11764 = _5293 & _11763;
    assign _11772 = _11764 ? _2996 : _11770;
    assign _11774 = _805 ? _3118 : _11772;
    assign _767 = _11774;
    always @(posedge _791) begin
        if (_789)
            _3177 <= _3118;
        else
            _3177 <= _767;
    end
    assign _11781 = _8620 == _3005;
    assign _11778 = ~ _3920;
    assign _11779 = _3135 & _11778;
    assign _11782 = _11779 & _11781;
    assign _11783 = _11782 ? _5304 : _3174;
    assign _11776 = _5296 == _3005;
    assign _11777 = _5293 & _11776;
    assign _11785 = _11777 ? _3005 : _11783;
    assign _11787 = _805 ? _3118 : _11785;
    assign _768 = _11787;
    always @(posedge _791) begin
        if (_789)
            _3174 <= _3118;
        else
            _3174 <= _768;
    end
    assign _11794 = _8620 == _3014;
    assign _11791 = ~ _3920;
    assign _11792 = _3135 & _11791;
    assign _11795 = _11792 & _11794;
    assign _11796 = _11795 ? _5304 : _3171;
    assign _11789 = _5296 == _3014;
    assign _11790 = _5293 & _11789;
    assign _11798 = _11790 ? _3014 : _11796;
    assign _11800 = _805 ? _3118 : _11798;
    assign _769 = _11800;
    always @(posedge _791) begin
        if (_789)
            _3171 <= _3118;
        else
            _3171 <= _769;
    end
    assign _11807 = _8620 == _3023;
    assign _11804 = ~ _3920;
    assign _11805 = _3135 & _11804;
    assign _11808 = _11805 & _11807;
    assign _11809 = _11808 ? _5304 : _3168;
    assign _11802 = _5296 == _3023;
    assign _11803 = _5293 & _11802;
    assign _11811 = _11803 ? _3023 : _11809;
    assign _11813 = _805 ? _3118 : _11811;
    assign _770 = _11813;
    always @(posedge _791) begin
        if (_789)
            _3168 <= _3118;
        else
            _3168 <= _770;
    end
    assign _11820 = _8620 == _3032;
    assign _11817 = ~ _3920;
    assign _11818 = _3135 & _11817;
    assign _11821 = _11818 & _11820;
    assign _11822 = _11821 ? _5304 : _3165;
    assign _11815 = _5296 == _3032;
    assign _11816 = _5293 & _11815;
    assign _11824 = _11816 ? _3032 : _11822;
    assign _11826 = _805 ? _3118 : _11824;
    assign _771 = _11826;
    always @(posedge _791) begin
        if (_789)
            _3165 <= _3118;
        else
            _3165 <= _771;
    end
    assign _11833 = _8620 == _3041;
    assign _11830 = ~ _3920;
    assign _11831 = _3135 & _11830;
    assign _11834 = _11831 & _11833;
    assign _11835 = _11834 ? _5304 : _3162;
    assign _11828 = _5296 == _3041;
    assign _11829 = _5293 & _11828;
    assign _11837 = _11829 ? _3041 : _11835;
    assign _11839 = _805 ? _3118 : _11837;
    assign _772 = _11839;
    always @(posedge _791) begin
        if (_789)
            _3162 <= _3118;
        else
            _3162 <= _772;
    end
    assign _11846 = _8620 == _3050;
    assign _11843 = ~ _3920;
    assign _11844 = _3135 & _11843;
    assign _11847 = _11844 & _11846;
    assign _11848 = _11847 ? _5304 : _3159;
    assign _11841 = _5296 == _3050;
    assign _11842 = _5293 & _11841;
    assign _11850 = _11842 ? _3050 : _11848;
    assign _11852 = _805 ? _3118 : _11850;
    assign _773 = _11852;
    always @(posedge _791) begin
        if (_789)
            _3159 <= _3118;
        else
            _3159 <= _773;
    end
    assign _11859 = _8620 == _3059;
    assign _11856 = ~ _3920;
    assign _11857 = _3135 & _11856;
    assign _11860 = _11857 & _11859;
    assign _11861 = _11860 ? _5304 : _3156;
    assign _11854 = _5296 == _3059;
    assign _11855 = _5293 & _11854;
    assign _11863 = _11855 ? _3059 : _11861;
    assign _11865 = _805 ? _3118 : _11863;
    assign _774 = _11865;
    always @(posedge _791) begin
        if (_789)
            _3156 <= _3118;
        else
            _3156 <= _774;
    end
    assign _11872 = _8620 == _3068;
    assign _11869 = ~ _3920;
    assign _11870 = _3135 & _11869;
    assign _11873 = _11870 & _11872;
    assign _11874 = _11873 ? _5304 : _3153;
    assign _11867 = _5296 == _3068;
    assign _11868 = _5293 & _11867;
    assign _11876 = _11868 ? _3068 : _11874;
    assign _11878 = _805 ? _3118 : _11876;
    assign _775 = _11878;
    always @(posedge _791) begin
        if (_789)
            _3153 <= _3118;
        else
            _3153 <= _775;
    end
    assign _11885 = _8620 == _3077;
    assign _11882 = ~ _3920;
    assign _11883 = _3135 & _11882;
    assign _11886 = _11883 & _11885;
    assign _11887 = _11886 ? _5304 : _3150;
    assign _11880 = _5296 == _3077;
    assign _11881 = _5293 & _11880;
    assign _11889 = _11881 ? _3077 : _11887;
    assign _11891 = _805 ? _3118 : _11889;
    assign _776 = _11891;
    always @(posedge _791) begin
        if (_789)
            _3150 <= _3118;
        else
            _3150 <= _776;
    end
    assign _11898 = _8620 == _3086;
    assign _11895 = ~ _3920;
    assign _11896 = _3135 & _11895;
    assign _11899 = _11896 & _11898;
    assign _11900 = _11899 ? _5304 : _3147;
    assign _11893 = _5296 == _3086;
    assign _11894 = _5293 & _11893;
    assign _11902 = _11894 ? _3086 : _11900;
    assign _11904 = _805 ? _3118 : _11902;
    assign _777 = _11904;
    always @(posedge _791) begin
        if (_789)
            _3147 <= _3118;
        else
            _3147 <= _777;
    end
    assign _11911 = _8620 == _3095;
    assign _11908 = ~ _3920;
    assign _11909 = _3135 & _11908;
    assign _11912 = _11909 & _11911;
    assign _11913 = _11912 ? _5304 : _3144;
    assign _11906 = _5296 == _3095;
    assign _11907 = _5293 & _11906;
    assign _11915 = _11907 ? _3095 : _11913;
    assign _11917 = _805 ? _3118 : _11915;
    assign _778 = _11917;
    always @(posedge _791) begin
        if (_789)
            _3144 <= _3118;
        else
            _3144 <= _778;
    end
    assign _11924 = _8620 == _3104;
    assign _11921 = ~ _3920;
    assign _11922 = _3135 & _11921;
    assign _11925 = _11922 & _11924;
    assign _11926 = _11925 ? _5304 : _3141;
    assign _11919 = _5296 == _3104;
    assign _11920 = _5293 & _11919;
    assign _11928 = _11920 ? _3104 : _11926;
    assign _11930 = _805 ? _3118 : _11928;
    assign _779 = _11930;
    always @(posedge _791) begin
        if (_789)
            _3141 <= _3118;
        else
            _3141 <= _779;
    end
    assign _781 = edge_j;
    always @* begin
        case (_781)
        0:
            _3912 <= _3138;
        1:
            _3912 <= _3141;
        2:
            _3912 <= _3144;
        3:
            _3912 <= _3147;
        4:
            _3912 <= _3150;
        5:
            _3912 <= _3153;
        6:
            _3912 <= _3156;
        7:
            _3912 <= _3159;
        8:
            _3912 <= _3162;
        9:
            _3912 <= _3165;
        10:
            _3912 <= _3168;
        11:
            _3912 <= _3171;
        12:
            _3912 <= _3174;
        13:
            _3912 <= _3177;
        14:
            _3912 <= _3180;
        15:
            _3912 <= _3183;
        16:
            _3912 <= _3186;
        17:
            _3912 <= _3189;
        18:
            _3912 <= _3192;
        19:
            _3912 <= _3195;
        20:
            _3912 <= _3198;
        21:
            _3912 <= _3201;
        22:
            _3912 <= _3204;
        23:
            _3912 <= _3207;
        24:
            _3912 <= _3210;
        25:
            _3912 <= _3213;
        26:
            _3912 <= _3216;
        27:
            _3912 <= _3219;
        28:
            _3912 <= _3222;
        29:
            _3912 <= _3225;
        30:
            _3912 <= _3228;
        31:
            _3912 <= _3231;
        32:
            _3912 <= _3234;
        33:
            _3912 <= _3237;
        34:
            _3912 <= _3240;
        35:
            _3912 <= _3243;
        36:
            _3912 <= _3246;
        37:
            _3912 <= _3249;
        38:
            _3912 <= _3252;
        39:
            _3912 <= _3255;
        40:
            _3912 <= _3258;
        41:
            _3912 <= _3261;
        42:
            _3912 <= _3264;
        43:
            _3912 <= _3267;
        44:
            _3912 <= _3270;
        45:
            _3912 <= _3273;
        46:
            _3912 <= _3276;
        47:
            _3912 <= _3279;
        48:
            _3912 <= _3282;
        49:
            _3912 <= _3285;
        50:
            _3912 <= _3288;
        51:
            _3912 <= _3291;
        52:
            _3912 <= _3294;
        53:
            _3912 <= _3297;
        54:
            _3912 <= _3300;
        55:
            _3912 <= _3303;
        56:
            _3912 <= _3306;
        57:
            _3912 <= _3309;
        58:
            _3912 <= _3312;
        59:
            _3912 <= _3315;
        60:
            _3912 <= _3318;
        61:
            _3912 <= _3321;
        62:
            _3912 <= _3324;
        63:
            _3912 <= _3327;
        64:
            _3912 <= _3330;
        65:
            _3912 <= _3333;
        66:
            _3912 <= _3336;
        67:
            _3912 <= _3339;
        68:
            _3912 <= _3342;
        69:
            _3912 <= _3345;
        70:
            _3912 <= _3348;
        71:
            _3912 <= _3351;
        72:
            _3912 <= _3354;
        73:
            _3912 <= _3357;
        74:
            _3912 <= _3360;
        75:
            _3912 <= _3363;
        76:
            _3912 <= _3366;
        77:
            _3912 <= _3369;
        78:
            _3912 <= _3372;
        79:
            _3912 <= _3375;
        80:
            _3912 <= _3378;
        81:
            _3912 <= _3381;
        82:
            _3912 <= _3384;
        83:
            _3912 <= _3387;
        84:
            _3912 <= _3390;
        85:
            _3912 <= _3393;
        86:
            _3912 <= _3396;
        87:
            _3912 <= _3399;
        88:
            _3912 <= _3402;
        89:
            _3912 <= _3405;
        90:
            _3912 <= _3408;
        91:
            _3912 <= _3411;
        92:
            _3912 <= _3414;
        93:
            _3912 <= _3417;
        94:
            _3912 <= _3420;
        95:
            _3912 <= _3423;
        96:
            _3912 <= _3426;
        97:
            _3912 <= _3429;
        98:
            _3912 <= _3432;
        99:
            _3912 <= _3435;
        100:
            _3912 <= _3438;
        101:
            _3912 <= _3441;
        102:
            _3912 <= _3444;
        103:
            _3912 <= _3447;
        104:
            _3912 <= _3450;
        105:
            _3912 <= _3453;
        106:
            _3912 <= _3456;
        107:
            _3912 <= _3459;
        108:
            _3912 <= _3462;
        109:
            _3912 <= _3465;
        110:
            _3912 <= _3468;
        111:
            _3912 <= _3471;
        112:
            _3912 <= _3474;
        113:
            _3912 <= _3477;
        114:
            _3912 <= _3480;
        115:
            _3912 <= _3483;
        116:
            _3912 <= _3486;
        117:
            _3912 <= _3489;
        118:
            _3912 <= _3492;
        119:
            _3912 <= _3495;
        120:
            _3912 <= _3498;
        121:
            _3912 <= _3501;
        122:
            _3912 <= _3504;
        123:
            _3912 <= _3507;
        124:
            _3912 <= _3510;
        125:
            _3912 <= _3513;
        126:
            _3912 <= _3516;
        127:
            _3912 <= _3519;
        128:
            _3912 <= _3522;
        129:
            _3912 <= _3525;
        130:
            _3912 <= _3528;
        131:
            _3912 <= _3531;
        132:
            _3912 <= _3534;
        133:
            _3912 <= _3537;
        134:
            _3912 <= _3540;
        135:
            _3912 <= _3543;
        136:
            _3912 <= _3546;
        137:
            _3912 <= _3549;
        138:
            _3912 <= _3552;
        139:
            _3912 <= _3555;
        140:
            _3912 <= _3558;
        141:
            _3912 <= _3561;
        142:
            _3912 <= _3564;
        143:
            _3912 <= _3567;
        144:
            _3912 <= _3570;
        145:
            _3912 <= _3573;
        146:
            _3912 <= _3576;
        147:
            _3912 <= _3579;
        148:
            _3912 <= _3582;
        149:
            _3912 <= _3585;
        150:
            _3912 <= _3588;
        151:
            _3912 <= _3591;
        152:
            _3912 <= _3594;
        153:
            _3912 <= _3597;
        154:
            _3912 <= _3600;
        155:
            _3912 <= _3603;
        156:
            _3912 <= _3606;
        157:
            _3912 <= _3609;
        158:
            _3912 <= _3612;
        159:
            _3912 <= _3615;
        160:
            _3912 <= _3618;
        161:
            _3912 <= _3621;
        162:
            _3912 <= _3624;
        163:
            _3912 <= _3627;
        164:
            _3912 <= _3630;
        165:
            _3912 <= _3633;
        166:
            _3912 <= _3636;
        167:
            _3912 <= _3639;
        168:
            _3912 <= _3642;
        169:
            _3912 <= _3645;
        170:
            _3912 <= _3648;
        171:
            _3912 <= _3651;
        172:
            _3912 <= _3654;
        173:
            _3912 <= _3657;
        174:
            _3912 <= _3660;
        175:
            _3912 <= _3663;
        176:
            _3912 <= _3666;
        177:
            _3912 <= _3669;
        178:
            _3912 <= _3672;
        179:
            _3912 <= _3675;
        180:
            _3912 <= _3678;
        181:
            _3912 <= _3681;
        182:
            _3912 <= _3684;
        183:
            _3912 <= _3687;
        184:
            _3912 <= _3690;
        185:
            _3912 <= _3693;
        186:
            _3912 <= _3696;
        187:
            _3912 <= _3699;
        188:
            _3912 <= _3702;
        189:
            _3912 <= _3705;
        190:
            _3912 <= _3708;
        191:
            _3912 <= _3711;
        192:
            _3912 <= _3714;
        193:
            _3912 <= _3717;
        194:
            _3912 <= _3720;
        195:
            _3912 <= _3723;
        196:
            _3912 <= _3726;
        197:
            _3912 <= _3729;
        198:
            _3912 <= _3732;
        199:
            _3912 <= _3735;
        200:
            _3912 <= _3738;
        201:
            _3912 <= _3741;
        202:
            _3912 <= _3744;
        203:
            _3912 <= _3747;
        204:
            _3912 <= _3750;
        205:
            _3912 <= _3753;
        206:
            _3912 <= _3756;
        207:
            _3912 <= _3759;
        208:
            _3912 <= _3762;
        209:
            _3912 <= _3765;
        210:
            _3912 <= _3768;
        211:
            _3912 <= _3771;
        212:
            _3912 <= _3774;
        213:
            _3912 <= _3777;
        214:
            _3912 <= _3780;
        215:
            _3912 <= _3783;
        216:
            _3912 <= _3786;
        217:
            _3912 <= _3789;
        218:
            _3912 <= _3792;
        219:
            _3912 <= _3795;
        220:
            _3912 <= _3798;
        221:
            _3912 <= _3801;
        222:
            _3912 <= _3804;
        223:
            _3912 <= _3807;
        224:
            _3912 <= _3810;
        225:
            _3912 <= _3813;
        226:
            _3912 <= _3816;
        227:
            _3912 <= _3819;
        228:
            _3912 <= _3822;
        229:
            _3912 <= _3825;
        230:
            _3912 <= _3828;
        231:
            _3912 <= _3831;
        232:
            _3912 <= _3834;
        233:
            _3912 <= _3837;
        234:
            _3912 <= _3840;
        235:
            _3912 <= _3843;
        236:
            _3912 <= _3846;
        237:
            _3912 <= _3849;
        238:
            _3912 <= _3852;
        239:
            _3912 <= _3855;
        240:
            _3912 <= _3858;
        241:
            _3912 <= _3861;
        242:
            _3912 <= _3864;
        243:
            _3912 <= _3867;
        244:
            _3912 <= _3870;
        245:
            _3912 <= _3873;
        246:
            _3912 <= _3876;
        247:
            _3912 <= _3879;
        248:
            _3912 <= _3882;
        249:
            _3912 <= _3885;
        250:
            _3912 <= _3888;
        251:
            _3912 <= _3891;
        252:
            _3912 <= _3894;
        253:
            _3912 <= _3897;
        254:
            _3912 <= _3900;
        default:
            _3912 <= _3903;
        endcase
    end
    always @* begin
        case (_3912)
        0:
            _3913 <= _3138;
        1:
            _3913 <= _3141;
        2:
            _3913 <= _3144;
        3:
            _3913 <= _3147;
        4:
            _3913 <= _3150;
        5:
            _3913 <= _3153;
        6:
            _3913 <= _3156;
        7:
            _3913 <= _3159;
        8:
            _3913 <= _3162;
        9:
            _3913 <= _3165;
        10:
            _3913 <= _3168;
        11:
            _3913 <= _3171;
        12:
            _3913 <= _3174;
        13:
            _3913 <= _3177;
        14:
            _3913 <= _3180;
        15:
            _3913 <= _3183;
        16:
            _3913 <= _3186;
        17:
            _3913 <= _3189;
        18:
            _3913 <= _3192;
        19:
            _3913 <= _3195;
        20:
            _3913 <= _3198;
        21:
            _3913 <= _3201;
        22:
            _3913 <= _3204;
        23:
            _3913 <= _3207;
        24:
            _3913 <= _3210;
        25:
            _3913 <= _3213;
        26:
            _3913 <= _3216;
        27:
            _3913 <= _3219;
        28:
            _3913 <= _3222;
        29:
            _3913 <= _3225;
        30:
            _3913 <= _3228;
        31:
            _3913 <= _3231;
        32:
            _3913 <= _3234;
        33:
            _3913 <= _3237;
        34:
            _3913 <= _3240;
        35:
            _3913 <= _3243;
        36:
            _3913 <= _3246;
        37:
            _3913 <= _3249;
        38:
            _3913 <= _3252;
        39:
            _3913 <= _3255;
        40:
            _3913 <= _3258;
        41:
            _3913 <= _3261;
        42:
            _3913 <= _3264;
        43:
            _3913 <= _3267;
        44:
            _3913 <= _3270;
        45:
            _3913 <= _3273;
        46:
            _3913 <= _3276;
        47:
            _3913 <= _3279;
        48:
            _3913 <= _3282;
        49:
            _3913 <= _3285;
        50:
            _3913 <= _3288;
        51:
            _3913 <= _3291;
        52:
            _3913 <= _3294;
        53:
            _3913 <= _3297;
        54:
            _3913 <= _3300;
        55:
            _3913 <= _3303;
        56:
            _3913 <= _3306;
        57:
            _3913 <= _3309;
        58:
            _3913 <= _3312;
        59:
            _3913 <= _3315;
        60:
            _3913 <= _3318;
        61:
            _3913 <= _3321;
        62:
            _3913 <= _3324;
        63:
            _3913 <= _3327;
        64:
            _3913 <= _3330;
        65:
            _3913 <= _3333;
        66:
            _3913 <= _3336;
        67:
            _3913 <= _3339;
        68:
            _3913 <= _3342;
        69:
            _3913 <= _3345;
        70:
            _3913 <= _3348;
        71:
            _3913 <= _3351;
        72:
            _3913 <= _3354;
        73:
            _3913 <= _3357;
        74:
            _3913 <= _3360;
        75:
            _3913 <= _3363;
        76:
            _3913 <= _3366;
        77:
            _3913 <= _3369;
        78:
            _3913 <= _3372;
        79:
            _3913 <= _3375;
        80:
            _3913 <= _3378;
        81:
            _3913 <= _3381;
        82:
            _3913 <= _3384;
        83:
            _3913 <= _3387;
        84:
            _3913 <= _3390;
        85:
            _3913 <= _3393;
        86:
            _3913 <= _3396;
        87:
            _3913 <= _3399;
        88:
            _3913 <= _3402;
        89:
            _3913 <= _3405;
        90:
            _3913 <= _3408;
        91:
            _3913 <= _3411;
        92:
            _3913 <= _3414;
        93:
            _3913 <= _3417;
        94:
            _3913 <= _3420;
        95:
            _3913 <= _3423;
        96:
            _3913 <= _3426;
        97:
            _3913 <= _3429;
        98:
            _3913 <= _3432;
        99:
            _3913 <= _3435;
        100:
            _3913 <= _3438;
        101:
            _3913 <= _3441;
        102:
            _3913 <= _3444;
        103:
            _3913 <= _3447;
        104:
            _3913 <= _3450;
        105:
            _3913 <= _3453;
        106:
            _3913 <= _3456;
        107:
            _3913 <= _3459;
        108:
            _3913 <= _3462;
        109:
            _3913 <= _3465;
        110:
            _3913 <= _3468;
        111:
            _3913 <= _3471;
        112:
            _3913 <= _3474;
        113:
            _3913 <= _3477;
        114:
            _3913 <= _3480;
        115:
            _3913 <= _3483;
        116:
            _3913 <= _3486;
        117:
            _3913 <= _3489;
        118:
            _3913 <= _3492;
        119:
            _3913 <= _3495;
        120:
            _3913 <= _3498;
        121:
            _3913 <= _3501;
        122:
            _3913 <= _3504;
        123:
            _3913 <= _3507;
        124:
            _3913 <= _3510;
        125:
            _3913 <= _3513;
        126:
            _3913 <= _3516;
        127:
            _3913 <= _3519;
        128:
            _3913 <= _3522;
        129:
            _3913 <= _3525;
        130:
            _3913 <= _3528;
        131:
            _3913 <= _3531;
        132:
            _3913 <= _3534;
        133:
            _3913 <= _3537;
        134:
            _3913 <= _3540;
        135:
            _3913 <= _3543;
        136:
            _3913 <= _3546;
        137:
            _3913 <= _3549;
        138:
            _3913 <= _3552;
        139:
            _3913 <= _3555;
        140:
            _3913 <= _3558;
        141:
            _3913 <= _3561;
        142:
            _3913 <= _3564;
        143:
            _3913 <= _3567;
        144:
            _3913 <= _3570;
        145:
            _3913 <= _3573;
        146:
            _3913 <= _3576;
        147:
            _3913 <= _3579;
        148:
            _3913 <= _3582;
        149:
            _3913 <= _3585;
        150:
            _3913 <= _3588;
        151:
            _3913 <= _3591;
        152:
            _3913 <= _3594;
        153:
            _3913 <= _3597;
        154:
            _3913 <= _3600;
        155:
            _3913 <= _3603;
        156:
            _3913 <= _3606;
        157:
            _3913 <= _3609;
        158:
            _3913 <= _3612;
        159:
            _3913 <= _3615;
        160:
            _3913 <= _3618;
        161:
            _3913 <= _3621;
        162:
            _3913 <= _3624;
        163:
            _3913 <= _3627;
        164:
            _3913 <= _3630;
        165:
            _3913 <= _3633;
        166:
            _3913 <= _3636;
        167:
            _3913 <= _3639;
        168:
            _3913 <= _3642;
        169:
            _3913 <= _3645;
        170:
            _3913 <= _3648;
        171:
            _3913 <= _3651;
        172:
            _3913 <= _3654;
        173:
            _3913 <= _3657;
        174:
            _3913 <= _3660;
        175:
            _3913 <= _3663;
        176:
            _3913 <= _3666;
        177:
            _3913 <= _3669;
        178:
            _3913 <= _3672;
        179:
            _3913 <= _3675;
        180:
            _3913 <= _3678;
        181:
            _3913 <= _3681;
        182:
            _3913 <= _3684;
        183:
            _3913 <= _3687;
        184:
            _3913 <= _3690;
        185:
            _3913 <= _3693;
        186:
            _3913 <= _3696;
        187:
            _3913 <= _3699;
        188:
            _3913 <= _3702;
        189:
            _3913 <= _3705;
        190:
            _3913 <= _3708;
        191:
            _3913 <= _3711;
        192:
            _3913 <= _3714;
        193:
            _3913 <= _3717;
        194:
            _3913 <= _3720;
        195:
            _3913 <= _3723;
        196:
            _3913 <= _3726;
        197:
            _3913 <= _3729;
        198:
            _3913 <= _3732;
        199:
            _3913 <= _3735;
        200:
            _3913 <= _3738;
        201:
            _3913 <= _3741;
        202:
            _3913 <= _3744;
        203:
            _3913 <= _3747;
        204:
            _3913 <= _3750;
        205:
            _3913 <= _3753;
        206:
            _3913 <= _3756;
        207:
            _3913 <= _3759;
        208:
            _3913 <= _3762;
        209:
            _3913 <= _3765;
        210:
            _3913 <= _3768;
        211:
            _3913 <= _3771;
        212:
            _3913 <= _3774;
        213:
            _3913 <= _3777;
        214:
            _3913 <= _3780;
        215:
            _3913 <= _3783;
        216:
            _3913 <= _3786;
        217:
            _3913 <= _3789;
        218:
            _3913 <= _3792;
        219:
            _3913 <= _3795;
        220:
            _3913 <= _3798;
        221:
            _3913 <= _3801;
        222:
            _3913 <= _3804;
        223:
            _3913 <= _3807;
        224:
            _3913 <= _3810;
        225:
            _3913 <= _3813;
        226:
            _3913 <= _3816;
        227:
            _3913 <= _3819;
        228:
            _3913 <= _3822;
        229:
            _3913 <= _3825;
        230:
            _3913 <= _3828;
        231:
            _3913 <= _3831;
        232:
            _3913 <= _3834;
        233:
            _3913 <= _3837;
        234:
            _3913 <= _3840;
        235:
            _3913 <= _3843;
        236:
            _3913 <= _3846;
        237:
            _3913 <= _3849;
        238:
            _3913 <= _3852;
        239:
            _3913 <= _3855;
        240:
            _3913 <= _3858;
        241:
            _3913 <= _3861;
        242:
            _3913 <= _3864;
        243:
            _3913 <= _3867;
        244:
            _3913 <= _3870;
        245:
            _3913 <= _3873;
        246:
            _3913 <= _3876;
        247:
            _3913 <= _3879;
        248:
            _3913 <= _3882;
        249:
            _3913 <= _3885;
        250:
            _3913 <= _3888;
        251:
            _3913 <= _3891;
        252:
            _3913 <= _3894;
        253:
            _3913 <= _3897;
        254:
            _3913 <= _3900;
        default:
            _3913 <= _3903;
        endcase
    end
    always @* begin
        case (_3913)
        0:
            _3914 <= _3138;
        1:
            _3914 <= _3141;
        2:
            _3914 <= _3144;
        3:
            _3914 <= _3147;
        4:
            _3914 <= _3150;
        5:
            _3914 <= _3153;
        6:
            _3914 <= _3156;
        7:
            _3914 <= _3159;
        8:
            _3914 <= _3162;
        9:
            _3914 <= _3165;
        10:
            _3914 <= _3168;
        11:
            _3914 <= _3171;
        12:
            _3914 <= _3174;
        13:
            _3914 <= _3177;
        14:
            _3914 <= _3180;
        15:
            _3914 <= _3183;
        16:
            _3914 <= _3186;
        17:
            _3914 <= _3189;
        18:
            _3914 <= _3192;
        19:
            _3914 <= _3195;
        20:
            _3914 <= _3198;
        21:
            _3914 <= _3201;
        22:
            _3914 <= _3204;
        23:
            _3914 <= _3207;
        24:
            _3914 <= _3210;
        25:
            _3914 <= _3213;
        26:
            _3914 <= _3216;
        27:
            _3914 <= _3219;
        28:
            _3914 <= _3222;
        29:
            _3914 <= _3225;
        30:
            _3914 <= _3228;
        31:
            _3914 <= _3231;
        32:
            _3914 <= _3234;
        33:
            _3914 <= _3237;
        34:
            _3914 <= _3240;
        35:
            _3914 <= _3243;
        36:
            _3914 <= _3246;
        37:
            _3914 <= _3249;
        38:
            _3914 <= _3252;
        39:
            _3914 <= _3255;
        40:
            _3914 <= _3258;
        41:
            _3914 <= _3261;
        42:
            _3914 <= _3264;
        43:
            _3914 <= _3267;
        44:
            _3914 <= _3270;
        45:
            _3914 <= _3273;
        46:
            _3914 <= _3276;
        47:
            _3914 <= _3279;
        48:
            _3914 <= _3282;
        49:
            _3914 <= _3285;
        50:
            _3914 <= _3288;
        51:
            _3914 <= _3291;
        52:
            _3914 <= _3294;
        53:
            _3914 <= _3297;
        54:
            _3914 <= _3300;
        55:
            _3914 <= _3303;
        56:
            _3914 <= _3306;
        57:
            _3914 <= _3309;
        58:
            _3914 <= _3312;
        59:
            _3914 <= _3315;
        60:
            _3914 <= _3318;
        61:
            _3914 <= _3321;
        62:
            _3914 <= _3324;
        63:
            _3914 <= _3327;
        64:
            _3914 <= _3330;
        65:
            _3914 <= _3333;
        66:
            _3914 <= _3336;
        67:
            _3914 <= _3339;
        68:
            _3914 <= _3342;
        69:
            _3914 <= _3345;
        70:
            _3914 <= _3348;
        71:
            _3914 <= _3351;
        72:
            _3914 <= _3354;
        73:
            _3914 <= _3357;
        74:
            _3914 <= _3360;
        75:
            _3914 <= _3363;
        76:
            _3914 <= _3366;
        77:
            _3914 <= _3369;
        78:
            _3914 <= _3372;
        79:
            _3914 <= _3375;
        80:
            _3914 <= _3378;
        81:
            _3914 <= _3381;
        82:
            _3914 <= _3384;
        83:
            _3914 <= _3387;
        84:
            _3914 <= _3390;
        85:
            _3914 <= _3393;
        86:
            _3914 <= _3396;
        87:
            _3914 <= _3399;
        88:
            _3914 <= _3402;
        89:
            _3914 <= _3405;
        90:
            _3914 <= _3408;
        91:
            _3914 <= _3411;
        92:
            _3914 <= _3414;
        93:
            _3914 <= _3417;
        94:
            _3914 <= _3420;
        95:
            _3914 <= _3423;
        96:
            _3914 <= _3426;
        97:
            _3914 <= _3429;
        98:
            _3914 <= _3432;
        99:
            _3914 <= _3435;
        100:
            _3914 <= _3438;
        101:
            _3914 <= _3441;
        102:
            _3914 <= _3444;
        103:
            _3914 <= _3447;
        104:
            _3914 <= _3450;
        105:
            _3914 <= _3453;
        106:
            _3914 <= _3456;
        107:
            _3914 <= _3459;
        108:
            _3914 <= _3462;
        109:
            _3914 <= _3465;
        110:
            _3914 <= _3468;
        111:
            _3914 <= _3471;
        112:
            _3914 <= _3474;
        113:
            _3914 <= _3477;
        114:
            _3914 <= _3480;
        115:
            _3914 <= _3483;
        116:
            _3914 <= _3486;
        117:
            _3914 <= _3489;
        118:
            _3914 <= _3492;
        119:
            _3914 <= _3495;
        120:
            _3914 <= _3498;
        121:
            _3914 <= _3501;
        122:
            _3914 <= _3504;
        123:
            _3914 <= _3507;
        124:
            _3914 <= _3510;
        125:
            _3914 <= _3513;
        126:
            _3914 <= _3516;
        127:
            _3914 <= _3519;
        128:
            _3914 <= _3522;
        129:
            _3914 <= _3525;
        130:
            _3914 <= _3528;
        131:
            _3914 <= _3531;
        132:
            _3914 <= _3534;
        133:
            _3914 <= _3537;
        134:
            _3914 <= _3540;
        135:
            _3914 <= _3543;
        136:
            _3914 <= _3546;
        137:
            _3914 <= _3549;
        138:
            _3914 <= _3552;
        139:
            _3914 <= _3555;
        140:
            _3914 <= _3558;
        141:
            _3914 <= _3561;
        142:
            _3914 <= _3564;
        143:
            _3914 <= _3567;
        144:
            _3914 <= _3570;
        145:
            _3914 <= _3573;
        146:
            _3914 <= _3576;
        147:
            _3914 <= _3579;
        148:
            _3914 <= _3582;
        149:
            _3914 <= _3585;
        150:
            _3914 <= _3588;
        151:
            _3914 <= _3591;
        152:
            _3914 <= _3594;
        153:
            _3914 <= _3597;
        154:
            _3914 <= _3600;
        155:
            _3914 <= _3603;
        156:
            _3914 <= _3606;
        157:
            _3914 <= _3609;
        158:
            _3914 <= _3612;
        159:
            _3914 <= _3615;
        160:
            _3914 <= _3618;
        161:
            _3914 <= _3621;
        162:
            _3914 <= _3624;
        163:
            _3914 <= _3627;
        164:
            _3914 <= _3630;
        165:
            _3914 <= _3633;
        166:
            _3914 <= _3636;
        167:
            _3914 <= _3639;
        168:
            _3914 <= _3642;
        169:
            _3914 <= _3645;
        170:
            _3914 <= _3648;
        171:
            _3914 <= _3651;
        172:
            _3914 <= _3654;
        173:
            _3914 <= _3657;
        174:
            _3914 <= _3660;
        175:
            _3914 <= _3663;
        176:
            _3914 <= _3666;
        177:
            _3914 <= _3669;
        178:
            _3914 <= _3672;
        179:
            _3914 <= _3675;
        180:
            _3914 <= _3678;
        181:
            _3914 <= _3681;
        182:
            _3914 <= _3684;
        183:
            _3914 <= _3687;
        184:
            _3914 <= _3690;
        185:
            _3914 <= _3693;
        186:
            _3914 <= _3696;
        187:
            _3914 <= _3699;
        188:
            _3914 <= _3702;
        189:
            _3914 <= _3705;
        190:
            _3914 <= _3708;
        191:
            _3914 <= _3711;
        192:
            _3914 <= _3714;
        193:
            _3914 <= _3717;
        194:
            _3914 <= _3720;
        195:
            _3914 <= _3723;
        196:
            _3914 <= _3726;
        197:
            _3914 <= _3729;
        198:
            _3914 <= _3732;
        199:
            _3914 <= _3735;
        200:
            _3914 <= _3738;
        201:
            _3914 <= _3741;
        202:
            _3914 <= _3744;
        203:
            _3914 <= _3747;
        204:
            _3914 <= _3750;
        205:
            _3914 <= _3753;
        206:
            _3914 <= _3756;
        207:
            _3914 <= _3759;
        208:
            _3914 <= _3762;
        209:
            _3914 <= _3765;
        210:
            _3914 <= _3768;
        211:
            _3914 <= _3771;
        212:
            _3914 <= _3774;
        213:
            _3914 <= _3777;
        214:
            _3914 <= _3780;
        215:
            _3914 <= _3783;
        216:
            _3914 <= _3786;
        217:
            _3914 <= _3789;
        218:
            _3914 <= _3792;
        219:
            _3914 <= _3795;
        220:
            _3914 <= _3798;
        221:
            _3914 <= _3801;
        222:
            _3914 <= _3804;
        223:
            _3914 <= _3807;
        224:
            _3914 <= _3810;
        225:
            _3914 <= _3813;
        226:
            _3914 <= _3816;
        227:
            _3914 <= _3819;
        228:
            _3914 <= _3822;
        229:
            _3914 <= _3825;
        230:
            _3914 <= _3828;
        231:
            _3914 <= _3831;
        232:
            _3914 <= _3834;
        233:
            _3914 <= _3837;
        234:
            _3914 <= _3840;
        235:
            _3914 <= _3843;
        236:
            _3914 <= _3846;
        237:
            _3914 <= _3849;
        238:
            _3914 <= _3852;
        239:
            _3914 <= _3855;
        240:
            _3914 <= _3858;
        241:
            _3914 <= _3861;
        242:
            _3914 <= _3864;
        243:
            _3914 <= _3867;
        244:
            _3914 <= _3870;
        245:
            _3914 <= _3873;
        246:
            _3914 <= _3876;
        247:
            _3914 <= _3879;
        248:
            _3914 <= _3882;
        249:
            _3914 <= _3885;
        250:
            _3914 <= _3888;
        251:
            _3914 <= _3891;
        252:
            _3914 <= _3894;
        253:
            _3914 <= _3897;
        254:
            _3914 <= _3900;
        default:
            _3914 <= _3903;
        endcase
    end
    always @* begin
        case (_3914)
        0:
            _3915 <= _3138;
        1:
            _3915 <= _3141;
        2:
            _3915 <= _3144;
        3:
            _3915 <= _3147;
        4:
            _3915 <= _3150;
        5:
            _3915 <= _3153;
        6:
            _3915 <= _3156;
        7:
            _3915 <= _3159;
        8:
            _3915 <= _3162;
        9:
            _3915 <= _3165;
        10:
            _3915 <= _3168;
        11:
            _3915 <= _3171;
        12:
            _3915 <= _3174;
        13:
            _3915 <= _3177;
        14:
            _3915 <= _3180;
        15:
            _3915 <= _3183;
        16:
            _3915 <= _3186;
        17:
            _3915 <= _3189;
        18:
            _3915 <= _3192;
        19:
            _3915 <= _3195;
        20:
            _3915 <= _3198;
        21:
            _3915 <= _3201;
        22:
            _3915 <= _3204;
        23:
            _3915 <= _3207;
        24:
            _3915 <= _3210;
        25:
            _3915 <= _3213;
        26:
            _3915 <= _3216;
        27:
            _3915 <= _3219;
        28:
            _3915 <= _3222;
        29:
            _3915 <= _3225;
        30:
            _3915 <= _3228;
        31:
            _3915 <= _3231;
        32:
            _3915 <= _3234;
        33:
            _3915 <= _3237;
        34:
            _3915 <= _3240;
        35:
            _3915 <= _3243;
        36:
            _3915 <= _3246;
        37:
            _3915 <= _3249;
        38:
            _3915 <= _3252;
        39:
            _3915 <= _3255;
        40:
            _3915 <= _3258;
        41:
            _3915 <= _3261;
        42:
            _3915 <= _3264;
        43:
            _3915 <= _3267;
        44:
            _3915 <= _3270;
        45:
            _3915 <= _3273;
        46:
            _3915 <= _3276;
        47:
            _3915 <= _3279;
        48:
            _3915 <= _3282;
        49:
            _3915 <= _3285;
        50:
            _3915 <= _3288;
        51:
            _3915 <= _3291;
        52:
            _3915 <= _3294;
        53:
            _3915 <= _3297;
        54:
            _3915 <= _3300;
        55:
            _3915 <= _3303;
        56:
            _3915 <= _3306;
        57:
            _3915 <= _3309;
        58:
            _3915 <= _3312;
        59:
            _3915 <= _3315;
        60:
            _3915 <= _3318;
        61:
            _3915 <= _3321;
        62:
            _3915 <= _3324;
        63:
            _3915 <= _3327;
        64:
            _3915 <= _3330;
        65:
            _3915 <= _3333;
        66:
            _3915 <= _3336;
        67:
            _3915 <= _3339;
        68:
            _3915 <= _3342;
        69:
            _3915 <= _3345;
        70:
            _3915 <= _3348;
        71:
            _3915 <= _3351;
        72:
            _3915 <= _3354;
        73:
            _3915 <= _3357;
        74:
            _3915 <= _3360;
        75:
            _3915 <= _3363;
        76:
            _3915 <= _3366;
        77:
            _3915 <= _3369;
        78:
            _3915 <= _3372;
        79:
            _3915 <= _3375;
        80:
            _3915 <= _3378;
        81:
            _3915 <= _3381;
        82:
            _3915 <= _3384;
        83:
            _3915 <= _3387;
        84:
            _3915 <= _3390;
        85:
            _3915 <= _3393;
        86:
            _3915 <= _3396;
        87:
            _3915 <= _3399;
        88:
            _3915 <= _3402;
        89:
            _3915 <= _3405;
        90:
            _3915 <= _3408;
        91:
            _3915 <= _3411;
        92:
            _3915 <= _3414;
        93:
            _3915 <= _3417;
        94:
            _3915 <= _3420;
        95:
            _3915 <= _3423;
        96:
            _3915 <= _3426;
        97:
            _3915 <= _3429;
        98:
            _3915 <= _3432;
        99:
            _3915 <= _3435;
        100:
            _3915 <= _3438;
        101:
            _3915 <= _3441;
        102:
            _3915 <= _3444;
        103:
            _3915 <= _3447;
        104:
            _3915 <= _3450;
        105:
            _3915 <= _3453;
        106:
            _3915 <= _3456;
        107:
            _3915 <= _3459;
        108:
            _3915 <= _3462;
        109:
            _3915 <= _3465;
        110:
            _3915 <= _3468;
        111:
            _3915 <= _3471;
        112:
            _3915 <= _3474;
        113:
            _3915 <= _3477;
        114:
            _3915 <= _3480;
        115:
            _3915 <= _3483;
        116:
            _3915 <= _3486;
        117:
            _3915 <= _3489;
        118:
            _3915 <= _3492;
        119:
            _3915 <= _3495;
        120:
            _3915 <= _3498;
        121:
            _3915 <= _3501;
        122:
            _3915 <= _3504;
        123:
            _3915 <= _3507;
        124:
            _3915 <= _3510;
        125:
            _3915 <= _3513;
        126:
            _3915 <= _3516;
        127:
            _3915 <= _3519;
        128:
            _3915 <= _3522;
        129:
            _3915 <= _3525;
        130:
            _3915 <= _3528;
        131:
            _3915 <= _3531;
        132:
            _3915 <= _3534;
        133:
            _3915 <= _3537;
        134:
            _3915 <= _3540;
        135:
            _3915 <= _3543;
        136:
            _3915 <= _3546;
        137:
            _3915 <= _3549;
        138:
            _3915 <= _3552;
        139:
            _3915 <= _3555;
        140:
            _3915 <= _3558;
        141:
            _3915 <= _3561;
        142:
            _3915 <= _3564;
        143:
            _3915 <= _3567;
        144:
            _3915 <= _3570;
        145:
            _3915 <= _3573;
        146:
            _3915 <= _3576;
        147:
            _3915 <= _3579;
        148:
            _3915 <= _3582;
        149:
            _3915 <= _3585;
        150:
            _3915 <= _3588;
        151:
            _3915 <= _3591;
        152:
            _3915 <= _3594;
        153:
            _3915 <= _3597;
        154:
            _3915 <= _3600;
        155:
            _3915 <= _3603;
        156:
            _3915 <= _3606;
        157:
            _3915 <= _3609;
        158:
            _3915 <= _3612;
        159:
            _3915 <= _3615;
        160:
            _3915 <= _3618;
        161:
            _3915 <= _3621;
        162:
            _3915 <= _3624;
        163:
            _3915 <= _3627;
        164:
            _3915 <= _3630;
        165:
            _3915 <= _3633;
        166:
            _3915 <= _3636;
        167:
            _3915 <= _3639;
        168:
            _3915 <= _3642;
        169:
            _3915 <= _3645;
        170:
            _3915 <= _3648;
        171:
            _3915 <= _3651;
        172:
            _3915 <= _3654;
        173:
            _3915 <= _3657;
        174:
            _3915 <= _3660;
        175:
            _3915 <= _3663;
        176:
            _3915 <= _3666;
        177:
            _3915 <= _3669;
        178:
            _3915 <= _3672;
        179:
            _3915 <= _3675;
        180:
            _3915 <= _3678;
        181:
            _3915 <= _3681;
        182:
            _3915 <= _3684;
        183:
            _3915 <= _3687;
        184:
            _3915 <= _3690;
        185:
            _3915 <= _3693;
        186:
            _3915 <= _3696;
        187:
            _3915 <= _3699;
        188:
            _3915 <= _3702;
        189:
            _3915 <= _3705;
        190:
            _3915 <= _3708;
        191:
            _3915 <= _3711;
        192:
            _3915 <= _3714;
        193:
            _3915 <= _3717;
        194:
            _3915 <= _3720;
        195:
            _3915 <= _3723;
        196:
            _3915 <= _3726;
        197:
            _3915 <= _3729;
        198:
            _3915 <= _3732;
        199:
            _3915 <= _3735;
        200:
            _3915 <= _3738;
        201:
            _3915 <= _3741;
        202:
            _3915 <= _3744;
        203:
            _3915 <= _3747;
        204:
            _3915 <= _3750;
        205:
            _3915 <= _3753;
        206:
            _3915 <= _3756;
        207:
            _3915 <= _3759;
        208:
            _3915 <= _3762;
        209:
            _3915 <= _3765;
        210:
            _3915 <= _3768;
        211:
            _3915 <= _3771;
        212:
            _3915 <= _3774;
        213:
            _3915 <= _3777;
        214:
            _3915 <= _3780;
        215:
            _3915 <= _3783;
        216:
            _3915 <= _3786;
        217:
            _3915 <= _3789;
        218:
            _3915 <= _3792;
        219:
            _3915 <= _3795;
        220:
            _3915 <= _3798;
        221:
            _3915 <= _3801;
        222:
            _3915 <= _3804;
        223:
            _3915 <= _3807;
        224:
            _3915 <= _3810;
        225:
            _3915 <= _3813;
        226:
            _3915 <= _3816;
        227:
            _3915 <= _3819;
        228:
            _3915 <= _3822;
        229:
            _3915 <= _3825;
        230:
            _3915 <= _3828;
        231:
            _3915 <= _3831;
        232:
            _3915 <= _3834;
        233:
            _3915 <= _3837;
        234:
            _3915 <= _3840;
        235:
            _3915 <= _3843;
        236:
            _3915 <= _3846;
        237:
            _3915 <= _3849;
        238:
            _3915 <= _3852;
        239:
            _3915 <= _3855;
        240:
            _3915 <= _3858;
        241:
            _3915 <= _3861;
        242:
            _3915 <= _3864;
        243:
            _3915 <= _3867;
        244:
            _3915 <= _3870;
        245:
            _3915 <= _3873;
        246:
            _3915 <= _3876;
        247:
            _3915 <= _3879;
        248:
            _3915 <= _3882;
        249:
            _3915 <= _3885;
        250:
            _3915 <= _3888;
        251:
            _3915 <= _3891;
        252:
            _3915 <= _3894;
        253:
            _3915 <= _3897;
        254:
            _3915 <= _3900;
        default:
            _3915 <= _3903;
        endcase
    end
    always @* begin
        case (_3915)
        0:
            _3916 <= _3138;
        1:
            _3916 <= _3141;
        2:
            _3916 <= _3144;
        3:
            _3916 <= _3147;
        4:
            _3916 <= _3150;
        5:
            _3916 <= _3153;
        6:
            _3916 <= _3156;
        7:
            _3916 <= _3159;
        8:
            _3916 <= _3162;
        9:
            _3916 <= _3165;
        10:
            _3916 <= _3168;
        11:
            _3916 <= _3171;
        12:
            _3916 <= _3174;
        13:
            _3916 <= _3177;
        14:
            _3916 <= _3180;
        15:
            _3916 <= _3183;
        16:
            _3916 <= _3186;
        17:
            _3916 <= _3189;
        18:
            _3916 <= _3192;
        19:
            _3916 <= _3195;
        20:
            _3916 <= _3198;
        21:
            _3916 <= _3201;
        22:
            _3916 <= _3204;
        23:
            _3916 <= _3207;
        24:
            _3916 <= _3210;
        25:
            _3916 <= _3213;
        26:
            _3916 <= _3216;
        27:
            _3916 <= _3219;
        28:
            _3916 <= _3222;
        29:
            _3916 <= _3225;
        30:
            _3916 <= _3228;
        31:
            _3916 <= _3231;
        32:
            _3916 <= _3234;
        33:
            _3916 <= _3237;
        34:
            _3916 <= _3240;
        35:
            _3916 <= _3243;
        36:
            _3916 <= _3246;
        37:
            _3916 <= _3249;
        38:
            _3916 <= _3252;
        39:
            _3916 <= _3255;
        40:
            _3916 <= _3258;
        41:
            _3916 <= _3261;
        42:
            _3916 <= _3264;
        43:
            _3916 <= _3267;
        44:
            _3916 <= _3270;
        45:
            _3916 <= _3273;
        46:
            _3916 <= _3276;
        47:
            _3916 <= _3279;
        48:
            _3916 <= _3282;
        49:
            _3916 <= _3285;
        50:
            _3916 <= _3288;
        51:
            _3916 <= _3291;
        52:
            _3916 <= _3294;
        53:
            _3916 <= _3297;
        54:
            _3916 <= _3300;
        55:
            _3916 <= _3303;
        56:
            _3916 <= _3306;
        57:
            _3916 <= _3309;
        58:
            _3916 <= _3312;
        59:
            _3916 <= _3315;
        60:
            _3916 <= _3318;
        61:
            _3916 <= _3321;
        62:
            _3916 <= _3324;
        63:
            _3916 <= _3327;
        64:
            _3916 <= _3330;
        65:
            _3916 <= _3333;
        66:
            _3916 <= _3336;
        67:
            _3916 <= _3339;
        68:
            _3916 <= _3342;
        69:
            _3916 <= _3345;
        70:
            _3916 <= _3348;
        71:
            _3916 <= _3351;
        72:
            _3916 <= _3354;
        73:
            _3916 <= _3357;
        74:
            _3916 <= _3360;
        75:
            _3916 <= _3363;
        76:
            _3916 <= _3366;
        77:
            _3916 <= _3369;
        78:
            _3916 <= _3372;
        79:
            _3916 <= _3375;
        80:
            _3916 <= _3378;
        81:
            _3916 <= _3381;
        82:
            _3916 <= _3384;
        83:
            _3916 <= _3387;
        84:
            _3916 <= _3390;
        85:
            _3916 <= _3393;
        86:
            _3916 <= _3396;
        87:
            _3916 <= _3399;
        88:
            _3916 <= _3402;
        89:
            _3916 <= _3405;
        90:
            _3916 <= _3408;
        91:
            _3916 <= _3411;
        92:
            _3916 <= _3414;
        93:
            _3916 <= _3417;
        94:
            _3916 <= _3420;
        95:
            _3916 <= _3423;
        96:
            _3916 <= _3426;
        97:
            _3916 <= _3429;
        98:
            _3916 <= _3432;
        99:
            _3916 <= _3435;
        100:
            _3916 <= _3438;
        101:
            _3916 <= _3441;
        102:
            _3916 <= _3444;
        103:
            _3916 <= _3447;
        104:
            _3916 <= _3450;
        105:
            _3916 <= _3453;
        106:
            _3916 <= _3456;
        107:
            _3916 <= _3459;
        108:
            _3916 <= _3462;
        109:
            _3916 <= _3465;
        110:
            _3916 <= _3468;
        111:
            _3916 <= _3471;
        112:
            _3916 <= _3474;
        113:
            _3916 <= _3477;
        114:
            _3916 <= _3480;
        115:
            _3916 <= _3483;
        116:
            _3916 <= _3486;
        117:
            _3916 <= _3489;
        118:
            _3916 <= _3492;
        119:
            _3916 <= _3495;
        120:
            _3916 <= _3498;
        121:
            _3916 <= _3501;
        122:
            _3916 <= _3504;
        123:
            _3916 <= _3507;
        124:
            _3916 <= _3510;
        125:
            _3916 <= _3513;
        126:
            _3916 <= _3516;
        127:
            _3916 <= _3519;
        128:
            _3916 <= _3522;
        129:
            _3916 <= _3525;
        130:
            _3916 <= _3528;
        131:
            _3916 <= _3531;
        132:
            _3916 <= _3534;
        133:
            _3916 <= _3537;
        134:
            _3916 <= _3540;
        135:
            _3916 <= _3543;
        136:
            _3916 <= _3546;
        137:
            _3916 <= _3549;
        138:
            _3916 <= _3552;
        139:
            _3916 <= _3555;
        140:
            _3916 <= _3558;
        141:
            _3916 <= _3561;
        142:
            _3916 <= _3564;
        143:
            _3916 <= _3567;
        144:
            _3916 <= _3570;
        145:
            _3916 <= _3573;
        146:
            _3916 <= _3576;
        147:
            _3916 <= _3579;
        148:
            _3916 <= _3582;
        149:
            _3916 <= _3585;
        150:
            _3916 <= _3588;
        151:
            _3916 <= _3591;
        152:
            _3916 <= _3594;
        153:
            _3916 <= _3597;
        154:
            _3916 <= _3600;
        155:
            _3916 <= _3603;
        156:
            _3916 <= _3606;
        157:
            _3916 <= _3609;
        158:
            _3916 <= _3612;
        159:
            _3916 <= _3615;
        160:
            _3916 <= _3618;
        161:
            _3916 <= _3621;
        162:
            _3916 <= _3624;
        163:
            _3916 <= _3627;
        164:
            _3916 <= _3630;
        165:
            _3916 <= _3633;
        166:
            _3916 <= _3636;
        167:
            _3916 <= _3639;
        168:
            _3916 <= _3642;
        169:
            _3916 <= _3645;
        170:
            _3916 <= _3648;
        171:
            _3916 <= _3651;
        172:
            _3916 <= _3654;
        173:
            _3916 <= _3657;
        174:
            _3916 <= _3660;
        175:
            _3916 <= _3663;
        176:
            _3916 <= _3666;
        177:
            _3916 <= _3669;
        178:
            _3916 <= _3672;
        179:
            _3916 <= _3675;
        180:
            _3916 <= _3678;
        181:
            _3916 <= _3681;
        182:
            _3916 <= _3684;
        183:
            _3916 <= _3687;
        184:
            _3916 <= _3690;
        185:
            _3916 <= _3693;
        186:
            _3916 <= _3696;
        187:
            _3916 <= _3699;
        188:
            _3916 <= _3702;
        189:
            _3916 <= _3705;
        190:
            _3916 <= _3708;
        191:
            _3916 <= _3711;
        192:
            _3916 <= _3714;
        193:
            _3916 <= _3717;
        194:
            _3916 <= _3720;
        195:
            _3916 <= _3723;
        196:
            _3916 <= _3726;
        197:
            _3916 <= _3729;
        198:
            _3916 <= _3732;
        199:
            _3916 <= _3735;
        200:
            _3916 <= _3738;
        201:
            _3916 <= _3741;
        202:
            _3916 <= _3744;
        203:
            _3916 <= _3747;
        204:
            _3916 <= _3750;
        205:
            _3916 <= _3753;
        206:
            _3916 <= _3756;
        207:
            _3916 <= _3759;
        208:
            _3916 <= _3762;
        209:
            _3916 <= _3765;
        210:
            _3916 <= _3768;
        211:
            _3916 <= _3771;
        212:
            _3916 <= _3774;
        213:
            _3916 <= _3777;
        214:
            _3916 <= _3780;
        215:
            _3916 <= _3783;
        216:
            _3916 <= _3786;
        217:
            _3916 <= _3789;
        218:
            _3916 <= _3792;
        219:
            _3916 <= _3795;
        220:
            _3916 <= _3798;
        221:
            _3916 <= _3801;
        222:
            _3916 <= _3804;
        223:
            _3916 <= _3807;
        224:
            _3916 <= _3810;
        225:
            _3916 <= _3813;
        226:
            _3916 <= _3816;
        227:
            _3916 <= _3819;
        228:
            _3916 <= _3822;
        229:
            _3916 <= _3825;
        230:
            _3916 <= _3828;
        231:
            _3916 <= _3831;
        232:
            _3916 <= _3834;
        233:
            _3916 <= _3837;
        234:
            _3916 <= _3840;
        235:
            _3916 <= _3843;
        236:
            _3916 <= _3846;
        237:
            _3916 <= _3849;
        238:
            _3916 <= _3852;
        239:
            _3916 <= _3855;
        240:
            _3916 <= _3858;
        241:
            _3916 <= _3861;
        242:
            _3916 <= _3864;
        243:
            _3916 <= _3867;
        244:
            _3916 <= _3870;
        245:
            _3916 <= _3873;
        246:
            _3916 <= _3876;
        247:
            _3916 <= _3879;
        248:
            _3916 <= _3882;
        249:
            _3916 <= _3885;
        250:
            _3916 <= _3888;
        251:
            _3916 <= _3891;
        252:
            _3916 <= _3894;
        253:
            _3916 <= _3897;
        254:
            _3916 <= _3900;
        default:
            _3916 <= _3903;
        endcase
    end
    always @* begin
        case (_3916)
        0:
            _3917 <= _3138;
        1:
            _3917 <= _3141;
        2:
            _3917 <= _3144;
        3:
            _3917 <= _3147;
        4:
            _3917 <= _3150;
        5:
            _3917 <= _3153;
        6:
            _3917 <= _3156;
        7:
            _3917 <= _3159;
        8:
            _3917 <= _3162;
        9:
            _3917 <= _3165;
        10:
            _3917 <= _3168;
        11:
            _3917 <= _3171;
        12:
            _3917 <= _3174;
        13:
            _3917 <= _3177;
        14:
            _3917 <= _3180;
        15:
            _3917 <= _3183;
        16:
            _3917 <= _3186;
        17:
            _3917 <= _3189;
        18:
            _3917 <= _3192;
        19:
            _3917 <= _3195;
        20:
            _3917 <= _3198;
        21:
            _3917 <= _3201;
        22:
            _3917 <= _3204;
        23:
            _3917 <= _3207;
        24:
            _3917 <= _3210;
        25:
            _3917 <= _3213;
        26:
            _3917 <= _3216;
        27:
            _3917 <= _3219;
        28:
            _3917 <= _3222;
        29:
            _3917 <= _3225;
        30:
            _3917 <= _3228;
        31:
            _3917 <= _3231;
        32:
            _3917 <= _3234;
        33:
            _3917 <= _3237;
        34:
            _3917 <= _3240;
        35:
            _3917 <= _3243;
        36:
            _3917 <= _3246;
        37:
            _3917 <= _3249;
        38:
            _3917 <= _3252;
        39:
            _3917 <= _3255;
        40:
            _3917 <= _3258;
        41:
            _3917 <= _3261;
        42:
            _3917 <= _3264;
        43:
            _3917 <= _3267;
        44:
            _3917 <= _3270;
        45:
            _3917 <= _3273;
        46:
            _3917 <= _3276;
        47:
            _3917 <= _3279;
        48:
            _3917 <= _3282;
        49:
            _3917 <= _3285;
        50:
            _3917 <= _3288;
        51:
            _3917 <= _3291;
        52:
            _3917 <= _3294;
        53:
            _3917 <= _3297;
        54:
            _3917 <= _3300;
        55:
            _3917 <= _3303;
        56:
            _3917 <= _3306;
        57:
            _3917 <= _3309;
        58:
            _3917 <= _3312;
        59:
            _3917 <= _3315;
        60:
            _3917 <= _3318;
        61:
            _3917 <= _3321;
        62:
            _3917 <= _3324;
        63:
            _3917 <= _3327;
        64:
            _3917 <= _3330;
        65:
            _3917 <= _3333;
        66:
            _3917 <= _3336;
        67:
            _3917 <= _3339;
        68:
            _3917 <= _3342;
        69:
            _3917 <= _3345;
        70:
            _3917 <= _3348;
        71:
            _3917 <= _3351;
        72:
            _3917 <= _3354;
        73:
            _3917 <= _3357;
        74:
            _3917 <= _3360;
        75:
            _3917 <= _3363;
        76:
            _3917 <= _3366;
        77:
            _3917 <= _3369;
        78:
            _3917 <= _3372;
        79:
            _3917 <= _3375;
        80:
            _3917 <= _3378;
        81:
            _3917 <= _3381;
        82:
            _3917 <= _3384;
        83:
            _3917 <= _3387;
        84:
            _3917 <= _3390;
        85:
            _3917 <= _3393;
        86:
            _3917 <= _3396;
        87:
            _3917 <= _3399;
        88:
            _3917 <= _3402;
        89:
            _3917 <= _3405;
        90:
            _3917 <= _3408;
        91:
            _3917 <= _3411;
        92:
            _3917 <= _3414;
        93:
            _3917 <= _3417;
        94:
            _3917 <= _3420;
        95:
            _3917 <= _3423;
        96:
            _3917 <= _3426;
        97:
            _3917 <= _3429;
        98:
            _3917 <= _3432;
        99:
            _3917 <= _3435;
        100:
            _3917 <= _3438;
        101:
            _3917 <= _3441;
        102:
            _3917 <= _3444;
        103:
            _3917 <= _3447;
        104:
            _3917 <= _3450;
        105:
            _3917 <= _3453;
        106:
            _3917 <= _3456;
        107:
            _3917 <= _3459;
        108:
            _3917 <= _3462;
        109:
            _3917 <= _3465;
        110:
            _3917 <= _3468;
        111:
            _3917 <= _3471;
        112:
            _3917 <= _3474;
        113:
            _3917 <= _3477;
        114:
            _3917 <= _3480;
        115:
            _3917 <= _3483;
        116:
            _3917 <= _3486;
        117:
            _3917 <= _3489;
        118:
            _3917 <= _3492;
        119:
            _3917 <= _3495;
        120:
            _3917 <= _3498;
        121:
            _3917 <= _3501;
        122:
            _3917 <= _3504;
        123:
            _3917 <= _3507;
        124:
            _3917 <= _3510;
        125:
            _3917 <= _3513;
        126:
            _3917 <= _3516;
        127:
            _3917 <= _3519;
        128:
            _3917 <= _3522;
        129:
            _3917 <= _3525;
        130:
            _3917 <= _3528;
        131:
            _3917 <= _3531;
        132:
            _3917 <= _3534;
        133:
            _3917 <= _3537;
        134:
            _3917 <= _3540;
        135:
            _3917 <= _3543;
        136:
            _3917 <= _3546;
        137:
            _3917 <= _3549;
        138:
            _3917 <= _3552;
        139:
            _3917 <= _3555;
        140:
            _3917 <= _3558;
        141:
            _3917 <= _3561;
        142:
            _3917 <= _3564;
        143:
            _3917 <= _3567;
        144:
            _3917 <= _3570;
        145:
            _3917 <= _3573;
        146:
            _3917 <= _3576;
        147:
            _3917 <= _3579;
        148:
            _3917 <= _3582;
        149:
            _3917 <= _3585;
        150:
            _3917 <= _3588;
        151:
            _3917 <= _3591;
        152:
            _3917 <= _3594;
        153:
            _3917 <= _3597;
        154:
            _3917 <= _3600;
        155:
            _3917 <= _3603;
        156:
            _3917 <= _3606;
        157:
            _3917 <= _3609;
        158:
            _3917 <= _3612;
        159:
            _3917 <= _3615;
        160:
            _3917 <= _3618;
        161:
            _3917 <= _3621;
        162:
            _3917 <= _3624;
        163:
            _3917 <= _3627;
        164:
            _3917 <= _3630;
        165:
            _3917 <= _3633;
        166:
            _3917 <= _3636;
        167:
            _3917 <= _3639;
        168:
            _3917 <= _3642;
        169:
            _3917 <= _3645;
        170:
            _3917 <= _3648;
        171:
            _3917 <= _3651;
        172:
            _3917 <= _3654;
        173:
            _3917 <= _3657;
        174:
            _3917 <= _3660;
        175:
            _3917 <= _3663;
        176:
            _3917 <= _3666;
        177:
            _3917 <= _3669;
        178:
            _3917 <= _3672;
        179:
            _3917 <= _3675;
        180:
            _3917 <= _3678;
        181:
            _3917 <= _3681;
        182:
            _3917 <= _3684;
        183:
            _3917 <= _3687;
        184:
            _3917 <= _3690;
        185:
            _3917 <= _3693;
        186:
            _3917 <= _3696;
        187:
            _3917 <= _3699;
        188:
            _3917 <= _3702;
        189:
            _3917 <= _3705;
        190:
            _3917 <= _3708;
        191:
            _3917 <= _3711;
        192:
            _3917 <= _3714;
        193:
            _3917 <= _3717;
        194:
            _3917 <= _3720;
        195:
            _3917 <= _3723;
        196:
            _3917 <= _3726;
        197:
            _3917 <= _3729;
        198:
            _3917 <= _3732;
        199:
            _3917 <= _3735;
        200:
            _3917 <= _3738;
        201:
            _3917 <= _3741;
        202:
            _3917 <= _3744;
        203:
            _3917 <= _3747;
        204:
            _3917 <= _3750;
        205:
            _3917 <= _3753;
        206:
            _3917 <= _3756;
        207:
            _3917 <= _3759;
        208:
            _3917 <= _3762;
        209:
            _3917 <= _3765;
        210:
            _3917 <= _3768;
        211:
            _3917 <= _3771;
        212:
            _3917 <= _3774;
        213:
            _3917 <= _3777;
        214:
            _3917 <= _3780;
        215:
            _3917 <= _3783;
        216:
            _3917 <= _3786;
        217:
            _3917 <= _3789;
        218:
            _3917 <= _3792;
        219:
            _3917 <= _3795;
        220:
            _3917 <= _3798;
        221:
            _3917 <= _3801;
        222:
            _3917 <= _3804;
        223:
            _3917 <= _3807;
        224:
            _3917 <= _3810;
        225:
            _3917 <= _3813;
        226:
            _3917 <= _3816;
        227:
            _3917 <= _3819;
        228:
            _3917 <= _3822;
        229:
            _3917 <= _3825;
        230:
            _3917 <= _3828;
        231:
            _3917 <= _3831;
        232:
            _3917 <= _3834;
        233:
            _3917 <= _3837;
        234:
            _3917 <= _3840;
        235:
            _3917 <= _3843;
        236:
            _3917 <= _3846;
        237:
            _3917 <= _3849;
        238:
            _3917 <= _3852;
        239:
            _3917 <= _3855;
        240:
            _3917 <= _3858;
        241:
            _3917 <= _3861;
        242:
            _3917 <= _3864;
        243:
            _3917 <= _3867;
        244:
            _3917 <= _3870;
        245:
            _3917 <= _3873;
        246:
            _3917 <= _3876;
        247:
            _3917 <= _3879;
        248:
            _3917 <= _3882;
        249:
            _3917 <= _3885;
        250:
            _3917 <= _3888;
        251:
            _3917 <= _3891;
        252:
            _3917 <= _3894;
        253:
            _3917 <= _3897;
        254:
            _3917 <= _3900;
        default:
            _3917 <= _3903;
        endcase
    end
    always @* begin
        case (_3917)
        0:
            _3918 <= _3138;
        1:
            _3918 <= _3141;
        2:
            _3918 <= _3144;
        3:
            _3918 <= _3147;
        4:
            _3918 <= _3150;
        5:
            _3918 <= _3153;
        6:
            _3918 <= _3156;
        7:
            _3918 <= _3159;
        8:
            _3918 <= _3162;
        9:
            _3918 <= _3165;
        10:
            _3918 <= _3168;
        11:
            _3918 <= _3171;
        12:
            _3918 <= _3174;
        13:
            _3918 <= _3177;
        14:
            _3918 <= _3180;
        15:
            _3918 <= _3183;
        16:
            _3918 <= _3186;
        17:
            _3918 <= _3189;
        18:
            _3918 <= _3192;
        19:
            _3918 <= _3195;
        20:
            _3918 <= _3198;
        21:
            _3918 <= _3201;
        22:
            _3918 <= _3204;
        23:
            _3918 <= _3207;
        24:
            _3918 <= _3210;
        25:
            _3918 <= _3213;
        26:
            _3918 <= _3216;
        27:
            _3918 <= _3219;
        28:
            _3918 <= _3222;
        29:
            _3918 <= _3225;
        30:
            _3918 <= _3228;
        31:
            _3918 <= _3231;
        32:
            _3918 <= _3234;
        33:
            _3918 <= _3237;
        34:
            _3918 <= _3240;
        35:
            _3918 <= _3243;
        36:
            _3918 <= _3246;
        37:
            _3918 <= _3249;
        38:
            _3918 <= _3252;
        39:
            _3918 <= _3255;
        40:
            _3918 <= _3258;
        41:
            _3918 <= _3261;
        42:
            _3918 <= _3264;
        43:
            _3918 <= _3267;
        44:
            _3918 <= _3270;
        45:
            _3918 <= _3273;
        46:
            _3918 <= _3276;
        47:
            _3918 <= _3279;
        48:
            _3918 <= _3282;
        49:
            _3918 <= _3285;
        50:
            _3918 <= _3288;
        51:
            _3918 <= _3291;
        52:
            _3918 <= _3294;
        53:
            _3918 <= _3297;
        54:
            _3918 <= _3300;
        55:
            _3918 <= _3303;
        56:
            _3918 <= _3306;
        57:
            _3918 <= _3309;
        58:
            _3918 <= _3312;
        59:
            _3918 <= _3315;
        60:
            _3918 <= _3318;
        61:
            _3918 <= _3321;
        62:
            _3918 <= _3324;
        63:
            _3918 <= _3327;
        64:
            _3918 <= _3330;
        65:
            _3918 <= _3333;
        66:
            _3918 <= _3336;
        67:
            _3918 <= _3339;
        68:
            _3918 <= _3342;
        69:
            _3918 <= _3345;
        70:
            _3918 <= _3348;
        71:
            _3918 <= _3351;
        72:
            _3918 <= _3354;
        73:
            _3918 <= _3357;
        74:
            _3918 <= _3360;
        75:
            _3918 <= _3363;
        76:
            _3918 <= _3366;
        77:
            _3918 <= _3369;
        78:
            _3918 <= _3372;
        79:
            _3918 <= _3375;
        80:
            _3918 <= _3378;
        81:
            _3918 <= _3381;
        82:
            _3918 <= _3384;
        83:
            _3918 <= _3387;
        84:
            _3918 <= _3390;
        85:
            _3918 <= _3393;
        86:
            _3918 <= _3396;
        87:
            _3918 <= _3399;
        88:
            _3918 <= _3402;
        89:
            _3918 <= _3405;
        90:
            _3918 <= _3408;
        91:
            _3918 <= _3411;
        92:
            _3918 <= _3414;
        93:
            _3918 <= _3417;
        94:
            _3918 <= _3420;
        95:
            _3918 <= _3423;
        96:
            _3918 <= _3426;
        97:
            _3918 <= _3429;
        98:
            _3918 <= _3432;
        99:
            _3918 <= _3435;
        100:
            _3918 <= _3438;
        101:
            _3918 <= _3441;
        102:
            _3918 <= _3444;
        103:
            _3918 <= _3447;
        104:
            _3918 <= _3450;
        105:
            _3918 <= _3453;
        106:
            _3918 <= _3456;
        107:
            _3918 <= _3459;
        108:
            _3918 <= _3462;
        109:
            _3918 <= _3465;
        110:
            _3918 <= _3468;
        111:
            _3918 <= _3471;
        112:
            _3918 <= _3474;
        113:
            _3918 <= _3477;
        114:
            _3918 <= _3480;
        115:
            _3918 <= _3483;
        116:
            _3918 <= _3486;
        117:
            _3918 <= _3489;
        118:
            _3918 <= _3492;
        119:
            _3918 <= _3495;
        120:
            _3918 <= _3498;
        121:
            _3918 <= _3501;
        122:
            _3918 <= _3504;
        123:
            _3918 <= _3507;
        124:
            _3918 <= _3510;
        125:
            _3918 <= _3513;
        126:
            _3918 <= _3516;
        127:
            _3918 <= _3519;
        128:
            _3918 <= _3522;
        129:
            _3918 <= _3525;
        130:
            _3918 <= _3528;
        131:
            _3918 <= _3531;
        132:
            _3918 <= _3534;
        133:
            _3918 <= _3537;
        134:
            _3918 <= _3540;
        135:
            _3918 <= _3543;
        136:
            _3918 <= _3546;
        137:
            _3918 <= _3549;
        138:
            _3918 <= _3552;
        139:
            _3918 <= _3555;
        140:
            _3918 <= _3558;
        141:
            _3918 <= _3561;
        142:
            _3918 <= _3564;
        143:
            _3918 <= _3567;
        144:
            _3918 <= _3570;
        145:
            _3918 <= _3573;
        146:
            _3918 <= _3576;
        147:
            _3918 <= _3579;
        148:
            _3918 <= _3582;
        149:
            _3918 <= _3585;
        150:
            _3918 <= _3588;
        151:
            _3918 <= _3591;
        152:
            _3918 <= _3594;
        153:
            _3918 <= _3597;
        154:
            _3918 <= _3600;
        155:
            _3918 <= _3603;
        156:
            _3918 <= _3606;
        157:
            _3918 <= _3609;
        158:
            _3918 <= _3612;
        159:
            _3918 <= _3615;
        160:
            _3918 <= _3618;
        161:
            _3918 <= _3621;
        162:
            _3918 <= _3624;
        163:
            _3918 <= _3627;
        164:
            _3918 <= _3630;
        165:
            _3918 <= _3633;
        166:
            _3918 <= _3636;
        167:
            _3918 <= _3639;
        168:
            _3918 <= _3642;
        169:
            _3918 <= _3645;
        170:
            _3918 <= _3648;
        171:
            _3918 <= _3651;
        172:
            _3918 <= _3654;
        173:
            _3918 <= _3657;
        174:
            _3918 <= _3660;
        175:
            _3918 <= _3663;
        176:
            _3918 <= _3666;
        177:
            _3918 <= _3669;
        178:
            _3918 <= _3672;
        179:
            _3918 <= _3675;
        180:
            _3918 <= _3678;
        181:
            _3918 <= _3681;
        182:
            _3918 <= _3684;
        183:
            _3918 <= _3687;
        184:
            _3918 <= _3690;
        185:
            _3918 <= _3693;
        186:
            _3918 <= _3696;
        187:
            _3918 <= _3699;
        188:
            _3918 <= _3702;
        189:
            _3918 <= _3705;
        190:
            _3918 <= _3708;
        191:
            _3918 <= _3711;
        192:
            _3918 <= _3714;
        193:
            _3918 <= _3717;
        194:
            _3918 <= _3720;
        195:
            _3918 <= _3723;
        196:
            _3918 <= _3726;
        197:
            _3918 <= _3729;
        198:
            _3918 <= _3732;
        199:
            _3918 <= _3735;
        200:
            _3918 <= _3738;
        201:
            _3918 <= _3741;
        202:
            _3918 <= _3744;
        203:
            _3918 <= _3747;
        204:
            _3918 <= _3750;
        205:
            _3918 <= _3753;
        206:
            _3918 <= _3756;
        207:
            _3918 <= _3759;
        208:
            _3918 <= _3762;
        209:
            _3918 <= _3765;
        210:
            _3918 <= _3768;
        211:
            _3918 <= _3771;
        212:
            _3918 <= _3774;
        213:
            _3918 <= _3777;
        214:
            _3918 <= _3780;
        215:
            _3918 <= _3783;
        216:
            _3918 <= _3786;
        217:
            _3918 <= _3789;
        218:
            _3918 <= _3792;
        219:
            _3918 <= _3795;
        220:
            _3918 <= _3798;
        221:
            _3918 <= _3801;
        222:
            _3918 <= _3804;
        223:
            _3918 <= _3807;
        224:
            _3918 <= _3810;
        225:
            _3918 <= _3813;
        226:
            _3918 <= _3816;
        227:
            _3918 <= _3819;
        228:
            _3918 <= _3822;
        229:
            _3918 <= _3825;
        230:
            _3918 <= _3828;
        231:
            _3918 <= _3831;
        232:
            _3918 <= _3834;
        233:
            _3918 <= _3837;
        234:
            _3918 <= _3840;
        235:
            _3918 <= _3843;
        236:
            _3918 <= _3846;
        237:
            _3918 <= _3849;
        238:
            _3918 <= _3852;
        239:
            _3918 <= _3855;
        240:
            _3918 <= _3858;
        241:
            _3918 <= _3861;
        242:
            _3918 <= _3864;
        243:
            _3918 <= _3867;
        244:
            _3918 <= _3870;
        245:
            _3918 <= _3873;
        246:
            _3918 <= _3876;
        247:
            _3918 <= _3879;
        248:
            _3918 <= _3882;
        249:
            _3918 <= _3885;
        250:
            _3918 <= _3888;
        251:
            _3918 <= _3891;
        252:
            _3918 <= _3894;
        253:
            _3918 <= _3897;
        254:
            _3918 <= _3900;
        default:
            _3918 <= _3903;
        endcase
    end
    always @* begin
        case (_3918)
        0:
            _3919 <= _3138;
        1:
            _3919 <= _3141;
        2:
            _3919 <= _3144;
        3:
            _3919 <= _3147;
        4:
            _3919 <= _3150;
        5:
            _3919 <= _3153;
        6:
            _3919 <= _3156;
        7:
            _3919 <= _3159;
        8:
            _3919 <= _3162;
        9:
            _3919 <= _3165;
        10:
            _3919 <= _3168;
        11:
            _3919 <= _3171;
        12:
            _3919 <= _3174;
        13:
            _3919 <= _3177;
        14:
            _3919 <= _3180;
        15:
            _3919 <= _3183;
        16:
            _3919 <= _3186;
        17:
            _3919 <= _3189;
        18:
            _3919 <= _3192;
        19:
            _3919 <= _3195;
        20:
            _3919 <= _3198;
        21:
            _3919 <= _3201;
        22:
            _3919 <= _3204;
        23:
            _3919 <= _3207;
        24:
            _3919 <= _3210;
        25:
            _3919 <= _3213;
        26:
            _3919 <= _3216;
        27:
            _3919 <= _3219;
        28:
            _3919 <= _3222;
        29:
            _3919 <= _3225;
        30:
            _3919 <= _3228;
        31:
            _3919 <= _3231;
        32:
            _3919 <= _3234;
        33:
            _3919 <= _3237;
        34:
            _3919 <= _3240;
        35:
            _3919 <= _3243;
        36:
            _3919 <= _3246;
        37:
            _3919 <= _3249;
        38:
            _3919 <= _3252;
        39:
            _3919 <= _3255;
        40:
            _3919 <= _3258;
        41:
            _3919 <= _3261;
        42:
            _3919 <= _3264;
        43:
            _3919 <= _3267;
        44:
            _3919 <= _3270;
        45:
            _3919 <= _3273;
        46:
            _3919 <= _3276;
        47:
            _3919 <= _3279;
        48:
            _3919 <= _3282;
        49:
            _3919 <= _3285;
        50:
            _3919 <= _3288;
        51:
            _3919 <= _3291;
        52:
            _3919 <= _3294;
        53:
            _3919 <= _3297;
        54:
            _3919 <= _3300;
        55:
            _3919 <= _3303;
        56:
            _3919 <= _3306;
        57:
            _3919 <= _3309;
        58:
            _3919 <= _3312;
        59:
            _3919 <= _3315;
        60:
            _3919 <= _3318;
        61:
            _3919 <= _3321;
        62:
            _3919 <= _3324;
        63:
            _3919 <= _3327;
        64:
            _3919 <= _3330;
        65:
            _3919 <= _3333;
        66:
            _3919 <= _3336;
        67:
            _3919 <= _3339;
        68:
            _3919 <= _3342;
        69:
            _3919 <= _3345;
        70:
            _3919 <= _3348;
        71:
            _3919 <= _3351;
        72:
            _3919 <= _3354;
        73:
            _3919 <= _3357;
        74:
            _3919 <= _3360;
        75:
            _3919 <= _3363;
        76:
            _3919 <= _3366;
        77:
            _3919 <= _3369;
        78:
            _3919 <= _3372;
        79:
            _3919 <= _3375;
        80:
            _3919 <= _3378;
        81:
            _3919 <= _3381;
        82:
            _3919 <= _3384;
        83:
            _3919 <= _3387;
        84:
            _3919 <= _3390;
        85:
            _3919 <= _3393;
        86:
            _3919 <= _3396;
        87:
            _3919 <= _3399;
        88:
            _3919 <= _3402;
        89:
            _3919 <= _3405;
        90:
            _3919 <= _3408;
        91:
            _3919 <= _3411;
        92:
            _3919 <= _3414;
        93:
            _3919 <= _3417;
        94:
            _3919 <= _3420;
        95:
            _3919 <= _3423;
        96:
            _3919 <= _3426;
        97:
            _3919 <= _3429;
        98:
            _3919 <= _3432;
        99:
            _3919 <= _3435;
        100:
            _3919 <= _3438;
        101:
            _3919 <= _3441;
        102:
            _3919 <= _3444;
        103:
            _3919 <= _3447;
        104:
            _3919 <= _3450;
        105:
            _3919 <= _3453;
        106:
            _3919 <= _3456;
        107:
            _3919 <= _3459;
        108:
            _3919 <= _3462;
        109:
            _3919 <= _3465;
        110:
            _3919 <= _3468;
        111:
            _3919 <= _3471;
        112:
            _3919 <= _3474;
        113:
            _3919 <= _3477;
        114:
            _3919 <= _3480;
        115:
            _3919 <= _3483;
        116:
            _3919 <= _3486;
        117:
            _3919 <= _3489;
        118:
            _3919 <= _3492;
        119:
            _3919 <= _3495;
        120:
            _3919 <= _3498;
        121:
            _3919 <= _3501;
        122:
            _3919 <= _3504;
        123:
            _3919 <= _3507;
        124:
            _3919 <= _3510;
        125:
            _3919 <= _3513;
        126:
            _3919 <= _3516;
        127:
            _3919 <= _3519;
        128:
            _3919 <= _3522;
        129:
            _3919 <= _3525;
        130:
            _3919 <= _3528;
        131:
            _3919 <= _3531;
        132:
            _3919 <= _3534;
        133:
            _3919 <= _3537;
        134:
            _3919 <= _3540;
        135:
            _3919 <= _3543;
        136:
            _3919 <= _3546;
        137:
            _3919 <= _3549;
        138:
            _3919 <= _3552;
        139:
            _3919 <= _3555;
        140:
            _3919 <= _3558;
        141:
            _3919 <= _3561;
        142:
            _3919 <= _3564;
        143:
            _3919 <= _3567;
        144:
            _3919 <= _3570;
        145:
            _3919 <= _3573;
        146:
            _3919 <= _3576;
        147:
            _3919 <= _3579;
        148:
            _3919 <= _3582;
        149:
            _3919 <= _3585;
        150:
            _3919 <= _3588;
        151:
            _3919 <= _3591;
        152:
            _3919 <= _3594;
        153:
            _3919 <= _3597;
        154:
            _3919 <= _3600;
        155:
            _3919 <= _3603;
        156:
            _3919 <= _3606;
        157:
            _3919 <= _3609;
        158:
            _3919 <= _3612;
        159:
            _3919 <= _3615;
        160:
            _3919 <= _3618;
        161:
            _3919 <= _3621;
        162:
            _3919 <= _3624;
        163:
            _3919 <= _3627;
        164:
            _3919 <= _3630;
        165:
            _3919 <= _3633;
        166:
            _3919 <= _3636;
        167:
            _3919 <= _3639;
        168:
            _3919 <= _3642;
        169:
            _3919 <= _3645;
        170:
            _3919 <= _3648;
        171:
            _3919 <= _3651;
        172:
            _3919 <= _3654;
        173:
            _3919 <= _3657;
        174:
            _3919 <= _3660;
        175:
            _3919 <= _3663;
        176:
            _3919 <= _3666;
        177:
            _3919 <= _3669;
        178:
            _3919 <= _3672;
        179:
            _3919 <= _3675;
        180:
            _3919 <= _3678;
        181:
            _3919 <= _3681;
        182:
            _3919 <= _3684;
        183:
            _3919 <= _3687;
        184:
            _3919 <= _3690;
        185:
            _3919 <= _3693;
        186:
            _3919 <= _3696;
        187:
            _3919 <= _3699;
        188:
            _3919 <= _3702;
        189:
            _3919 <= _3705;
        190:
            _3919 <= _3708;
        191:
            _3919 <= _3711;
        192:
            _3919 <= _3714;
        193:
            _3919 <= _3717;
        194:
            _3919 <= _3720;
        195:
            _3919 <= _3723;
        196:
            _3919 <= _3726;
        197:
            _3919 <= _3729;
        198:
            _3919 <= _3732;
        199:
            _3919 <= _3735;
        200:
            _3919 <= _3738;
        201:
            _3919 <= _3741;
        202:
            _3919 <= _3744;
        203:
            _3919 <= _3747;
        204:
            _3919 <= _3750;
        205:
            _3919 <= _3753;
        206:
            _3919 <= _3756;
        207:
            _3919 <= _3759;
        208:
            _3919 <= _3762;
        209:
            _3919 <= _3765;
        210:
            _3919 <= _3768;
        211:
            _3919 <= _3771;
        212:
            _3919 <= _3774;
        213:
            _3919 <= _3777;
        214:
            _3919 <= _3780;
        215:
            _3919 <= _3783;
        216:
            _3919 <= _3786;
        217:
            _3919 <= _3789;
        218:
            _3919 <= _3792;
        219:
            _3919 <= _3795;
        220:
            _3919 <= _3798;
        221:
            _3919 <= _3801;
        222:
            _3919 <= _3804;
        223:
            _3919 <= _3807;
        224:
            _3919 <= _3810;
        225:
            _3919 <= _3813;
        226:
            _3919 <= _3816;
        227:
            _3919 <= _3819;
        228:
            _3919 <= _3822;
        229:
            _3919 <= _3825;
        230:
            _3919 <= _3828;
        231:
            _3919 <= _3831;
        232:
            _3919 <= _3834;
        233:
            _3919 <= _3837;
        234:
            _3919 <= _3840;
        235:
            _3919 <= _3843;
        236:
            _3919 <= _3846;
        237:
            _3919 <= _3849;
        238:
            _3919 <= _3852;
        239:
            _3919 <= _3855;
        240:
            _3919 <= _3858;
        241:
            _3919 <= _3861;
        242:
            _3919 <= _3864;
        243:
            _3919 <= _3867;
        244:
            _3919 <= _3870;
        245:
            _3919 <= _3873;
        246:
            _3919 <= _3876;
        247:
            _3919 <= _3879;
        248:
            _3919 <= _3882;
        249:
            _3919 <= _3885;
        250:
            _3919 <= _3888;
        251:
            _3919 <= _3891;
        252:
            _3919 <= _3894;
        253:
            _3919 <= _3897;
        254:
            _3919 <= _3900;
        default:
            _3919 <= _3903;
        endcase
    end
    assign _5304 = _5303 ? _3911 : _3919;
    assign _11937 = _5304 == _3118;
    assign _11934 = ~ _3920;
    assign _11935 = _3135 & _11934;
    assign _11938 = _11935 & _11937;
    assign _11939 = _11938 ? _4693 : _3925;
    assign _11932 = _5296 == _3118;
    assign _11933 = _5293 & _11932;
    assign _11941 = _11933 ? _11940 : _11939;
    assign _11943 = _805 ? _4718 : _11941;
    assign _782 = _11943;
    always @(posedge _791) begin
        if (_789)
            _3925 <= _4718;
        else
            _3925 <= _782;
    end
    always @* begin
        case (_3911)
        0:
            _4691 <= _3925;
        1:
            _4691 <= _3928;
        2:
            _4691 <= _3931;
        3:
            _4691 <= _3934;
        4:
            _4691 <= _3937;
        5:
            _4691 <= _3940;
        6:
            _4691 <= _3943;
        7:
            _4691 <= _3946;
        8:
            _4691 <= _3949;
        9:
            _4691 <= _3952;
        10:
            _4691 <= _3955;
        11:
            _4691 <= _3958;
        12:
            _4691 <= _3961;
        13:
            _4691 <= _3964;
        14:
            _4691 <= _3967;
        15:
            _4691 <= _3970;
        16:
            _4691 <= _3973;
        17:
            _4691 <= _3976;
        18:
            _4691 <= _3979;
        19:
            _4691 <= _3982;
        20:
            _4691 <= _3985;
        21:
            _4691 <= _3988;
        22:
            _4691 <= _3991;
        23:
            _4691 <= _3994;
        24:
            _4691 <= _3997;
        25:
            _4691 <= _4000;
        26:
            _4691 <= _4003;
        27:
            _4691 <= _4006;
        28:
            _4691 <= _4009;
        29:
            _4691 <= _4012;
        30:
            _4691 <= _4015;
        31:
            _4691 <= _4018;
        32:
            _4691 <= _4021;
        33:
            _4691 <= _4024;
        34:
            _4691 <= _4027;
        35:
            _4691 <= _4030;
        36:
            _4691 <= _4033;
        37:
            _4691 <= _4036;
        38:
            _4691 <= _4039;
        39:
            _4691 <= _4042;
        40:
            _4691 <= _4045;
        41:
            _4691 <= _4048;
        42:
            _4691 <= _4051;
        43:
            _4691 <= _4054;
        44:
            _4691 <= _4057;
        45:
            _4691 <= _4060;
        46:
            _4691 <= _4063;
        47:
            _4691 <= _4066;
        48:
            _4691 <= _4069;
        49:
            _4691 <= _4072;
        50:
            _4691 <= _4075;
        51:
            _4691 <= _4078;
        52:
            _4691 <= _4081;
        53:
            _4691 <= _4084;
        54:
            _4691 <= _4087;
        55:
            _4691 <= _4090;
        56:
            _4691 <= _4093;
        57:
            _4691 <= _4096;
        58:
            _4691 <= _4099;
        59:
            _4691 <= _4102;
        60:
            _4691 <= _4105;
        61:
            _4691 <= _4108;
        62:
            _4691 <= _4111;
        63:
            _4691 <= _4114;
        64:
            _4691 <= _4117;
        65:
            _4691 <= _4120;
        66:
            _4691 <= _4123;
        67:
            _4691 <= _4126;
        68:
            _4691 <= _4129;
        69:
            _4691 <= _4132;
        70:
            _4691 <= _4135;
        71:
            _4691 <= _4138;
        72:
            _4691 <= _4141;
        73:
            _4691 <= _4144;
        74:
            _4691 <= _4147;
        75:
            _4691 <= _4150;
        76:
            _4691 <= _4153;
        77:
            _4691 <= _4156;
        78:
            _4691 <= _4159;
        79:
            _4691 <= _4162;
        80:
            _4691 <= _4165;
        81:
            _4691 <= _4168;
        82:
            _4691 <= _4171;
        83:
            _4691 <= _4174;
        84:
            _4691 <= _4177;
        85:
            _4691 <= _4180;
        86:
            _4691 <= _4183;
        87:
            _4691 <= _4186;
        88:
            _4691 <= _4189;
        89:
            _4691 <= _4192;
        90:
            _4691 <= _4195;
        91:
            _4691 <= _4198;
        92:
            _4691 <= _4201;
        93:
            _4691 <= _4204;
        94:
            _4691 <= _4207;
        95:
            _4691 <= _4210;
        96:
            _4691 <= _4213;
        97:
            _4691 <= _4216;
        98:
            _4691 <= _4219;
        99:
            _4691 <= _4222;
        100:
            _4691 <= _4225;
        101:
            _4691 <= _4228;
        102:
            _4691 <= _4231;
        103:
            _4691 <= _4234;
        104:
            _4691 <= _4237;
        105:
            _4691 <= _4240;
        106:
            _4691 <= _4243;
        107:
            _4691 <= _4246;
        108:
            _4691 <= _4249;
        109:
            _4691 <= _4252;
        110:
            _4691 <= _4255;
        111:
            _4691 <= _4258;
        112:
            _4691 <= _4261;
        113:
            _4691 <= _4264;
        114:
            _4691 <= _4267;
        115:
            _4691 <= _4270;
        116:
            _4691 <= _4273;
        117:
            _4691 <= _4276;
        118:
            _4691 <= _4279;
        119:
            _4691 <= _4282;
        120:
            _4691 <= _4285;
        121:
            _4691 <= _4288;
        122:
            _4691 <= _4291;
        123:
            _4691 <= _4294;
        124:
            _4691 <= _4297;
        125:
            _4691 <= _4300;
        126:
            _4691 <= _4303;
        127:
            _4691 <= _4306;
        128:
            _4691 <= _4309;
        129:
            _4691 <= _4312;
        130:
            _4691 <= _4315;
        131:
            _4691 <= _4318;
        132:
            _4691 <= _4321;
        133:
            _4691 <= _4324;
        134:
            _4691 <= _4327;
        135:
            _4691 <= _4330;
        136:
            _4691 <= _4333;
        137:
            _4691 <= _4336;
        138:
            _4691 <= _4339;
        139:
            _4691 <= _4342;
        140:
            _4691 <= _4345;
        141:
            _4691 <= _4348;
        142:
            _4691 <= _4351;
        143:
            _4691 <= _4354;
        144:
            _4691 <= _4357;
        145:
            _4691 <= _4360;
        146:
            _4691 <= _4363;
        147:
            _4691 <= _4366;
        148:
            _4691 <= _4369;
        149:
            _4691 <= _4372;
        150:
            _4691 <= _4375;
        151:
            _4691 <= _4378;
        152:
            _4691 <= _4381;
        153:
            _4691 <= _4384;
        154:
            _4691 <= _4387;
        155:
            _4691 <= _4390;
        156:
            _4691 <= _4393;
        157:
            _4691 <= _4396;
        158:
            _4691 <= _4399;
        159:
            _4691 <= _4402;
        160:
            _4691 <= _4405;
        161:
            _4691 <= _4408;
        162:
            _4691 <= _4411;
        163:
            _4691 <= _4414;
        164:
            _4691 <= _4417;
        165:
            _4691 <= _4420;
        166:
            _4691 <= _4423;
        167:
            _4691 <= _4426;
        168:
            _4691 <= _4429;
        169:
            _4691 <= _4432;
        170:
            _4691 <= _4435;
        171:
            _4691 <= _4438;
        172:
            _4691 <= _4441;
        173:
            _4691 <= _4444;
        174:
            _4691 <= _4447;
        175:
            _4691 <= _4450;
        176:
            _4691 <= _4453;
        177:
            _4691 <= _4456;
        178:
            _4691 <= _4459;
        179:
            _4691 <= _4462;
        180:
            _4691 <= _4465;
        181:
            _4691 <= _4468;
        182:
            _4691 <= _4471;
        183:
            _4691 <= _4474;
        184:
            _4691 <= _4477;
        185:
            _4691 <= _4480;
        186:
            _4691 <= _4483;
        187:
            _4691 <= _4486;
        188:
            _4691 <= _4489;
        189:
            _4691 <= _4492;
        190:
            _4691 <= _4495;
        191:
            _4691 <= _4498;
        192:
            _4691 <= _4501;
        193:
            _4691 <= _4504;
        194:
            _4691 <= _4507;
        195:
            _4691 <= _4510;
        196:
            _4691 <= _4513;
        197:
            _4691 <= _4516;
        198:
            _4691 <= _4519;
        199:
            _4691 <= _4522;
        200:
            _4691 <= _4525;
        201:
            _4691 <= _4528;
        202:
            _4691 <= _4531;
        203:
            _4691 <= _4534;
        204:
            _4691 <= _4537;
        205:
            _4691 <= _4540;
        206:
            _4691 <= _4543;
        207:
            _4691 <= _4546;
        208:
            _4691 <= _4549;
        209:
            _4691 <= _4552;
        210:
            _4691 <= _4555;
        211:
            _4691 <= _4558;
        212:
            _4691 <= _4561;
        213:
            _4691 <= _4564;
        214:
            _4691 <= _4567;
        215:
            _4691 <= _4570;
        216:
            _4691 <= _4573;
        217:
            _4691 <= _4576;
        218:
            _4691 <= _4579;
        219:
            _4691 <= _4582;
        220:
            _4691 <= _4585;
        221:
            _4691 <= _4588;
        222:
            _4691 <= _4591;
        223:
            _4691 <= _4594;
        224:
            _4691 <= _4597;
        225:
            _4691 <= _4600;
        226:
            _4691 <= _4603;
        227:
            _4691 <= _4606;
        228:
            _4691 <= _4609;
        229:
            _4691 <= _4612;
        230:
            _4691 <= _4615;
        231:
            _4691 <= _4618;
        232:
            _4691 <= _4621;
        233:
            _4691 <= _4624;
        234:
            _4691 <= _4627;
        235:
            _4691 <= _4630;
        236:
            _4691 <= _4633;
        237:
            _4691 <= _4636;
        238:
            _4691 <= _4639;
        239:
            _4691 <= _4642;
        240:
            _4691 <= _4645;
        241:
            _4691 <= _4648;
        242:
            _4691 <= _4651;
        243:
            _4691 <= _4654;
        244:
            _4691 <= _4657;
        245:
            _4691 <= _4660;
        246:
            _4691 <= _4663;
        247:
            _4691 <= _4666;
        248:
            _4691 <= _4669;
        249:
            _4691 <= _4672;
        250:
            _4691 <= _4675;
        251:
            _4691 <= _4678;
        252:
            _4691 <= _4681;
        253:
            _4691 <= _4684;
        254:
            _4691 <= _4687;
        default:
            _4691 <= _4690;
        endcase
    end
    assign _5302 = _4691 < _4692;
    assign _5303 = ~ _5302;
    assign _8620 = _5303 ? _3919 : _3911;
    assign _11950 = _8620 == _3118;
    assign _11947 = ~ _3920;
    assign _11948 = _3135 & _11947;
    assign _11951 = _11948 & _11950;
    assign _11952 = _11951 ? _5304 : _3138;
    assign _11945 = _5296 == _3118;
    assign _11946 = _5293 & _11945;
    assign _11954 = _11946 ? _3118 : _11952;
    assign _11956 = _805 ? _3118 : _11954;
    assign _783 = _11956;
    always @(posedge _791) begin
        if (_789)
            _3138 <= _3118;
        else
            _3138 <= _783;
    end
    assign _785 = edge_i;
    always @* begin
        case (_785)
        0:
            _3904 <= _3138;
        1:
            _3904 <= _3141;
        2:
            _3904 <= _3144;
        3:
            _3904 <= _3147;
        4:
            _3904 <= _3150;
        5:
            _3904 <= _3153;
        6:
            _3904 <= _3156;
        7:
            _3904 <= _3159;
        8:
            _3904 <= _3162;
        9:
            _3904 <= _3165;
        10:
            _3904 <= _3168;
        11:
            _3904 <= _3171;
        12:
            _3904 <= _3174;
        13:
            _3904 <= _3177;
        14:
            _3904 <= _3180;
        15:
            _3904 <= _3183;
        16:
            _3904 <= _3186;
        17:
            _3904 <= _3189;
        18:
            _3904 <= _3192;
        19:
            _3904 <= _3195;
        20:
            _3904 <= _3198;
        21:
            _3904 <= _3201;
        22:
            _3904 <= _3204;
        23:
            _3904 <= _3207;
        24:
            _3904 <= _3210;
        25:
            _3904 <= _3213;
        26:
            _3904 <= _3216;
        27:
            _3904 <= _3219;
        28:
            _3904 <= _3222;
        29:
            _3904 <= _3225;
        30:
            _3904 <= _3228;
        31:
            _3904 <= _3231;
        32:
            _3904 <= _3234;
        33:
            _3904 <= _3237;
        34:
            _3904 <= _3240;
        35:
            _3904 <= _3243;
        36:
            _3904 <= _3246;
        37:
            _3904 <= _3249;
        38:
            _3904 <= _3252;
        39:
            _3904 <= _3255;
        40:
            _3904 <= _3258;
        41:
            _3904 <= _3261;
        42:
            _3904 <= _3264;
        43:
            _3904 <= _3267;
        44:
            _3904 <= _3270;
        45:
            _3904 <= _3273;
        46:
            _3904 <= _3276;
        47:
            _3904 <= _3279;
        48:
            _3904 <= _3282;
        49:
            _3904 <= _3285;
        50:
            _3904 <= _3288;
        51:
            _3904 <= _3291;
        52:
            _3904 <= _3294;
        53:
            _3904 <= _3297;
        54:
            _3904 <= _3300;
        55:
            _3904 <= _3303;
        56:
            _3904 <= _3306;
        57:
            _3904 <= _3309;
        58:
            _3904 <= _3312;
        59:
            _3904 <= _3315;
        60:
            _3904 <= _3318;
        61:
            _3904 <= _3321;
        62:
            _3904 <= _3324;
        63:
            _3904 <= _3327;
        64:
            _3904 <= _3330;
        65:
            _3904 <= _3333;
        66:
            _3904 <= _3336;
        67:
            _3904 <= _3339;
        68:
            _3904 <= _3342;
        69:
            _3904 <= _3345;
        70:
            _3904 <= _3348;
        71:
            _3904 <= _3351;
        72:
            _3904 <= _3354;
        73:
            _3904 <= _3357;
        74:
            _3904 <= _3360;
        75:
            _3904 <= _3363;
        76:
            _3904 <= _3366;
        77:
            _3904 <= _3369;
        78:
            _3904 <= _3372;
        79:
            _3904 <= _3375;
        80:
            _3904 <= _3378;
        81:
            _3904 <= _3381;
        82:
            _3904 <= _3384;
        83:
            _3904 <= _3387;
        84:
            _3904 <= _3390;
        85:
            _3904 <= _3393;
        86:
            _3904 <= _3396;
        87:
            _3904 <= _3399;
        88:
            _3904 <= _3402;
        89:
            _3904 <= _3405;
        90:
            _3904 <= _3408;
        91:
            _3904 <= _3411;
        92:
            _3904 <= _3414;
        93:
            _3904 <= _3417;
        94:
            _3904 <= _3420;
        95:
            _3904 <= _3423;
        96:
            _3904 <= _3426;
        97:
            _3904 <= _3429;
        98:
            _3904 <= _3432;
        99:
            _3904 <= _3435;
        100:
            _3904 <= _3438;
        101:
            _3904 <= _3441;
        102:
            _3904 <= _3444;
        103:
            _3904 <= _3447;
        104:
            _3904 <= _3450;
        105:
            _3904 <= _3453;
        106:
            _3904 <= _3456;
        107:
            _3904 <= _3459;
        108:
            _3904 <= _3462;
        109:
            _3904 <= _3465;
        110:
            _3904 <= _3468;
        111:
            _3904 <= _3471;
        112:
            _3904 <= _3474;
        113:
            _3904 <= _3477;
        114:
            _3904 <= _3480;
        115:
            _3904 <= _3483;
        116:
            _3904 <= _3486;
        117:
            _3904 <= _3489;
        118:
            _3904 <= _3492;
        119:
            _3904 <= _3495;
        120:
            _3904 <= _3498;
        121:
            _3904 <= _3501;
        122:
            _3904 <= _3504;
        123:
            _3904 <= _3507;
        124:
            _3904 <= _3510;
        125:
            _3904 <= _3513;
        126:
            _3904 <= _3516;
        127:
            _3904 <= _3519;
        128:
            _3904 <= _3522;
        129:
            _3904 <= _3525;
        130:
            _3904 <= _3528;
        131:
            _3904 <= _3531;
        132:
            _3904 <= _3534;
        133:
            _3904 <= _3537;
        134:
            _3904 <= _3540;
        135:
            _3904 <= _3543;
        136:
            _3904 <= _3546;
        137:
            _3904 <= _3549;
        138:
            _3904 <= _3552;
        139:
            _3904 <= _3555;
        140:
            _3904 <= _3558;
        141:
            _3904 <= _3561;
        142:
            _3904 <= _3564;
        143:
            _3904 <= _3567;
        144:
            _3904 <= _3570;
        145:
            _3904 <= _3573;
        146:
            _3904 <= _3576;
        147:
            _3904 <= _3579;
        148:
            _3904 <= _3582;
        149:
            _3904 <= _3585;
        150:
            _3904 <= _3588;
        151:
            _3904 <= _3591;
        152:
            _3904 <= _3594;
        153:
            _3904 <= _3597;
        154:
            _3904 <= _3600;
        155:
            _3904 <= _3603;
        156:
            _3904 <= _3606;
        157:
            _3904 <= _3609;
        158:
            _3904 <= _3612;
        159:
            _3904 <= _3615;
        160:
            _3904 <= _3618;
        161:
            _3904 <= _3621;
        162:
            _3904 <= _3624;
        163:
            _3904 <= _3627;
        164:
            _3904 <= _3630;
        165:
            _3904 <= _3633;
        166:
            _3904 <= _3636;
        167:
            _3904 <= _3639;
        168:
            _3904 <= _3642;
        169:
            _3904 <= _3645;
        170:
            _3904 <= _3648;
        171:
            _3904 <= _3651;
        172:
            _3904 <= _3654;
        173:
            _3904 <= _3657;
        174:
            _3904 <= _3660;
        175:
            _3904 <= _3663;
        176:
            _3904 <= _3666;
        177:
            _3904 <= _3669;
        178:
            _3904 <= _3672;
        179:
            _3904 <= _3675;
        180:
            _3904 <= _3678;
        181:
            _3904 <= _3681;
        182:
            _3904 <= _3684;
        183:
            _3904 <= _3687;
        184:
            _3904 <= _3690;
        185:
            _3904 <= _3693;
        186:
            _3904 <= _3696;
        187:
            _3904 <= _3699;
        188:
            _3904 <= _3702;
        189:
            _3904 <= _3705;
        190:
            _3904 <= _3708;
        191:
            _3904 <= _3711;
        192:
            _3904 <= _3714;
        193:
            _3904 <= _3717;
        194:
            _3904 <= _3720;
        195:
            _3904 <= _3723;
        196:
            _3904 <= _3726;
        197:
            _3904 <= _3729;
        198:
            _3904 <= _3732;
        199:
            _3904 <= _3735;
        200:
            _3904 <= _3738;
        201:
            _3904 <= _3741;
        202:
            _3904 <= _3744;
        203:
            _3904 <= _3747;
        204:
            _3904 <= _3750;
        205:
            _3904 <= _3753;
        206:
            _3904 <= _3756;
        207:
            _3904 <= _3759;
        208:
            _3904 <= _3762;
        209:
            _3904 <= _3765;
        210:
            _3904 <= _3768;
        211:
            _3904 <= _3771;
        212:
            _3904 <= _3774;
        213:
            _3904 <= _3777;
        214:
            _3904 <= _3780;
        215:
            _3904 <= _3783;
        216:
            _3904 <= _3786;
        217:
            _3904 <= _3789;
        218:
            _3904 <= _3792;
        219:
            _3904 <= _3795;
        220:
            _3904 <= _3798;
        221:
            _3904 <= _3801;
        222:
            _3904 <= _3804;
        223:
            _3904 <= _3807;
        224:
            _3904 <= _3810;
        225:
            _3904 <= _3813;
        226:
            _3904 <= _3816;
        227:
            _3904 <= _3819;
        228:
            _3904 <= _3822;
        229:
            _3904 <= _3825;
        230:
            _3904 <= _3828;
        231:
            _3904 <= _3831;
        232:
            _3904 <= _3834;
        233:
            _3904 <= _3837;
        234:
            _3904 <= _3840;
        235:
            _3904 <= _3843;
        236:
            _3904 <= _3846;
        237:
            _3904 <= _3849;
        238:
            _3904 <= _3852;
        239:
            _3904 <= _3855;
        240:
            _3904 <= _3858;
        241:
            _3904 <= _3861;
        242:
            _3904 <= _3864;
        243:
            _3904 <= _3867;
        244:
            _3904 <= _3870;
        245:
            _3904 <= _3873;
        246:
            _3904 <= _3876;
        247:
            _3904 <= _3879;
        248:
            _3904 <= _3882;
        249:
            _3904 <= _3885;
        250:
            _3904 <= _3888;
        251:
            _3904 <= _3891;
        252:
            _3904 <= _3894;
        253:
            _3904 <= _3897;
        254:
            _3904 <= _3900;
        default:
            _3904 <= _3903;
        endcase
    end
    always @* begin
        case (_3904)
        0:
            _3905 <= _3138;
        1:
            _3905 <= _3141;
        2:
            _3905 <= _3144;
        3:
            _3905 <= _3147;
        4:
            _3905 <= _3150;
        5:
            _3905 <= _3153;
        6:
            _3905 <= _3156;
        7:
            _3905 <= _3159;
        8:
            _3905 <= _3162;
        9:
            _3905 <= _3165;
        10:
            _3905 <= _3168;
        11:
            _3905 <= _3171;
        12:
            _3905 <= _3174;
        13:
            _3905 <= _3177;
        14:
            _3905 <= _3180;
        15:
            _3905 <= _3183;
        16:
            _3905 <= _3186;
        17:
            _3905 <= _3189;
        18:
            _3905 <= _3192;
        19:
            _3905 <= _3195;
        20:
            _3905 <= _3198;
        21:
            _3905 <= _3201;
        22:
            _3905 <= _3204;
        23:
            _3905 <= _3207;
        24:
            _3905 <= _3210;
        25:
            _3905 <= _3213;
        26:
            _3905 <= _3216;
        27:
            _3905 <= _3219;
        28:
            _3905 <= _3222;
        29:
            _3905 <= _3225;
        30:
            _3905 <= _3228;
        31:
            _3905 <= _3231;
        32:
            _3905 <= _3234;
        33:
            _3905 <= _3237;
        34:
            _3905 <= _3240;
        35:
            _3905 <= _3243;
        36:
            _3905 <= _3246;
        37:
            _3905 <= _3249;
        38:
            _3905 <= _3252;
        39:
            _3905 <= _3255;
        40:
            _3905 <= _3258;
        41:
            _3905 <= _3261;
        42:
            _3905 <= _3264;
        43:
            _3905 <= _3267;
        44:
            _3905 <= _3270;
        45:
            _3905 <= _3273;
        46:
            _3905 <= _3276;
        47:
            _3905 <= _3279;
        48:
            _3905 <= _3282;
        49:
            _3905 <= _3285;
        50:
            _3905 <= _3288;
        51:
            _3905 <= _3291;
        52:
            _3905 <= _3294;
        53:
            _3905 <= _3297;
        54:
            _3905 <= _3300;
        55:
            _3905 <= _3303;
        56:
            _3905 <= _3306;
        57:
            _3905 <= _3309;
        58:
            _3905 <= _3312;
        59:
            _3905 <= _3315;
        60:
            _3905 <= _3318;
        61:
            _3905 <= _3321;
        62:
            _3905 <= _3324;
        63:
            _3905 <= _3327;
        64:
            _3905 <= _3330;
        65:
            _3905 <= _3333;
        66:
            _3905 <= _3336;
        67:
            _3905 <= _3339;
        68:
            _3905 <= _3342;
        69:
            _3905 <= _3345;
        70:
            _3905 <= _3348;
        71:
            _3905 <= _3351;
        72:
            _3905 <= _3354;
        73:
            _3905 <= _3357;
        74:
            _3905 <= _3360;
        75:
            _3905 <= _3363;
        76:
            _3905 <= _3366;
        77:
            _3905 <= _3369;
        78:
            _3905 <= _3372;
        79:
            _3905 <= _3375;
        80:
            _3905 <= _3378;
        81:
            _3905 <= _3381;
        82:
            _3905 <= _3384;
        83:
            _3905 <= _3387;
        84:
            _3905 <= _3390;
        85:
            _3905 <= _3393;
        86:
            _3905 <= _3396;
        87:
            _3905 <= _3399;
        88:
            _3905 <= _3402;
        89:
            _3905 <= _3405;
        90:
            _3905 <= _3408;
        91:
            _3905 <= _3411;
        92:
            _3905 <= _3414;
        93:
            _3905 <= _3417;
        94:
            _3905 <= _3420;
        95:
            _3905 <= _3423;
        96:
            _3905 <= _3426;
        97:
            _3905 <= _3429;
        98:
            _3905 <= _3432;
        99:
            _3905 <= _3435;
        100:
            _3905 <= _3438;
        101:
            _3905 <= _3441;
        102:
            _3905 <= _3444;
        103:
            _3905 <= _3447;
        104:
            _3905 <= _3450;
        105:
            _3905 <= _3453;
        106:
            _3905 <= _3456;
        107:
            _3905 <= _3459;
        108:
            _3905 <= _3462;
        109:
            _3905 <= _3465;
        110:
            _3905 <= _3468;
        111:
            _3905 <= _3471;
        112:
            _3905 <= _3474;
        113:
            _3905 <= _3477;
        114:
            _3905 <= _3480;
        115:
            _3905 <= _3483;
        116:
            _3905 <= _3486;
        117:
            _3905 <= _3489;
        118:
            _3905 <= _3492;
        119:
            _3905 <= _3495;
        120:
            _3905 <= _3498;
        121:
            _3905 <= _3501;
        122:
            _3905 <= _3504;
        123:
            _3905 <= _3507;
        124:
            _3905 <= _3510;
        125:
            _3905 <= _3513;
        126:
            _3905 <= _3516;
        127:
            _3905 <= _3519;
        128:
            _3905 <= _3522;
        129:
            _3905 <= _3525;
        130:
            _3905 <= _3528;
        131:
            _3905 <= _3531;
        132:
            _3905 <= _3534;
        133:
            _3905 <= _3537;
        134:
            _3905 <= _3540;
        135:
            _3905 <= _3543;
        136:
            _3905 <= _3546;
        137:
            _3905 <= _3549;
        138:
            _3905 <= _3552;
        139:
            _3905 <= _3555;
        140:
            _3905 <= _3558;
        141:
            _3905 <= _3561;
        142:
            _3905 <= _3564;
        143:
            _3905 <= _3567;
        144:
            _3905 <= _3570;
        145:
            _3905 <= _3573;
        146:
            _3905 <= _3576;
        147:
            _3905 <= _3579;
        148:
            _3905 <= _3582;
        149:
            _3905 <= _3585;
        150:
            _3905 <= _3588;
        151:
            _3905 <= _3591;
        152:
            _3905 <= _3594;
        153:
            _3905 <= _3597;
        154:
            _3905 <= _3600;
        155:
            _3905 <= _3603;
        156:
            _3905 <= _3606;
        157:
            _3905 <= _3609;
        158:
            _3905 <= _3612;
        159:
            _3905 <= _3615;
        160:
            _3905 <= _3618;
        161:
            _3905 <= _3621;
        162:
            _3905 <= _3624;
        163:
            _3905 <= _3627;
        164:
            _3905 <= _3630;
        165:
            _3905 <= _3633;
        166:
            _3905 <= _3636;
        167:
            _3905 <= _3639;
        168:
            _3905 <= _3642;
        169:
            _3905 <= _3645;
        170:
            _3905 <= _3648;
        171:
            _3905 <= _3651;
        172:
            _3905 <= _3654;
        173:
            _3905 <= _3657;
        174:
            _3905 <= _3660;
        175:
            _3905 <= _3663;
        176:
            _3905 <= _3666;
        177:
            _3905 <= _3669;
        178:
            _3905 <= _3672;
        179:
            _3905 <= _3675;
        180:
            _3905 <= _3678;
        181:
            _3905 <= _3681;
        182:
            _3905 <= _3684;
        183:
            _3905 <= _3687;
        184:
            _3905 <= _3690;
        185:
            _3905 <= _3693;
        186:
            _3905 <= _3696;
        187:
            _3905 <= _3699;
        188:
            _3905 <= _3702;
        189:
            _3905 <= _3705;
        190:
            _3905 <= _3708;
        191:
            _3905 <= _3711;
        192:
            _3905 <= _3714;
        193:
            _3905 <= _3717;
        194:
            _3905 <= _3720;
        195:
            _3905 <= _3723;
        196:
            _3905 <= _3726;
        197:
            _3905 <= _3729;
        198:
            _3905 <= _3732;
        199:
            _3905 <= _3735;
        200:
            _3905 <= _3738;
        201:
            _3905 <= _3741;
        202:
            _3905 <= _3744;
        203:
            _3905 <= _3747;
        204:
            _3905 <= _3750;
        205:
            _3905 <= _3753;
        206:
            _3905 <= _3756;
        207:
            _3905 <= _3759;
        208:
            _3905 <= _3762;
        209:
            _3905 <= _3765;
        210:
            _3905 <= _3768;
        211:
            _3905 <= _3771;
        212:
            _3905 <= _3774;
        213:
            _3905 <= _3777;
        214:
            _3905 <= _3780;
        215:
            _3905 <= _3783;
        216:
            _3905 <= _3786;
        217:
            _3905 <= _3789;
        218:
            _3905 <= _3792;
        219:
            _3905 <= _3795;
        220:
            _3905 <= _3798;
        221:
            _3905 <= _3801;
        222:
            _3905 <= _3804;
        223:
            _3905 <= _3807;
        224:
            _3905 <= _3810;
        225:
            _3905 <= _3813;
        226:
            _3905 <= _3816;
        227:
            _3905 <= _3819;
        228:
            _3905 <= _3822;
        229:
            _3905 <= _3825;
        230:
            _3905 <= _3828;
        231:
            _3905 <= _3831;
        232:
            _3905 <= _3834;
        233:
            _3905 <= _3837;
        234:
            _3905 <= _3840;
        235:
            _3905 <= _3843;
        236:
            _3905 <= _3846;
        237:
            _3905 <= _3849;
        238:
            _3905 <= _3852;
        239:
            _3905 <= _3855;
        240:
            _3905 <= _3858;
        241:
            _3905 <= _3861;
        242:
            _3905 <= _3864;
        243:
            _3905 <= _3867;
        244:
            _3905 <= _3870;
        245:
            _3905 <= _3873;
        246:
            _3905 <= _3876;
        247:
            _3905 <= _3879;
        248:
            _3905 <= _3882;
        249:
            _3905 <= _3885;
        250:
            _3905 <= _3888;
        251:
            _3905 <= _3891;
        252:
            _3905 <= _3894;
        253:
            _3905 <= _3897;
        254:
            _3905 <= _3900;
        default:
            _3905 <= _3903;
        endcase
    end
    always @* begin
        case (_3905)
        0:
            _3906 <= _3138;
        1:
            _3906 <= _3141;
        2:
            _3906 <= _3144;
        3:
            _3906 <= _3147;
        4:
            _3906 <= _3150;
        5:
            _3906 <= _3153;
        6:
            _3906 <= _3156;
        7:
            _3906 <= _3159;
        8:
            _3906 <= _3162;
        9:
            _3906 <= _3165;
        10:
            _3906 <= _3168;
        11:
            _3906 <= _3171;
        12:
            _3906 <= _3174;
        13:
            _3906 <= _3177;
        14:
            _3906 <= _3180;
        15:
            _3906 <= _3183;
        16:
            _3906 <= _3186;
        17:
            _3906 <= _3189;
        18:
            _3906 <= _3192;
        19:
            _3906 <= _3195;
        20:
            _3906 <= _3198;
        21:
            _3906 <= _3201;
        22:
            _3906 <= _3204;
        23:
            _3906 <= _3207;
        24:
            _3906 <= _3210;
        25:
            _3906 <= _3213;
        26:
            _3906 <= _3216;
        27:
            _3906 <= _3219;
        28:
            _3906 <= _3222;
        29:
            _3906 <= _3225;
        30:
            _3906 <= _3228;
        31:
            _3906 <= _3231;
        32:
            _3906 <= _3234;
        33:
            _3906 <= _3237;
        34:
            _3906 <= _3240;
        35:
            _3906 <= _3243;
        36:
            _3906 <= _3246;
        37:
            _3906 <= _3249;
        38:
            _3906 <= _3252;
        39:
            _3906 <= _3255;
        40:
            _3906 <= _3258;
        41:
            _3906 <= _3261;
        42:
            _3906 <= _3264;
        43:
            _3906 <= _3267;
        44:
            _3906 <= _3270;
        45:
            _3906 <= _3273;
        46:
            _3906 <= _3276;
        47:
            _3906 <= _3279;
        48:
            _3906 <= _3282;
        49:
            _3906 <= _3285;
        50:
            _3906 <= _3288;
        51:
            _3906 <= _3291;
        52:
            _3906 <= _3294;
        53:
            _3906 <= _3297;
        54:
            _3906 <= _3300;
        55:
            _3906 <= _3303;
        56:
            _3906 <= _3306;
        57:
            _3906 <= _3309;
        58:
            _3906 <= _3312;
        59:
            _3906 <= _3315;
        60:
            _3906 <= _3318;
        61:
            _3906 <= _3321;
        62:
            _3906 <= _3324;
        63:
            _3906 <= _3327;
        64:
            _3906 <= _3330;
        65:
            _3906 <= _3333;
        66:
            _3906 <= _3336;
        67:
            _3906 <= _3339;
        68:
            _3906 <= _3342;
        69:
            _3906 <= _3345;
        70:
            _3906 <= _3348;
        71:
            _3906 <= _3351;
        72:
            _3906 <= _3354;
        73:
            _3906 <= _3357;
        74:
            _3906 <= _3360;
        75:
            _3906 <= _3363;
        76:
            _3906 <= _3366;
        77:
            _3906 <= _3369;
        78:
            _3906 <= _3372;
        79:
            _3906 <= _3375;
        80:
            _3906 <= _3378;
        81:
            _3906 <= _3381;
        82:
            _3906 <= _3384;
        83:
            _3906 <= _3387;
        84:
            _3906 <= _3390;
        85:
            _3906 <= _3393;
        86:
            _3906 <= _3396;
        87:
            _3906 <= _3399;
        88:
            _3906 <= _3402;
        89:
            _3906 <= _3405;
        90:
            _3906 <= _3408;
        91:
            _3906 <= _3411;
        92:
            _3906 <= _3414;
        93:
            _3906 <= _3417;
        94:
            _3906 <= _3420;
        95:
            _3906 <= _3423;
        96:
            _3906 <= _3426;
        97:
            _3906 <= _3429;
        98:
            _3906 <= _3432;
        99:
            _3906 <= _3435;
        100:
            _3906 <= _3438;
        101:
            _3906 <= _3441;
        102:
            _3906 <= _3444;
        103:
            _3906 <= _3447;
        104:
            _3906 <= _3450;
        105:
            _3906 <= _3453;
        106:
            _3906 <= _3456;
        107:
            _3906 <= _3459;
        108:
            _3906 <= _3462;
        109:
            _3906 <= _3465;
        110:
            _3906 <= _3468;
        111:
            _3906 <= _3471;
        112:
            _3906 <= _3474;
        113:
            _3906 <= _3477;
        114:
            _3906 <= _3480;
        115:
            _3906 <= _3483;
        116:
            _3906 <= _3486;
        117:
            _3906 <= _3489;
        118:
            _3906 <= _3492;
        119:
            _3906 <= _3495;
        120:
            _3906 <= _3498;
        121:
            _3906 <= _3501;
        122:
            _3906 <= _3504;
        123:
            _3906 <= _3507;
        124:
            _3906 <= _3510;
        125:
            _3906 <= _3513;
        126:
            _3906 <= _3516;
        127:
            _3906 <= _3519;
        128:
            _3906 <= _3522;
        129:
            _3906 <= _3525;
        130:
            _3906 <= _3528;
        131:
            _3906 <= _3531;
        132:
            _3906 <= _3534;
        133:
            _3906 <= _3537;
        134:
            _3906 <= _3540;
        135:
            _3906 <= _3543;
        136:
            _3906 <= _3546;
        137:
            _3906 <= _3549;
        138:
            _3906 <= _3552;
        139:
            _3906 <= _3555;
        140:
            _3906 <= _3558;
        141:
            _3906 <= _3561;
        142:
            _3906 <= _3564;
        143:
            _3906 <= _3567;
        144:
            _3906 <= _3570;
        145:
            _3906 <= _3573;
        146:
            _3906 <= _3576;
        147:
            _3906 <= _3579;
        148:
            _3906 <= _3582;
        149:
            _3906 <= _3585;
        150:
            _3906 <= _3588;
        151:
            _3906 <= _3591;
        152:
            _3906 <= _3594;
        153:
            _3906 <= _3597;
        154:
            _3906 <= _3600;
        155:
            _3906 <= _3603;
        156:
            _3906 <= _3606;
        157:
            _3906 <= _3609;
        158:
            _3906 <= _3612;
        159:
            _3906 <= _3615;
        160:
            _3906 <= _3618;
        161:
            _3906 <= _3621;
        162:
            _3906 <= _3624;
        163:
            _3906 <= _3627;
        164:
            _3906 <= _3630;
        165:
            _3906 <= _3633;
        166:
            _3906 <= _3636;
        167:
            _3906 <= _3639;
        168:
            _3906 <= _3642;
        169:
            _3906 <= _3645;
        170:
            _3906 <= _3648;
        171:
            _3906 <= _3651;
        172:
            _3906 <= _3654;
        173:
            _3906 <= _3657;
        174:
            _3906 <= _3660;
        175:
            _3906 <= _3663;
        176:
            _3906 <= _3666;
        177:
            _3906 <= _3669;
        178:
            _3906 <= _3672;
        179:
            _3906 <= _3675;
        180:
            _3906 <= _3678;
        181:
            _3906 <= _3681;
        182:
            _3906 <= _3684;
        183:
            _3906 <= _3687;
        184:
            _3906 <= _3690;
        185:
            _3906 <= _3693;
        186:
            _3906 <= _3696;
        187:
            _3906 <= _3699;
        188:
            _3906 <= _3702;
        189:
            _3906 <= _3705;
        190:
            _3906 <= _3708;
        191:
            _3906 <= _3711;
        192:
            _3906 <= _3714;
        193:
            _3906 <= _3717;
        194:
            _3906 <= _3720;
        195:
            _3906 <= _3723;
        196:
            _3906 <= _3726;
        197:
            _3906 <= _3729;
        198:
            _3906 <= _3732;
        199:
            _3906 <= _3735;
        200:
            _3906 <= _3738;
        201:
            _3906 <= _3741;
        202:
            _3906 <= _3744;
        203:
            _3906 <= _3747;
        204:
            _3906 <= _3750;
        205:
            _3906 <= _3753;
        206:
            _3906 <= _3756;
        207:
            _3906 <= _3759;
        208:
            _3906 <= _3762;
        209:
            _3906 <= _3765;
        210:
            _3906 <= _3768;
        211:
            _3906 <= _3771;
        212:
            _3906 <= _3774;
        213:
            _3906 <= _3777;
        214:
            _3906 <= _3780;
        215:
            _3906 <= _3783;
        216:
            _3906 <= _3786;
        217:
            _3906 <= _3789;
        218:
            _3906 <= _3792;
        219:
            _3906 <= _3795;
        220:
            _3906 <= _3798;
        221:
            _3906 <= _3801;
        222:
            _3906 <= _3804;
        223:
            _3906 <= _3807;
        224:
            _3906 <= _3810;
        225:
            _3906 <= _3813;
        226:
            _3906 <= _3816;
        227:
            _3906 <= _3819;
        228:
            _3906 <= _3822;
        229:
            _3906 <= _3825;
        230:
            _3906 <= _3828;
        231:
            _3906 <= _3831;
        232:
            _3906 <= _3834;
        233:
            _3906 <= _3837;
        234:
            _3906 <= _3840;
        235:
            _3906 <= _3843;
        236:
            _3906 <= _3846;
        237:
            _3906 <= _3849;
        238:
            _3906 <= _3852;
        239:
            _3906 <= _3855;
        240:
            _3906 <= _3858;
        241:
            _3906 <= _3861;
        242:
            _3906 <= _3864;
        243:
            _3906 <= _3867;
        244:
            _3906 <= _3870;
        245:
            _3906 <= _3873;
        246:
            _3906 <= _3876;
        247:
            _3906 <= _3879;
        248:
            _3906 <= _3882;
        249:
            _3906 <= _3885;
        250:
            _3906 <= _3888;
        251:
            _3906 <= _3891;
        252:
            _3906 <= _3894;
        253:
            _3906 <= _3897;
        254:
            _3906 <= _3900;
        default:
            _3906 <= _3903;
        endcase
    end
    always @* begin
        case (_3906)
        0:
            _3907 <= _3138;
        1:
            _3907 <= _3141;
        2:
            _3907 <= _3144;
        3:
            _3907 <= _3147;
        4:
            _3907 <= _3150;
        5:
            _3907 <= _3153;
        6:
            _3907 <= _3156;
        7:
            _3907 <= _3159;
        8:
            _3907 <= _3162;
        9:
            _3907 <= _3165;
        10:
            _3907 <= _3168;
        11:
            _3907 <= _3171;
        12:
            _3907 <= _3174;
        13:
            _3907 <= _3177;
        14:
            _3907 <= _3180;
        15:
            _3907 <= _3183;
        16:
            _3907 <= _3186;
        17:
            _3907 <= _3189;
        18:
            _3907 <= _3192;
        19:
            _3907 <= _3195;
        20:
            _3907 <= _3198;
        21:
            _3907 <= _3201;
        22:
            _3907 <= _3204;
        23:
            _3907 <= _3207;
        24:
            _3907 <= _3210;
        25:
            _3907 <= _3213;
        26:
            _3907 <= _3216;
        27:
            _3907 <= _3219;
        28:
            _3907 <= _3222;
        29:
            _3907 <= _3225;
        30:
            _3907 <= _3228;
        31:
            _3907 <= _3231;
        32:
            _3907 <= _3234;
        33:
            _3907 <= _3237;
        34:
            _3907 <= _3240;
        35:
            _3907 <= _3243;
        36:
            _3907 <= _3246;
        37:
            _3907 <= _3249;
        38:
            _3907 <= _3252;
        39:
            _3907 <= _3255;
        40:
            _3907 <= _3258;
        41:
            _3907 <= _3261;
        42:
            _3907 <= _3264;
        43:
            _3907 <= _3267;
        44:
            _3907 <= _3270;
        45:
            _3907 <= _3273;
        46:
            _3907 <= _3276;
        47:
            _3907 <= _3279;
        48:
            _3907 <= _3282;
        49:
            _3907 <= _3285;
        50:
            _3907 <= _3288;
        51:
            _3907 <= _3291;
        52:
            _3907 <= _3294;
        53:
            _3907 <= _3297;
        54:
            _3907 <= _3300;
        55:
            _3907 <= _3303;
        56:
            _3907 <= _3306;
        57:
            _3907 <= _3309;
        58:
            _3907 <= _3312;
        59:
            _3907 <= _3315;
        60:
            _3907 <= _3318;
        61:
            _3907 <= _3321;
        62:
            _3907 <= _3324;
        63:
            _3907 <= _3327;
        64:
            _3907 <= _3330;
        65:
            _3907 <= _3333;
        66:
            _3907 <= _3336;
        67:
            _3907 <= _3339;
        68:
            _3907 <= _3342;
        69:
            _3907 <= _3345;
        70:
            _3907 <= _3348;
        71:
            _3907 <= _3351;
        72:
            _3907 <= _3354;
        73:
            _3907 <= _3357;
        74:
            _3907 <= _3360;
        75:
            _3907 <= _3363;
        76:
            _3907 <= _3366;
        77:
            _3907 <= _3369;
        78:
            _3907 <= _3372;
        79:
            _3907 <= _3375;
        80:
            _3907 <= _3378;
        81:
            _3907 <= _3381;
        82:
            _3907 <= _3384;
        83:
            _3907 <= _3387;
        84:
            _3907 <= _3390;
        85:
            _3907 <= _3393;
        86:
            _3907 <= _3396;
        87:
            _3907 <= _3399;
        88:
            _3907 <= _3402;
        89:
            _3907 <= _3405;
        90:
            _3907 <= _3408;
        91:
            _3907 <= _3411;
        92:
            _3907 <= _3414;
        93:
            _3907 <= _3417;
        94:
            _3907 <= _3420;
        95:
            _3907 <= _3423;
        96:
            _3907 <= _3426;
        97:
            _3907 <= _3429;
        98:
            _3907 <= _3432;
        99:
            _3907 <= _3435;
        100:
            _3907 <= _3438;
        101:
            _3907 <= _3441;
        102:
            _3907 <= _3444;
        103:
            _3907 <= _3447;
        104:
            _3907 <= _3450;
        105:
            _3907 <= _3453;
        106:
            _3907 <= _3456;
        107:
            _3907 <= _3459;
        108:
            _3907 <= _3462;
        109:
            _3907 <= _3465;
        110:
            _3907 <= _3468;
        111:
            _3907 <= _3471;
        112:
            _3907 <= _3474;
        113:
            _3907 <= _3477;
        114:
            _3907 <= _3480;
        115:
            _3907 <= _3483;
        116:
            _3907 <= _3486;
        117:
            _3907 <= _3489;
        118:
            _3907 <= _3492;
        119:
            _3907 <= _3495;
        120:
            _3907 <= _3498;
        121:
            _3907 <= _3501;
        122:
            _3907 <= _3504;
        123:
            _3907 <= _3507;
        124:
            _3907 <= _3510;
        125:
            _3907 <= _3513;
        126:
            _3907 <= _3516;
        127:
            _3907 <= _3519;
        128:
            _3907 <= _3522;
        129:
            _3907 <= _3525;
        130:
            _3907 <= _3528;
        131:
            _3907 <= _3531;
        132:
            _3907 <= _3534;
        133:
            _3907 <= _3537;
        134:
            _3907 <= _3540;
        135:
            _3907 <= _3543;
        136:
            _3907 <= _3546;
        137:
            _3907 <= _3549;
        138:
            _3907 <= _3552;
        139:
            _3907 <= _3555;
        140:
            _3907 <= _3558;
        141:
            _3907 <= _3561;
        142:
            _3907 <= _3564;
        143:
            _3907 <= _3567;
        144:
            _3907 <= _3570;
        145:
            _3907 <= _3573;
        146:
            _3907 <= _3576;
        147:
            _3907 <= _3579;
        148:
            _3907 <= _3582;
        149:
            _3907 <= _3585;
        150:
            _3907 <= _3588;
        151:
            _3907 <= _3591;
        152:
            _3907 <= _3594;
        153:
            _3907 <= _3597;
        154:
            _3907 <= _3600;
        155:
            _3907 <= _3603;
        156:
            _3907 <= _3606;
        157:
            _3907 <= _3609;
        158:
            _3907 <= _3612;
        159:
            _3907 <= _3615;
        160:
            _3907 <= _3618;
        161:
            _3907 <= _3621;
        162:
            _3907 <= _3624;
        163:
            _3907 <= _3627;
        164:
            _3907 <= _3630;
        165:
            _3907 <= _3633;
        166:
            _3907 <= _3636;
        167:
            _3907 <= _3639;
        168:
            _3907 <= _3642;
        169:
            _3907 <= _3645;
        170:
            _3907 <= _3648;
        171:
            _3907 <= _3651;
        172:
            _3907 <= _3654;
        173:
            _3907 <= _3657;
        174:
            _3907 <= _3660;
        175:
            _3907 <= _3663;
        176:
            _3907 <= _3666;
        177:
            _3907 <= _3669;
        178:
            _3907 <= _3672;
        179:
            _3907 <= _3675;
        180:
            _3907 <= _3678;
        181:
            _3907 <= _3681;
        182:
            _3907 <= _3684;
        183:
            _3907 <= _3687;
        184:
            _3907 <= _3690;
        185:
            _3907 <= _3693;
        186:
            _3907 <= _3696;
        187:
            _3907 <= _3699;
        188:
            _3907 <= _3702;
        189:
            _3907 <= _3705;
        190:
            _3907 <= _3708;
        191:
            _3907 <= _3711;
        192:
            _3907 <= _3714;
        193:
            _3907 <= _3717;
        194:
            _3907 <= _3720;
        195:
            _3907 <= _3723;
        196:
            _3907 <= _3726;
        197:
            _3907 <= _3729;
        198:
            _3907 <= _3732;
        199:
            _3907 <= _3735;
        200:
            _3907 <= _3738;
        201:
            _3907 <= _3741;
        202:
            _3907 <= _3744;
        203:
            _3907 <= _3747;
        204:
            _3907 <= _3750;
        205:
            _3907 <= _3753;
        206:
            _3907 <= _3756;
        207:
            _3907 <= _3759;
        208:
            _3907 <= _3762;
        209:
            _3907 <= _3765;
        210:
            _3907 <= _3768;
        211:
            _3907 <= _3771;
        212:
            _3907 <= _3774;
        213:
            _3907 <= _3777;
        214:
            _3907 <= _3780;
        215:
            _3907 <= _3783;
        216:
            _3907 <= _3786;
        217:
            _3907 <= _3789;
        218:
            _3907 <= _3792;
        219:
            _3907 <= _3795;
        220:
            _3907 <= _3798;
        221:
            _3907 <= _3801;
        222:
            _3907 <= _3804;
        223:
            _3907 <= _3807;
        224:
            _3907 <= _3810;
        225:
            _3907 <= _3813;
        226:
            _3907 <= _3816;
        227:
            _3907 <= _3819;
        228:
            _3907 <= _3822;
        229:
            _3907 <= _3825;
        230:
            _3907 <= _3828;
        231:
            _3907 <= _3831;
        232:
            _3907 <= _3834;
        233:
            _3907 <= _3837;
        234:
            _3907 <= _3840;
        235:
            _3907 <= _3843;
        236:
            _3907 <= _3846;
        237:
            _3907 <= _3849;
        238:
            _3907 <= _3852;
        239:
            _3907 <= _3855;
        240:
            _3907 <= _3858;
        241:
            _3907 <= _3861;
        242:
            _3907 <= _3864;
        243:
            _3907 <= _3867;
        244:
            _3907 <= _3870;
        245:
            _3907 <= _3873;
        246:
            _3907 <= _3876;
        247:
            _3907 <= _3879;
        248:
            _3907 <= _3882;
        249:
            _3907 <= _3885;
        250:
            _3907 <= _3888;
        251:
            _3907 <= _3891;
        252:
            _3907 <= _3894;
        253:
            _3907 <= _3897;
        254:
            _3907 <= _3900;
        default:
            _3907 <= _3903;
        endcase
    end
    always @* begin
        case (_3907)
        0:
            _3908 <= _3138;
        1:
            _3908 <= _3141;
        2:
            _3908 <= _3144;
        3:
            _3908 <= _3147;
        4:
            _3908 <= _3150;
        5:
            _3908 <= _3153;
        6:
            _3908 <= _3156;
        7:
            _3908 <= _3159;
        8:
            _3908 <= _3162;
        9:
            _3908 <= _3165;
        10:
            _3908 <= _3168;
        11:
            _3908 <= _3171;
        12:
            _3908 <= _3174;
        13:
            _3908 <= _3177;
        14:
            _3908 <= _3180;
        15:
            _3908 <= _3183;
        16:
            _3908 <= _3186;
        17:
            _3908 <= _3189;
        18:
            _3908 <= _3192;
        19:
            _3908 <= _3195;
        20:
            _3908 <= _3198;
        21:
            _3908 <= _3201;
        22:
            _3908 <= _3204;
        23:
            _3908 <= _3207;
        24:
            _3908 <= _3210;
        25:
            _3908 <= _3213;
        26:
            _3908 <= _3216;
        27:
            _3908 <= _3219;
        28:
            _3908 <= _3222;
        29:
            _3908 <= _3225;
        30:
            _3908 <= _3228;
        31:
            _3908 <= _3231;
        32:
            _3908 <= _3234;
        33:
            _3908 <= _3237;
        34:
            _3908 <= _3240;
        35:
            _3908 <= _3243;
        36:
            _3908 <= _3246;
        37:
            _3908 <= _3249;
        38:
            _3908 <= _3252;
        39:
            _3908 <= _3255;
        40:
            _3908 <= _3258;
        41:
            _3908 <= _3261;
        42:
            _3908 <= _3264;
        43:
            _3908 <= _3267;
        44:
            _3908 <= _3270;
        45:
            _3908 <= _3273;
        46:
            _3908 <= _3276;
        47:
            _3908 <= _3279;
        48:
            _3908 <= _3282;
        49:
            _3908 <= _3285;
        50:
            _3908 <= _3288;
        51:
            _3908 <= _3291;
        52:
            _3908 <= _3294;
        53:
            _3908 <= _3297;
        54:
            _3908 <= _3300;
        55:
            _3908 <= _3303;
        56:
            _3908 <= _3306;
        57:
            _3908 <= _3309;
        58:
            _3908 <= _3312;
        59:
            _3908 <= _3315;
        60:
            _3908 <= _3318;
        61:
            _3908 <= _3321;
        62:
            _3908 <= _3324;
        63:
            _3908 <= _3327;
        64:
            _3908 <= _3330;
        65:
            _3908 <= _3333;
        66:
            _3908 <= _3336;
        67:
            _3908 <= _3339;
        68:
            _3908 <= _3342;
        69:
            _3908 <= _3345;
        70:
            _3908 <= _3348;
        71:
            _3908 <= _3351;
        72:
            _3908 <= _3354;
        73:
            _3908 <= _3357;
        74:
            _3908 <= _3360;
        75:
            _3908 <= _3363;
        76:
            _3908 <= _3366;
        77:
            _3908 <= _3369;
        78:
            _3908 <= _3372;
        79:
            _3908 <= _3375;
        80:
            _3908 <= _3378;
        81:
            _3908 <= _3381;
        82:
            _3908 <= _3384;
        83:
            _3908 <= _3387;
        84:
            _3908 <= _3390;
        85:
            _3908 <= _3393;
        86:
            _3908 <= _3396;
        87:
            _3908 <= _3399;
        88:
            _3908 <= _3402;
        89:
            _3908 <= _3405;
        90:
            _3908 <= _3408;
        91:
            _3908 <= _3411;
        92:
            _3908 <= _3414;
        93:
            _3908 <= _3417;
        94:
            _3908 <= _3420;
        95:
            _3908 <= _3423;
        96:
            _3908 <= _3426;
        97:
            _3908 <= _3429;
        98:
            _3908 <= _3432;
        99:
            _3908 <= _3435;
        100:
            _3908 <= _3438;
        101:
            _3908 <= _3441;
        102:
            _3908 <= _3444;
        103:
            _3908 <= _3447;
        104:
            _3908 <= _3450;
        105:
            _3908 <= _3453;
        106:
            _3908 <= _3456;
        107:
            _3908 <= _3459;
        108:
            _3908 <= _3462;
        109:
            _3908 <= _3465;
        110:
            _3908 <= _3468;
        111:
            _3908 <= _3471;
        112:
            _3908 <= _3474;
        113:
            _3908 <= _3477;
        114:
            _3908 <= _3480;
        115:
            _3908 <= _3483;
        116:
            _3908 <= _3486;
        117:
            _3908 <= _3489;
        118:
            _3908 <= _3492;
        119:
            _3908 <= _3495;
        120:
            _3908 <= _3498;
        121:
            _3908 <= _3501;
        122:
            _3908 <= _3504;
        123:
            _3908 <= _3507;
        124:
            _3908 <= _3510;
        125:
            _3908 <= _3513;
        126:
            _3908 <= _3516;
        127:
            _3908 <= _3519;
        128:
            _3908 <= _3522;
        129:
            _3908 <= _3525;
        130:
            _3908 <= _3528;
        131:
            _3908 <= _3531;
        132:
            _3908 <= _3534;
        133:
            _3908 <= _3537;
        134:
            _3908 <= _3540;
        135:
            _3908 <= _3543;
        136:
            _3908 <= _3546;
        137:
            _3908 <= _3549;
        138:
            _3908 <= _3552;
        139:
            _3908 <= _3555;
        140:
            _3908 <= _3558;
        141:
            _3908 <= _3561;
        142:
            _3908 <= _3564;
        143:
            _3908 <= _3567;
        144:
            _3908 <= _3570;
        145:
            _3908 <= _3573;
        146:
            _3908 <= _3576;
        147:
            _3908 <= _3579;
        148:
            _3908 <= _3582;
        149:
            _3908 <= _3585;
        150:
            _3908 <= _3588;
        151:
            _3908 <= _3591;
        152:
            _3908 <= _3594;
        153:
            _3908 <= _3597;
        154:
            _3908 <= _3600;
        155:
            _3908 <= _3603;
        156:
            _3908 <= _3606;
        157:
            _3908 <= _3609;
        158:
            _3908 <= _3612;
        159:
            _3908 <= _3615;
        160:
            _3908 <= _3618;
        161:
            _3908 <= _3621;
        162:
            _3908 <= _3624;
        163:
            _3908 <= _3627;
        164:
            _3908 <= _3630;
        165:
            _3908 <= _3633;
        166:
            _3908 <= _3636;
        167:
            _3908 <= _3639;
        168:
            _3908 <= _3642;
        169:
            _3908 <= _3645;
        170:
            _3908 <= _3648;
        171:
            _3908 <= _3651;
        172:
            _3908 <= _3654;
        173:
            _3908 <= _3657;
        174:
            _3908 <= _3660;
        175:
            _3908 <= _3663;
        176:
            _3908 <= _3666;
        177:
            _3908 <= _3669;
        178:
            _3908 <= _3672;
        179:
            _3908 <= _3675;
        180:
            _3908 <= _3678;
        181:
            _3908 <= _3681;
        182:
            _3908 <= _3684;
        183:
            _3908 <= _3687;
        184:
            _3908 <= _3690;
        185:
            _3908 <= _3693;
        186:
            _3908 <= _3696;
        187:
            _3908 <= _3699;
        188:
            _3908 <= _3702;
        189:
            _3908 <= _3705;
        190:
            _3908 <= _3708;
        191:
            _3908 <= _3711;
        192:
            _3908 <= _3714;
        193:
            _3908 <= _3717;
        194:
            _3908 <= _3720;
        195:
            _3908 <= _3723;
        196:
            _3908 <= _3726;
        197:
            _3908 <= _3729;
        198:
            _3908 <= _3732;
        199:
            _3908 <= _3735;
        200:
            _3908 <= _3738;
        201:
            _3908 <= _3741;
        202:
            _3908 <= _3744;
        203:
            _3908 <= _3747;
        204:
            _3908 <= _3750;
        205:
            _3908 <= _3753;
        206:
            _3908 <= _3756;
        207:
            _3908 <= _3759;
        208:
            _3908 <= _3762;
        209:
            _3908 <= _3765;
        210:
            _3908 <= _3768;
        211:
            _3908 <= _3771;
        212:
            _3908 <= _3774;
        213:
            _3908 <= _3777;
        214:
            _3908 <= _3780;
        215:
            _3908 <= _3783;
        216:
            _3908 <= _3786;
        217:
            _3908 <= _3789;
        218:
            _3908 <= _3792;
        219:
            _3908 <= _3795;
        220:
            _3908 <= _3798;
        221:
            _3908 <= _3801;
        222:
            _3908 <= _3804;
        223:
            _3908 <= _3807;
        224:
            _3908 <= _3810;
        225:
            _3908 <= _3813;
        226:
            _3908 <= _3816;
        227:
            _3908 <= _3819;
        228:
            _3908 <= _3822;
        229:
            _3908 <= _3825;
        230:
            _3908 <= _3828;
        231:
            _3908 <= _3831;
        232:
            _3908 <= _3834;
        233:
            _3908 <= _3837;
        234:
            _3908 <= _3840;
        235:
            _3908 <= _3843;
        236:
            _3908 <= _3846;
        237:
            _3908 <= _3849;
        238:
            _3908 <= _3852;
        239:
            _3908 <= _3855;
        240:
            _3908 <= _3858;
        241:
            _3908 <= _3861;
        242:
            _3908 <= _3864;
        243:
            _3908 <= _3867;
        244:
            _3908 <= _3870;
        245:
            _3908 <= _3873;
        246:
            _3908 <= _3876;
        247:
            _3908 <= _3879;
        248:
            _3908 <= _3882;
        249:
            _3908 <= _3885;
        250:
            _3908 <= _3888;
        251:
            _3908 <= _3891;
        252:
            _3908 <= _3894;
        253:
            _3908 <= _3897;
        254:
            _3908 <= _3900;
        default:
            _3908 <= _3903;
        endcase
    end
    always @* begin
        case (_3908)
        0:
            _3909 <= _3138;
        1:
            _3909 <= _3141;
        2:
            _3909 <= _3144;
        3:
            _3909 <= _3147;
        4:
            _3909 <= _3150;
        5:
            _3909 <= _3153;
        6:
            _3909 <= _3156;
        7:
            _3909 <= _3159;
        8:
            _3909 <= _3162;
        9:
            _3909 <= _3165;
        10:
            _3909 <= _3168;
        11:
            _3909 <= _3171;
        12:
            _3909 <= _3174;
        13:
            _3909 <= _3177;
        14:
            _3909 <= _3180;
        15:
            _3909 <= _3183;
        16:
            _3909 <= _3186;
        17:
            _3909 <= _3189;
        18:
            _3909 <= _3192;
        19:
            _3909 <= _3195;
        20:
            _3909 <= _3198;
        21:
            _3909 <= _3201;
        22:
            _3909 <= _3204;
        23:
            _3909 <= _3207;
        24:
            _3909 <= _3210;
        25:
            _3909 <= _3213;
        26:
            _3909 <= _3216;
        27:
            _3909 <= _3219;
        28:
            _3909 <= _3222;
        29:
            _3909 <= _3225;
        30:
            _3909 <= _3228;
        31:
            _3909 <= _3231;
        32:
            _3909 <= _3234;
        33:
            _3909 <= _3237;
        34:
            _3909 <= _3240;
        35:
            _3909 <= _3243;
        36:
            _3909 <= _3246;
        37:
            _3909 <= _3249;
        38:
            _3909 <= _3252;
        39:
            _3909 <= _3255;
        40:
            _3909 <= _3258;
        41:
            _3909 <= _3261;
        42:
            _3909 <= _3264;
        43:
            _3909 <= _3267;
        44:
            _3909 <= _3270;
        45:
            _3909 <= _3273;
        46:
            _3909 <= _3276;
        47:
            _3909 <= _3279;
        48:
            _3909 <= _3282;
        49:
            _3909 <= _3285;
        50:
            _3909 <= _3288;
        51:
            _3909 <= _3291;
        52:
            _3909 <= _3294;
        53:
            _3909 <= _3297;
        54:
            _3909 <= _3300;
        55:
            _3909 <= _3303;
        56:
            _3909 <= _3306;
        57:
            _3909 <= _3309;
        58:
            _3909 <= _3312;
        59:
            _3909 <= _3315;
        60:
            _3909 <= _3318;
        61:
            _3909 <= _3321;
        62:
            _3909 <= _3324;
        63:
            _3909 <= _3327;
        64:
            _3909 <= _3330;
        65:
            _3909 <= _3333;
        66:
            _3909 <= _3336;
        67:
            _3909 <= _3339;
        68:
            _3909 <= _3342;
        69:
            _3909 <= _3345;
        70:
            _3909 <= _3348;
        71:
            _3909 <= _3351;
        72:
            _3909 <= _3354;
        73:
            _3909 <= _3357;
        74:
            _3909 <= _3360;
        75:
            _3909 <= _3363;
        76:
            _3909 <= _3366;
        77:
            _3909 <= _3369;
        78:
            _3909 <= _3372;
        79:
            _3909 <= _3375;
        80:
            _3909 <= _3378;
        81:
            _3909 <= _3381;
        82:
            _3909 <= _3384;
        83:
            _3909 <= _3387;
        84:
            _3909 <= _3390;
        85:
            _3909 <= _3393;
        86:
            _3909 <= _3396;
        87:
            _3909 <= _3399;
        88:
            _3909 <= _3402;
        89:
            _3909 <= _3405;
        90:
            _3909 <= _3408;
        91:
            _3909 <= _3411;
        92:
            _3909 <= _3414;
        93:
            _3909 <= _3417;
        94:
            _3909 <= _3420;
        95:
            _3909 <= _3423;
        96:
            _3909 <= _3426;
        97:
            _3909 <= _3429;
        98:
            _3909 <= _3432;
        99:
            _3909 <= _3435;
        100:
            _3909 <= _3438;
        101:
            _3909 <= _3441;
        102:
            _3909 <= _3444;
        103:
            _3909 <= _3447;
        104:
            _3909 <= _3450;
        105:
            _3909 <= _3453;
        106:
            _3909 <= _3456;
        107:
            _3909 <= _3459;
        108:
            _3909 <= _3462;
        109:
            _3909 <= _3465;
        110:
            _3909 <= _3468;
        111:
            _3909 <= _3471;
        112:
            _3909 <= _3474;
        113:
            _3909 <= _3477;
        114:
            _3909 <= _3480;
        115:
            _3909 <= _3483;
        116:
            _3909 <= _3486;
        117:
            _3909 <= _3489;
        118:
            _3909 <= _3492;
        119:
            _3909 <= _3495;
        120:
            _3909 <= _3498;
        121:
            _3909 <= _3501;
        122:
            _3909 <= _3504;
        123:
            _3909 <= _3507;
        124:
            _3909 <= _3510;
        125:
            _3909 <= _3513;
        126:
            _3909 <= _3516;
        127:
            _3909 <= _3519;
        128:
            _3909 <= _3522;
        129:
            _3909 <= _3525;
        130:
            _3909 <= _3528;
        131:
            _3909 <= _3531;
        132:
            _3909 <= _3534;
        133:
            _3909 <= _3537;
        134:
            _3909 <= _3540;
        135:
            _3909 <= _3543;
        136:
            _3909 <= _3546;
        137:
            _3909 <= _3549;
        138:
            _3909 <= _3552;
        139:
            _3909 <= _3555;
        140:
            _3909 <= _3558;
        141:
            _3909 <= _3561;
        142:
            _3909 <= _3564;
        143:
            _3909 <= _3567;
        144:
            _3909 <= _3570;
        145:
            _3909 <= _3573;
        146:
            _3909 <= _3576;
        147:
            _3909 <= _3579;
        148:
            _3909 <= _3582;
        149:
            _3909 <= _3585;
        150:
            _3909 <= _3588;
        151:
            _3909 <= _3591;
        152:
            _3909 <= _3594;
        153:
            _3909 <= _3597;
        154:
            _3909 <= _3600;
        155:
            _3909 <= _3603;
        156:
            _3909 <= _3606;
        157:
            _3909 <= _3609;
        158:
            _3909 <= _3612;
        159:
            _3909 <= _3615;
        160:
            _3909 <= _3618;
        161:
            _3909 <= _3621;
        162:
            _3909 <= _3624;
        163:
            _3909 <= _3627;
        164:
            _3909 <= _3630;
        165:
            _3909 <= _3633;
        166:
            _3909 <= _3636;
        167:
            _3909 <= _3639;
        168:
            _3909 <= _3642;
        169:
            _3909 <= _3645;
        170:
            _3909 <= _3648;
        171:
            _3909 <= _3651;
        172:
            _3909 <= _3654;
        173:
            _3909 <= _3657;
        174:
            _3909 <= _3660;
        175:
            _3909 <= _3663;
        176:
            _3909 <= _3666;
        177:
            _3909 <= _3669;
        178:
            _3909 <= _3672;
        179:
            _3909 <= _3675;
        180:
            _3909 <= _3678;
        181:
            _3909 <= _3681;
        182:
            _3909 <= _3684;
        183:
            _3909 <= _3687;
        184:
            _3909 <= _3690;
        185:
            _3909 <= _3693;
        186:
            _3909 <= _3696;
        187:
            _3909 <= _3699;
        188:
            _3909 <= _3702;
        189:
            _3909 <= _3705;
        190:
            _3909 <= _3708;
        191:
            _3909 <= _3711;
        192:
            _3909 <= _3714;
        193:
            _3909 <= _3717;
        194:
            _3909 <= _3720;
        195:
            _3909 <= _3723;
        196:
            _3909 <= _3726;
        197:
            _3909 <= _3729;
        198:
            _3909 <= _3732;
        199:
            _3909 <= _3735;
        200:
            _3909 <= _3738;
        201:
            _3909 <= _3741;
        202:
            _3909 <= _3744;
        203:
            _3909 <= _3747;
        204:
            _3909 <= _3750;
        205:
            _3909 <= _3753;
        206:
            _3909 <= _3756;
        207:
            _3909 <= _3759;
        208:
            _3909 <= _3762;
        209:
            _3909 <= _3765;
        210:
            _3909 <= _3768;
        211:
            _3909 <= _3771;
        212:
            _3909 <= _3774;
        213:
            _3909 <= _3777;
        214:
            _3909 <= _3780;
        215:
            _3909 <= _3783;
        216:
            _3909 <= _3786;
        217:
            _3909 <= _3789;
        218:
            _3909 <= _3792;
        219:
            _3909 <= _3795;
        220:
            _3909 <= _3798;
        221:
            _3909 <= _3801;
        222:
            _3909 <= _3804;
        223:
            _3909 <= _3807;
        224:
            _3909 <= _3810;
        225:
            _3909 <= _3813;
        226:
            _3909 <= _3816;
        227:
            _3909 <= _3819;
        228:
            _3909 <= _3822;
        229:
            _3909 <= _3825;
        230:
            _3909 <= _3828;
        231:
            _3909 <= _3831;
        232:
            _3909 <= _3834;
        233:
            _3909 <= _3837;
        234:
            _3909 <= _3840;
        235:
            _3909 <= _3843;
        236:
            _3909 <= _3846;
        237:
            _3909 <= _3849;
        238:
            _3909 <= _3852;
        239:
            _3909 <= _3855;
        240:
            _3909 <= _3858;
        241:
            _3909 <= _3861;
        242:
            _3909 <= _3864;
        243:
            _3909 <= _3867;
        244:
            _3909 <= _3870;
        245:
            _3909 <= _3873;
        246:
            _3909 <= _3876;
        247:
            _3909 <= _3879;
        248:
            _3909 <= _3882;
        249:
            _3909 <= _3885;
        250:
            _3909 <= _3888;
        251:
            _3909 <= _3891;
        252:
            _3909 <= _3894;
        253:
            _3909 <= _3897;
        254:
            _3909 <= _3900;
        default:
            _3909 <= _3903;
        endcase
    end
    always @* begin
        case (_3909)
        0:
            _3910 <= _3138;
        1:
            _3910 <= _3141;
        2:
            _3910 <= _3144;
        3:
            _3910 <= _3147;
        4:
            _3910 <= _3150;
        5:
            _3910 <= _3153;
        6:
            _3910 <= _3156;
        7:
            _3910 <= _3159;
        8:
            _3910 <= _3162;
        9:
            _3910 <= _3165;
        10:
            _3910 <= _3168;
        11:
            _3910 <= _3171;
        12:
            _3910 <= _3174;
        13:
            _3910 <= _3177;
        14:
            _3910 <= _3180;
        15:
            _3910 <= _3183;
        16:
            _3910 <= _3186;
        17:
            _3910 <= _3189;
        18:
            _3910 <= _3192;
        19:
            _3910 <= _3195;
        20:
            _3910 <= _3198;
        21:
            _3910 <= _3201;
        22:
            _3910 <= _3204;
        23:
            _3910 <= _3207;
        24:
            _3910 <= _3210;
        25:
            _3910 <= _3213;
        26:
            _3910 <= _3216;
        27:
            _3910 <= _3219;
        28:
            _3910 <= _3222;
        29:
            _3910 <= _3225;
        30:
            _3910 <= _3228;
        31:
            _3910 <= _3231;
        32:
            _3910 <= _3234;
        33:
            _3910 <= _3237;
        34:
            _3910 <= _3240;
        35:
            _3910 <= _3243;
        36:
            _3910 <= _3246;
        37:
            _3910 <= _3249;
        38:
            _3910 <= _3252;
        39:
            _3910 <= _3255;
        40:
            _3910 <= _3258;
        41:
            _3910 <= _3261;
        42:
            _3910 <= _3264;
        43:
            _3910 <= _3267;
        44:
            _3910 <= _3270;
        45:
            _3910 <= _3273;
        46:
            _3910 <= _3276;
        47:
            _3910 <= _3279;
        48:
            _3910 <= _3282;
        49:
            _3910 <= _3285;
        50:
            _3910 <= _3288;
        51:
            _3910 <= _3291;
        52:
            _3910 <= _3294;
        53:
            _3910 <= _3297;
        54:
            _3910 <= _3300;
        55:
            _3910 <= _3303;
        56:
            _3910 <= _3306;
        57:
            _3910 <= _3309;
        58:
            _3910 <= _3312;
        59:
            _3910 <= _3315;
        60:
            _3910 <= _3318;
        61:
            _3910 <= _3321;
        62:
            _3910 <= _3324;
        63:
            _3910 <= _3327;
        64:
            _3910 <= _3330;
        65:
            _3910 <= _3333;
        66:
            _3910 <= _3336;
        67:
            _3910 <= _3339;
        68:
            _3910 <= _3342;
        69:
            _3910 <= _3345;
        70:
            _3910 <= _3348;
        71:
            _3910 <= _3351;
        72:
            _3910 <= _3354;
        73:
            _3910 <= _3357;
        74:
            _3910 <= _3360;
        75:
            _3910 <= _3363;
        76:
            _3910 <= _3366;
        77:
            _3910 <= _3369;
        78:
            _3910 <= _3372;
        79:
            _3910 <= _3375;
        80:
            _3910 <= _3378;
        81:
            _3910 <= _3381;
        82:
            _3910 <= _3384;
        83:
            _3910 <= _3387;
        84:
            _3910 <= _3390;
        85:
            _3910 <= _3393;
        86:
            _3910 <= _3396;
        87:
            _3910 <= _3399;
        88:
            _3910 <= _3402;
        89:
            _3910 <= _3405;
        90:
            _3910 <= _3408;
        91:
            _3910 <= _3411;
        92:
            _3910 <= _3414;
        93:
            _3910 <= _3417;
        94:
            _3910 <= _3420;
        95:
            _3910 <= _3423;
        96:
            _3910 <= _3426;
        97:
            _3910 <= _3429;
        98:
            _3910 <= _3432;
        99:
            _3910 <= _3435;
        100:
            _3910 <= _3438;
        101:
            _3910 <= _3441;
        102:
            _3910 <= _3444;
        103:
            _3910 <= _3447;
        104:
            _3910 <= _3450;
        105:
            _3910 <= _3453;
        106:
            _3910 <= _3456;
        107:
            _3910 <= _3459;
        108:
            _3910 <= _3462;
        109:
            _3910 <= _3465;
        110:
            _3910 <= _3468;
        111:
            _3910 <= _3471;
        112:
            _3910 <= _3474;
        113:
            _3910 <= _3477;
        114:
            _3910 <= _3480;
        115:
            _3910 <= _3483;
        116:
            _3910 <= _3486;
        117:
            _3910 <= _3489;
        118:
            _3910 <= _3492;
        119:
            _3910 <= _3495;
        120:
            _3910 <= _3498;
        121:
            _3910 <= _3501;
        122:
            _3910 <= _3504;
        123:
            _3910 <= _3507;
        124:
            _3910 <= _3510;
        125:
            _3910 <= _3513;
        126:
            _3910 <= _3516;
        127:
            _3910 <= _3519;
        128:
            _3910 <= _3522;
        129:
            _3910 <= _3525;
        130:
            _3910 <= _3528;
        131:
            _3910 <= _3531;
        132:
            _3910 <= _3534;
        133:
            _3910 <= _3537;
        134:
            _3910 <= _3540;
        135:
            _3910 <= _3543;
        136:
            _3910 <= _3546;
        137:
            _3910 <= _3549;
        138:
            _3910 <= _3552;
        139:
            _3910 <= _3555;
        140:
            _3910 <= _3558;
        141:
            _3910 <= _3561;
        142:
            _3910 <= _3564;
        143:
            _3910 <= _3567;
        144:
            _3910 <= _3570;
        145:
            _3910 <= _3573;
        146:
            _3910 <= _3576;
        147:
            _3910 <= _3579;
        148:
            _3910 <= _3582;
        149:
            _3910 <= _3585;
        150:
            _3910 <= _3588;
        151:
            _3910 <= _3591;
        152:
            _3910 <= _3594;
        153:
            _3910 <= _3597;
        154:
            _3910 <= _3600;
        155:
            _3910 <= _3603;
        156:
            _3910 <= _3606;
        157:
            _3910 <= _3609;
        158:
            _3910 <= _3612;
        159:
            _3910 <= _3615;
        160:
            _3910 <= _3618;
        161:
            _3910 <= _3621;
        162:
            _3910 <= _3624;
        163:
            _3910 <= _3627;
        164:
            _3910 <= _3630;
        165:
            _3910 <= _3633;
        166:
            _3910 <= _3636;
        167:
            _3910 <= _3639;
        168:
            _3910 <= _3642;
        169:
            _3910 <= _3645;
        170:
            _3910 <= _3648;
        171:
            _3910 <= _3651;
        172:
            _3910 <= _3654;
        173:
            _3910 <= _3657;
        174:
            _3910 <= _3660;
        175:
            _3910 <= _3663;
        176:
            _3910 <= _3666;
        177:
            _3910 <= _3669;
        178:
            _3910 <= _3672;
        179:
            _3910 <= _3675;
        180:
            _3910 <= _3678;
        181:
            _3910 <= _3681;
        182:
            _3910 <= _3684;
        183:
            _3910 <= _3687;
        184:
            _3910 <= _3690;
        185:
            _3910 <= _3693;
        186:
            _3910 <= _3696;
        187:
            _3910 <= _3699;
        188:
            _3910 <= _3702;
        189:
            _3910 <= _3705;
        190:
            _3910 <= _3708;
        191:
            _3910 <= _3711;
        192:
            _3910 <= _3714;
        193:
            _3910 <= _3717;
        194:
            _3910 <= _3720;
        195:
            _3910 <= _3723;
        196:
            _3910 <= _3726;
        197:
            _3910 <= _3729;
        198:
            _3910 <= _3732;
        199:
            _3910 <= _3735;
        200:
            _3910 <= _3738;
        201:
            _3910 <= _3741;
        202:
            _3910 <= _3744;
        203:
            _3910 <= _3747;
        204:
            _3910 <= _3750;
        205:
            _3910 <= _3753;
        206:
            _3910 <= _3756;
        207:
            _3910 <= _3759;
        208:
            _3910 <= _3762;
        209:
            _3910 <= _3765;
        210:
            _3910 <= _3768;
        211:
            _3910 <= _3771;
        212:
            _3910 <= _3774;
        213:
            _3910 <= _3777;
        214:
            _3910 <= _3780;
        215:
            _3910 <= _3783;
        216:
            _3910 <= _3786;
        217:
            _3910 <= _3789;
        218:
            _3910 <= _3792;
        219:
            _3910 <= _3795;
        220:
            _3910 <= _3798;
        221:
            _3910 <= _3801;
        222:
            _3910 <= _3804;
        223:
            _3910 <= _3807;
        224:
            _3910 <= _3810;
        225:
            _3910 <= _3813;
        226:
            _3910 <= _3816;
        227:
            _3910 <= _3819;
        228:
            _3910 <= _3822;
        229:
            _3910 <= _3825;
        230:
            _3910 <= _3828;
        231:
            _3910 <= _3831;
        232:
            _3910 <= _3834;
        233:
            _3910 <= _3837;
        234:
            _3910 <= _3840;
        235:
            _3910 <= _3843;
        236:
            _3910 <= _3846;
        237:
            _3910 <= _3849;
        238:
            _3910 <= _3852;
        239:
            _3910 <= _3855;
        240:
            _3910 <= _3858;
        241:
            _3910 <= _3861;
        242:
            _3910 <= _3864;
        243:
            _3910 <= _3867;
        244:
            _3910 <= _3870;
        245:
            _3910 <= _3873;
        246:
            _3910 <= _3876;
        247:
            _3910 <= _3879;
        248:
            _3910 <= _3882;
        249:
            _3910 <= _3885;
        250:
            _3910 <= _3888;
        251:
            _3910 <= _3891;
        252:
            _3910 <= _3894;
        253:
            _3910 <= _3897;
        254:
            _3910 <= _3900;
        default:
            _3910 <= _3903;
        endcase
    end
    always @* begin
        case (_3910)
        0:
            _3911 <= _3138;
        1:
            _3911 <= _3141;
        2:
            _3911 <= _3144;
        3:
            _3911 <= _3147;
        4:
            _3911 <= _3150;
        5:
            _3911 <= _3153;
        6:
            _3911 <= _3156;
        7:
            _3911 <= _3159;
        8:
            _3911 <= _3162;
        9:
            _3911 <= _3165;
        10:
            _3911 <= _3168;
        11:
            _3911 <= _3171;
        12:
            _3911 <= _3174;
        13:
            _3911 <= _3177;
        14:
            _3911 <= _3180;
        15:
            _3911 <= _3183;
        16:
            _3911 <= _3186;
        17:
            _3911 <= _3189;
        18:
            _3911 <= _3192;
        19:
            _3911 <= _3195;
        20:
            _3911 <= _3198;
        21:
            _3911 <= _3201;
        22:
            _3911 <= _3204;
        23:
            _3911 <= _3207;
        24:
            _3911 <= _3210;
        25:
            _3911 <= _3213;
        26:
            _3911 <= _3216;
        27:
            _3911 <= _3219;
        28:
            _3911 <= _3222;
        29:
            _3911 <= _3225;
        30:
            _3911 <= _3228;
        31:
            _3911 <= _3231;
        32:
            _3911 <= _3234;
        33:
            _3911 <= _3237;
        34:
            _3911 <= _3240;
        35:
            _3911 <= _3243;
        36:
            _3911 <= _3246;
        37:
            _3911 <= _3249;
        38:
            _3911 <= _3252;
        39:
            _3911 <= _3255;
        40:
            _3911 <= _3258;
        41:
            _3911 <= _3261;
        42:
            _3911 <= _3264;
        43:
            _3911 <= _3267;
        44:
            _3911 <= _3270;
        45:
            _3911 <= _3273;
        46:
            _3911 <= _3276;
        47:
            _3911 <= _3279;
        48:
            _3911 <= _3282;
        49:
            _3911 <= _3285;
        50:
            _3911 <= _3288;
        51:
            _3911 <= _3291;
        52:
            _3911 <= _3294;
        53:
            _3911 <= _3297;
        54:
            _3911 <= _3300;
        55:
            _3911 <= _3303;
        56:
            _3911 <= _3306;
        57:
            _3911 <= _3309;
        58:
            _3911 <= _3312;
        59:
            _3911 <= _3315;
        60:
            _3911 <= _3318;
        61:
            _3911 <= _3321;
        62:
            _3911 <= _3324;
        63:
            _3911 <= _3327;
        64:
            _3911 <= _3330;
        65:
            _3911 <= _3333;
        66:
            _3911 <= _3336;
        67:
            _3911 <= _3339;
        68:
            _3911 <= _3342;
        69:
            _3911 <= _3345;
        70:
            _3911 <= _3348;
        71:
            _3911 <= _3351;
        72:
            _3911 <= _3354;
        73:
            _3911 <= _3357;
        74:
            _3911 <= _3360;
        75:
            _3911 <= _3363;
        76:
            _3911 <= _3366;
        77:
            _3911 <= _3369;
        78:
            _3911 <= _3372;
        79:
            _3911 <= _3375;
        80:
            _3911 <= _3378;
        81:
            _3911 <= _3381;
        82:
            _3911 <= _3384;
        83:
            _3911 <= _3387;
        84:
            _3911 <= _3390;
        85:
            _3911 <= _3393;
        86:
            _3911 <= _3396;
        87:
            _3911 <= _3399;
        88:
            _3911 <= _3402;
        89:
            _3911 <= _3405;
        90:
            _3911 <= _3408;
        91:
            _3911 <= _3411;
        92:
            _3911 <= _3414;
        93:
            _3911 <= _3417;
        94:
            _3911 <= _3420;
        95:
            _3911 <= _3423;
        96:
            _3911 <= _3426;
        97:
            _3911 <= _3429;
        98:
            _3911 <= _3432;
        99:
            _3911 <= _3435;
        100:
            _3911 <= _3438;
        101:
            _3911 <= _3441;
        102:
            _3911 <= _3444;
        103:
            _3911 <= _3447;
        104:
            _3911 <= _3450;
        105:
            _3911 <= _3453;
        106:
            _3911 <= _3456;
        107:
            _3911 <= _3459;
        108:
            _3911 <= _3462;
        109:
            _3911 <= _3465;
        110:
            _3911 <= _3468;
        111:
            _3911 <= _3471;
        112:
            _3911 <= _3474;
        113:
            _3911 <= _3477;
        114:
            _3911 <= _3480;
        115:
            _3911 <= _3483;
        116:
            _3911 <= _3486;
        117:
            _3911 <= _3489;
        118:
            _3911 <= _3492;
        119:
            _3911 <= _3495;
        120:
            _3911 <= _3498;
        121:
            _3911 <= _3501;
        122:
            _3911 <= _3504;
        123:
            _3911 <= _3507;
        124:
            _3911 <= _3510;
        125:
            _3911 <= _3513;
        126:
            _3911 <= _3516;
        127:
            _3911 <= _3519;
        128:
            _3911 <= _3522;
        129:
            _3911 <= _3525;
        130:
            _3911 <= _3528;
        131:
            _3911 <= _3531;
        132:
            _3911 <= _3534;
        133:
            _3911 <= _3537;
        134:
            _3911 <= _3540;
        135:
            _3911 <= _3543;
        136:
            _3911 <= _3546;
        137:
            _3911 <= _3549;
        138:
            _3911 <= _3552;
        139:
            _3911 <= _3555;
        140:
            _3911 <= _3558;
        141:
            _3911 <= _3561;
        142:
            _3911 <= _3564;
        143:
            _3911 <= _3567;
        144:
            _3911 <= _3570;
        145:
            _3911 <= _3573;
        146:
            _3911 <= _3576;
        147:
            _3911 <= _3579;
        148:
            _3911 <= _3582;
        149:
            _3911 <= _3585;
        150:
            _3911 <= _3588;
        151:
            _3911 <= _3591;
        152:
            _3911 <= _3594;
        153:
            _3911 <= _3597;
        154:
            _3911 <= _3600;
        155:
            _3911 <= _3603;
        156:
            _3911 <= _3606;
        157:
            _3911 <= _3609;
        158:
            _3911 <= _3612;
        159:
            _3911 <= _3615;
        160:
            _3911 <= _3618;
        161:
            _3911 <= _3621;
        162:
            _3911 <= _3624;
        163:
            _3911 <= _3627;
        164:
            _3911 <= _3630;
        165:
            _3911 <= _3633;
        166:
            _3911 <= _3636;
        167:
            _3911 <= _3639;
        168:
            _3911 <= _3642;
        169:
            _3911 <= _3645;
        170:
            _3911 <= _3648;
        171:
            _3911 <= _3651;
        172:
            _3911 <= _3654;
        173:
            _3911 <= _3657;
        174:
            _3911 <= _3660;
        175:
            _3911 <= _3663;
        176:
            _3911 <= _3666;
        177:
            _3911 <= _3669;
        178:
            _3911 <= _3672;
        179:
            _3911 <= _3675;
        180:
            _3911 <= _3678;
        181:
            _3911 <= _3681;
        182:
            _3911 <= _3684;
        183:
            _3911 <= _3687;
        184:
            _3911 <= _3690;
        185:
            _3911 <= _3693;
        186:
            _3911 <= _3696;
        187:
            _3911 <= _3699;
        188:
            _3911 <= _3702;
        189:
            _3911 <= _3705;
        190:
            _3911 <= _3708;
        191:
            _3911 <= _3711;
        192:
            _3911 <= _3714;
        193:
            _3911 <= _3717;
        194:
            _3911 <= _3720;
        195:
            _3911 <= _3723;
        196:
            _3911 <= _3726;
        197:
            _3911 <= _3729;
        198:
            _3911 <= _3732;
        199:
            _3911 <= _3735;
        200:
            _3911 <= _3738;
        201:
            _3911 <= _3741;
        202:
            _3911 <= _3744;
        203:
            _3911 <= _3747;
        204:
            _3911 <= _3750;
        205:
            _3911 <= _3753;
        206:
            _3911 <= _3756;
        207:
            _3911 <= _3759;
        208:
            _3911 <= _3762;
        209:
            _3911 <= _3765;
        210:
            _3911 <= _3768;
        211:
            _3911 <= _3771;
        212:
            _3911 <= _3774;
        213:
            _3911 <= _3777;
        214:
            _3911 <= _3780;
        215:
            _3911 <= _3783;
        216:
            _3911 <= _3786;
        217:
            _3911 <= _3789;
        218:
            _3911 <= _3792;
        219:
            _3911 <= _3795;
        220:
            _3911 <= _3798;
        221:
            _3911 <= _3801;
        222:
            _3911 <= _3804;
        223:
            _3911 <= _3807;
        224:
            _3911 <= _3810;
        225:
            _3911 <= _3813;
        226:
            _3911 <= _3816;
        227:
            _3911 <= _3819;
        228:
            _3911 <= _3822;
        229:
            _3911 <= _3825;
        230:
            _3911 <= _3828;
        231:
            _3911 <= _3831;
        232:
            _3911 <= _3834;
        233:
            _3911 <= _3837;
        234:
            _3911 <= _3840;
        235:
            _3911 <= _3843;
        236:
            _3911 <= _3846;
        237:
            _3911 <= _3849;
        238:
            _3911 <= _3852;
        239:
            _3911 <= _3855;
        240:
            _3911 <= _3858;
        241:
            _3911 <= _3861;
        242:
            _3911 <= _3864;
        243:
            _3911 <= _3867;
        244:
            _3911 <= _3870;
        245:
            _3911 <= _3873;
        246:
            _3911 <= _3876;
        247:
            _3911 <= _3879;
        248:
            _3911 <= _3882;
        249:
            _3911 <= _3885;
        250:
            _3911 <= _3888;
        251:
            _3911 <= _3891;
        252:
            _3911 <= _3894;
        253:
            _3911 <= _3897;
        254:
            _3911 <= _3900;
        default:
            _3911 <= _3903;
        endcase
    end
    assign _3920 = _3911 == _3919;
    assign _3921 = ~ _3920;
    assign _3922 = _3135 & _3921;
    assign _4698 = _3922 & _4697;
    assign _11989 = _3132 & _4698;
    assign _11993 = _11989 ? _5287 : _11992;
    assign _11988 = _5292 & _11965;
    assign _11994 = _11988 ? _3131 : _11993;
    assign _11986 = _4729 == _787;
    assign _11987 = _4714 & _11986;
    assign _11995 = _11987 ? _5291 : _11994;
    assign _11984 = _3128 & _3135;
    assign _11985 = _11984 & _793;
    assign _11996 = _11985 ? _4713 : _11995;
    assign _11978 = _5296 + _3104;
    assign _11972 = _805 ? _3118 : _5296;
    assign _11968 = _811 == _809;
    assign _11969 = _11968 & _814;
    assign _11970 = _11969 & _801;
    assign _11974 = _11970 ? _3118 : _11972;
    assign _787 = n_nodes;
    assign vdd = 1'b1;
    assign _789 = clear;
    assign _791 = clock;
    assign _11962 = _4729 + _3104;
    assign _11958 = _805 ? _3118 : _4729;
    assign _793 = edge_last;
    assign _795 = edge_valid;
    assign _3131 = 3'b101;
    assign _3132 = _811 == _3131;
    assign _3133 = _3132 & _797;
    assign _797 = edge_phase;
    assign _3129 = ~ _797;
    assign _3130 = _3128 & _3129;
    assign _3134 = _3130 | _3133;
    assign _3135 = _3134 & _795;
    assign _3127 = 3'b010;
    assign _3128 = _811 == _3127;
    assign _4715 = _3128 & _3135;
    assign _4716 = _4715 & _793;
    assign _11960 = _4716 ? _3118 : _11958;
    assign _11963 = _4714 ? _11962 : _11960;
    assign _798 = _11963;
    always @(posedge _791) begin
        if (_789)
            _4729 <= _3118;
        else
            _4729 <= _798;
    end
    assign _5269 = _4729 == _787;
    assign _4713 = 3'b011;
    assign _4714 = _811 == _4713;
    assign _5270 = _4714 & _5269;
    assign _11976 = _5270 ? _3118 : _11974;
    assign _11966 = ~ _11965;
    assign _11967 = _5293 & _11966;
    assign _11979 = _11967 ? _11978 : _11976;
    assign _799 = _11979;
    always @(posedge _791) begin
        if (_789)
            _5296 <= _3118;
        else
            _5296 <= _799;
    end
    assign _11964 = _5296 == _787;
    assign _5291 = 3'b100;
    assign _5292 = _811 == _5291;
    assign _5293 = _5290 | _5292;
    assign _11965 = _5293 & _11964;
    assign _5289 = 3'b001;
    assign _5290 = _811 == _5289;
    assign _11983 = _5290 & _11965;
    assign _11997 = _11983 ? _3127 : _11996;
    assign _801 = x0_last;
    assign _803 = x0_valid;
    assign _814 = _813 & _803;
    assign _11980 = _811 == _809;
    assign _11981 = _11980 & _814;
    assign _11982 = _11981 & _801;
    assign _11998 = _11982 ? _5289 : _11997;
    assign _805 = load;
    assign _11999 = _805 ? _809 : _11998;
    assign _806 = _11999;
    always @(posedge _791) begin
        if (_789)
            _811 <= _809;
        else
            _811 <= _806;
    end
    assign _813 = _811 == _809;
    assign x0_ready = _813;
    assign edge_ready = _3134;
    assign done_ = _5288;
    assign part1_result = _5273;
    assign part2_result = _4701;
    assign state = _811;

endmodule
