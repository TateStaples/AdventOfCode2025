module day3_opt_b (
    length,
    data,
    clear,
    clock,
    k,
    start,
    result,
    done_
);

    input [7:0] length;
    input [511:0] data;
    input clear;
    input clock;
    input [3:0] k;
    input start;
    output [63:0] result;
    output done_;

    wire _39;
    wire _42;
    reg _43;
    wire _1;
    reg _40;
    wire [63:0] _323;
    wire [59:0] _428;
    wire [63:0] _429;
    wire [63:0] _425;
    wire [127:0] _426;
    wire [63:0] _427;
    wire [63:0] _430;
    wire [63:0] _422;
    wire [127:0] _419;
    wire [63:0] _420;
    wire [63:0] _423;
    wire [63:0] _415;
    wire [127:0] _412;
    wire [63:0] _413;
    wire [63:0] _416;
    wire [63:0] _408;
    wire [127:0] _405;
    wire [63:0] _406;
    wire [63:0] _409;
    wire [63:0] _401;
    wire [127:0] _398;
    wire [63:0] _399;
    wire [63:0] _402;
    wire [63:0] _394;
    wire [127:0] _391;
    wire [63:0] _392;
    wire [63:0] _395;
    wire [63:0] _387;
    wire [127:0] _384;
    wire [63:0] _385;
    wire [63:0] _388;
    wire [63:0] _380;
    wire [127:0] _377;
    wire [63:0] _378;
    wire [63:0] _381;
    wire [63:0] _373;
    wire [127:0] _370;
    wire [63:0] _371;
    wire [63:0] _374;
    wire [63:0] _366;
    wire [127:0] _363;
    wire [63:0] _364;
    wire [63:0] _367;
    wire [63:0] _359;
    wire [127:0] _356;
    wire [63:0] _357;
    wire [63:0] _360;
    wire [63:0] _353;
    wire [3:0] _349;
    wire _350;
    wire [63:0] _354;
    wire [3:0] _347;
    wire _348;
    wire [63:0] _361;
    wire [3:0] _345;
    wire _346;
    wire [63:0] _368;
    wire [3:0] _343;
    wire _344;
    wire [63:0] _375;
    wire [3:0] _341;
    wire _342;
    wire [63:0] _382;
    wire [3:0] _339;
    wire _340;
    wire [63:0] _389;
    wire [3:0] _337;
    wire _338;
    wire [63:0] _396;
    wire [3:0] _335;
    wire _336;
    wire [63:0] _403;
    wire [3:0] _333;
    wire _334;
    wire [63:0] _410;
    wire [3:0] _331;
    wire _332;
    wire [63:0] _417;
    wire [3:0] _329;
    wire _330;
    wire [63:0] _424;
    wire [3:0] _327;
    wire _328;
    wire [63:0] _431;
    wire [63:0] _326;
    wire [2:0] _35;
    wire [2:0] _317;
    wire [2:0] _316;
    wire _314;
    wire _315;
    wire [2:0] _318;
    wire [2:0] _312;
    wire [2:0] _313;
    wire [2:0] _308;
    wire [7:0] _294;
    wire [7:0] _45;
    wire [7:0] _48;
    wire [7:0] _49;
    wire [7:0] _4;
    wire [7:0] _47;
    reg [7:0] _50;
    wire [7:0] _5;
    reg [7:0] _46;
    wire [3:0] _290;
    wire [7:0] _291;
    wire [7:0] _292;
    wire _295;
    wire _296;
    wire _59;
    wire _60;
    wire [3:0] _196;
    wire [3:0] _6;
    reg [3:0] _63;
    wire _198;
    wire _199;
    wire [3:0] _203;
    wire [3:0] _7;
    reg [3:0] _202;
    wire _205;
    wire _206;
    wire [3:0] _210;
    wire [3:0] _8;
    reg [3:0] _209;
    wire _212;
    wire _213;
    wire [3:0] _217;
    wire [3:0] _9;
    reg [3:0] _216;
    wire _219;
    wire _220;
    wire [3:0] _224;
    wire [3:0] _10;
    reg [3:0] _223;
    wire _226;
    wire _227;
    wire [3:0] _231;
    wire [3:0] _11;
    reg [3:0] _230;
    wire _233;
    wire _234;
    wire [3:0] _238;
    wire [3:0] _12;
    reg [3:0] _237;
    wire _240;
    wire _241;
    wire [3:0] _245;
    wire [3:0] _13;
    reg [3:0] _244;
    wire _247;
    wire _248;
    wire [3:0] _252;
    wire [3:0] _14;
    reg [3:0] _251;
    wire _254;
    wire _255;
    wire [3:0] _259;
    wire [3:0] _15;
    reg [3:0] _258;
    wire _261;
    wire _262;
    wire [3:0] _266;
    wire [3:0] _16;
    reg [3:0] _265;
    wire [3:0] _194;
    wire [3:0] _193;
    wire [3:0] _192;
    wire [3:0] _191;
    wire [3:0] _190;
    wire [3:0] _189;
    wire [3:0] _188;
    wire [3:0] _187;
    wire [3:0] _186;
    wire [3:0] _185;
    wire [3:0] _184;
    wire [3:0] _183;
    wire [3:0] _182;
    wire [3:0] _181;
    wire [3:0] _180;
    wire [3:0] _179;
    wire [3:0] _178;
    wire [3:0] _177;
    wire [3:0] _176;
    wire [3:0] _175;
    wire [3:0] _174;
    wire [3:0] _173;
    wire [3:0] _172;
    wire [3:0] _171;
    wire [3:0] _170;
    wire [3:0] _169;
    wire [3:0] _168;
    wire [3:0] _167;
    wire [3:0] _166;
    wire [3:0] _165;
    wire [3:0] _164;
    wire [3:0] _163;
    wire [3:0] _162;
    wire [3:0] _161;
    wire [3:0] _160;
    wire [3:0] _159;
    wire [3:0] _158;
    wire [3:0] _157;
    wire [3:0] _156;
    wire [3:0] _155;
    wire [3:0] _154;
    wire [3:0] _153;
    wire [3:0] _152;
    wire [3:0] _151;
    wire [3:0] _150;
    wire [3:0] _149;
    wire [3:0] _148;
    wire [3:0] _147;
    wire [3:0] _146;
    wire [3:0] _145;
    wire [3:0] _144;
    wire [3:0] _143;
    wire [3:0] _142;
    wire [3:0] _141;
    wire [3:0] _140;
    wire [3:0] _139;
    wire [3:0] _138;
    wire [3:0] _137;
    wire [3:0] _136;
    wire [3:0] _135;
    wire [3:0] _134;
    wire [3:0] _133;
    wire [3:0] _132;
    wire [3:0] _131;
    wire [3:0] _130;
    wire [3:0] _129;
    wire [3:0] _128;
    wire [3:0] _127;
    wire [3:0] _126;
    wire [3:0] _125;
    wire [3:0] _124;
    wire [3:0] _123;
    wire [3:0] _122;
    wire [3:0] _121;
    wire [3:0] _120;
    wire [3:0] _119;
    wire [3:0] _118;
    wire [3:0] _117;
    wire [3:0] _116;
    wire [3:0] _115;
    wire [3:0] _114;
    wire [3:0] _113;
    wire [3:0] _112;
    wire [3:0] _111;
    wire [3:0] _110;
    wire [3:0] _109;
    wire [3:0] _108;
    wire [3:0] _107;
    wire [3:0] _106;
    wire [3:0] _105;
    wire [3:0] _104;
    wire [3:0] _103;
    wire [3:0] _102;
    wire [3:0] _101;
    wire [3:0] _100;
    wire [3:0] _99;
    wire [3:0] _98;
    wire [3:0] _97;
    wire [3:0] _96;
    wire [3:0] _95;
    wire [3:0] _94;
    wire [3:0] _93;
    wire [3:0] _92;
    wire [3:0] _91;
    wire [3:0] _90;
    wire [3:0] _89;
    wire [3:0] _88;
    wire [3:0] _87;
    wire [3:0] _86;
    wire [3:0] _85;
    wire [3:0] _84;
    wire [3:0] _83;
    wire [3:0] _82;
    wire [3:0] _81;
    wire [3:0] _80;
    wire [3:0] _79;
    wire [3:0] _78;
    wire [3:0] _77;
    wire [3:0] _76;
    wire [3:0] _75;
    wire [3:0] _74;
    wire [3:0] _73;
    wire [3:0] _72;
    wire [3:0] _71;
    wire [3:0] _70;
    wire [3:0] _69;
    wire [3:0] _68;
    wire [511:0] _18;
    wire [3:0] _67;
    wire [7:0] _270;
    wire [7:0] _268;
    reg [7:0] _271;
    wire [7:0] _19;
    reg [7:0] _66;
    reg [3:0] _195;
    wire _273;
    wire _274;
    wire [3:0] _278;
    wire [3:0] _20;
    reg [3:0] _277;
    wire [3:0] _284;
    reg [3:0] _285;
    wire _286;
    wire [3:0] _302;
    wire vdd;
    wire _22;
    wire _24;
    wire [3:0] _26;
    wire [3:0] _279;
    wire [3:0] _27;
    reg [3:0] _56;
    wire _57;
    wire [3:0] _303;
    wire [3:0] _299;
    wire [3:0] _300;
    wire [3:0] _281;
    reg [3:0] _304;
    wire [3:0] _28;
    reg [3:0] _53;
    wire _282;
    wire _287;
    wire _297;
    wire [2:0] _310;
    wire _30;
    wire [2:0] _307;
    reg [2:0] _321;
    wire [2:0] _31;
    reg [2:0] _37;
    reg [63:0] _432;
    wire [63:0] _32;
    reg [63:0] _324;
    assign _39 = 1'b0;
    assign _42 = _30 ? _39 : _40;
    always @* begin
        case (_37)
        0:
            _43 <= _42;
        1:
            _43 <= _40;
        2:
            _43 <= _40;
        3:
            _43 <= _40;
        4:
            _43 <= vdd;
        5:
            _43 <= _40;
        6:
            _43 <= _40;
        default:
            _43 <= _40;
        endcase
    end
    assign _1 = _43;
    always @(posedge _24) begin
        if (_22)
            _40 <= _39;
        else
            _40 <= _1;
    end
    assign _323 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign _428 = 60'b000000000000000000000000000000000000000000000000000000000000;
    assign _429 = { _428,
                    _63 };
    assign _425 = 64'b0000000000000000000000000000000000000000000000000000000000001010;
    assign _426 = _424 * _425;
    assign _427 = _426[63:0];
    assign _430 = _427 + _429;
    assign _422 = { _428,
                    _202 };
    assign _419 = _417 * _425;
    assign _420 = _419[63:0];
    assign _423 = _420 + _422;
    assign _415 = { _428,
                    _209 };
    assign _412 = _410 * _425;
    assign _413 = _412[63:0];
    assign _416 = _413 + _415;
    assign _408 = { _428,
                    _216 };
    assign _405 = _403 * _425;
    assign _406 = _405[63:0];
    assign _409 = _406 + _408;
    assign _401 = { _428,
                    _223 };
    assign _398 = _396 * _425;
    assign _399 = _398[63:0];
    assign _402 = _399 + _401;
    assign _394 = { _428,
                    _230 };
    assign _391 = _389 * _425;
    assign _392 = _391[63:0];
    assign _395 = _392 + _394;
    assign _387 = { _428,
                    _237 };
    assign _384 = _382 * _425;
    assign _385 = _384[63:0];
    assign _388 = _385 + _387;
    assign _380 = { _428,
                    _244 };
    assign _377 = _375 * _425;
    assign _378 = _377[63:0];
    assign _381 = _378 + _380;
    assign _373 = { _428,
                    _251 };
    assign _370 = _368 * _425;
    assign _371 = _370[63:0];
    assign _374 = _371 + _373;
    assign _366 = { _428,
                    _258 };
    assign _363 = _361 * _425;
    assign _364 = _363[63:0];
    assign _367 = _364 + _366;
    assign _359 = { _428,
                    _265 };
    assign _356 = _354 * _425;
    assign _357 = _356[63:0];
    assign _360 = _357 + _359;
    assign _353 = { _428,
                    _277 };
    assign _349 = 4'b0000;
    assign _350 = _349 < _56;
    assign _354 = _350 ? _353 : _323;
    assign _347 = 4'b0001;
    assign _348 = _347 < _56;
    assign _361 = _348 ? _360 : _354;
    assign _345 = 4'b0010;
    assign _346 = _345 < _56;
    assign _368 = _346 ? _367 : _361;
    assign _343 = 4'b0011;
    assign _344 = _343 < _56;
    assign _375 = _344 ? _374 : _368;
    assign _341 = 4'b0100;
    assign _342 = _341 < _56;
    assign _382 = _342 ? _381 : _375;
    assign _339 = 4'b0101;
    assign _340 = _339 < _56;
    assign _389 = _340 ? _388 : _382;
    assign _337 = 4'b0110;
    assign _338 = _337 < _56;
    assign _396 = _338 ? _395 : _389;
    assign _335 = 4'b0111;
    assign _336 = _335 < _56;
    assign _403 = _336 ? _402 : _396;
    assign _333 = 4'b1000;
    assign _334 = _333 < _56;
    assign _410 = _334 ? _409 : _403;
    assign _331 = 4'b1001;
    assign _332 = _331 < _56;
    assign _417 = _332 ? _416 : _410;
    assign _329 = 4'b1010;
    assign _330 = _329 < _56;
    assign _424 = _330 ? _423 : _417;
    assign _327 = 4'b1011;
    assign _328 = _327 < _56;
    assign _431 = _328 ? _430 : _424;
    assign _326 = _30 ? _323 : _324;
    assign _35 = 3'b000;
    assign _317 = 3'b100;
    assign _316 = 3'b001;
    assign _314 = _66 < _4;
    assign _315 = ~ _314;
    assign _318 = _315 ? _317 : _316;
    assign _312 = 3'b011;
    assign _313 = _57 ? _312 : _312;
    assign _308 = 3'b010;
    assign _294 = { _349,
                    _56 };
    assign _45 = 8'b00000000;
    assign _48 = 8'b00000001;
    assign _49 = _46 - _48;
    assign _4 = length;
    assign _47 = _30 ? _4 : _46;
    always @* begin
        case (_37)
        0:
            _50 <= _47;
        1:
            _50 <= _46;
        2:
            _50 <= _46;
        3:
            _50 <= _49;
        4:
            _50 <= _46;
        5:
            _50 <= _46;
        6:
            _50 <= _46;
        default:
            _50 <= _46;
        endcase
    end
    assign _5 = _50;
    always @(posedge _24) begin
        if (_22)
            _46 <= _45;
        else
            _46 <= _5;
    end
    assign _290 = _53 - _347;
    assign _291 = { _349,
                    _290 };
    assign _292 = _291 + _46;
    assign _295 = _292 < _294;
    assign _296 = ~ _295;
    assign _59 = _327 == _53;
    assign _60 = _57 & _59;
    assign _196 = _60 ? _195 : _63;
    assign _6 = _196;
    always @(posedge _24) begin
        if (_22)
            _63 <= _349;
        else
            _63 <= _6;
    end
    assign _198 = _329 == _53;
    assign _199 = _57 & _198;
    assign _203 = _199 ? _195 : _202;
    assign _7 = _203;
    always @(posedge _24) begin
        if (_22)
            _202 <= _349;
        else
            _202 <= _7;
    end
    assign _205 = _331 == _53;
    assign _206 = _57 & _205;
    assign _210 = _206 ? _195 : _209;
    assign _8 = _210;
    always @(posedge _24) begin
        if (_22)
            _209 <= _349;
        else
            _209 <= _8;
    end
    assign _212 = _333 == _53;
    assign _213 = _57 & _212;
    assign _217 = _213 ? _195 : _216;
    assign _9 = _217;
    always @(posedge _24) begin
        if (_22)
            _216 <= _349;
        else
            _216 <= _9;
    end
    assign _219 = _335 == _53;
    assign _220 = _57 & _219;
    assign _224 = _220 ? _195 : _223;
    assign _10 = _224;
    always @(posedge _24) begin
        if (_22)
            _223 <= _349;
        else
            _223 <= _10;
    end
    assign _226 = _337 == _53;
    assign _227 = _57 & _226;
    assign _231 = _227 ? _195 : _230;
    assign _11 = _231;
    always @(posedge _24) begin
        if (_22)
            _230 <= _349;
        else
            _230 <= _11;
    end
    assign _233 = _339 == _53;
    assign _234 = _57 & _233;
    assign _238 = _234 ? _195 : _237;
    assign _12 = _238;
    always @(posedge _24) begin
        if (_22)
            _237 <= _349;
        else
            _237 <= _12;
    end
    assign _240 = _341 == _53;
    assign _241 = _57 & _240;
    assign _245 = _241 ? _195 : _244;
    assign _13 = _245;
    always @(posedge _24) begin
        if (_22)
            _244 <= _349;
        else
            _244 <= _13;
    end
    assign _247 = _343 == _53;
    assign _248 = _57 & _247;
    assign _252 = _248 ? _195 : _251;
    assign _14 = _252;
    always @(posedge _24) begin
        if (_22)
            _251 <= _349;
        else
            _251 <= _14;
    end
    assign _254 = _345 == _53;
    assign _255 = _57 & _254;
    assign _259 = _255 ? _195 : _258;
    assign _15 = _259;
    always @(posedge _24) begin
        if (_22)
            _258 <= _349;
        else
            _258 <= _15;
    end
    assign _261 = _347 == _53;
    assign _262 = _57 & _261;
    assign _266 = _262 ? _195 : _265;
    assign _16 = _266;
    always @(posedge _24) begin
        if (_22)
            _265 <= _349;
        else
            _265 <= _16;
    end
    assign _194 = _18[511:508];
    assign _193 = _18[507:504];
    assign _192 = _18[503:500];
    assign _191 = _18[499:496];
    assign _190 = _18[495:492];
    assign _189 = _18[491:488];
    assign _188 = _18[487:484];
    assign _187 = _18[483:480];
    assign _186 = _18[479:476];
    assign _185 = _18[475:472];
    assign _184 = _18[471:468];
    assign _183 = _18[467:464];
    assign _182 = _18[463:460];
    assign _181 = _18[459:456];
    assign _180 = _18[455:452];
    assign _179 = _18[451:448];
    assign _178 = _18[447:444];
    assign _177 = _18[443:440];
    assign _176 = _18[439:436];
    assign _175 = _18[435:432];
    assign _174 = _18[431:428];
    assign _173 = _18[427:424];
    assign _172 = _18[423:420];
    assign _171 = _18[419:416];
    assign _170 = _18[415:412];
    assign _169 = _18[411:408];
    assign _168 = _18[407:404];
    assign _167 = _18[403:400];
    assign _166 = _18[399:396];
    assign _165 = _18[395:392];
    assign _164 = _18[391:388];
    assign _163 = _18[387:384];
    assign _162 = _18[383:380];
    assign _161 = _18[379:376];
    assign _160 = _18[375:372];
    assign _159 = _18[371:368];
    assign _158 = _18[367:364];
    assign _157 = _18[363:360];
    assign _156 = _18[359:356];
    assign _155 = _18[355:352];
    assign _154 = _18[351:348];
    assign _153 = _18[347:344];
    assign _152 = _18[343:340];
    assign _151 = _18[339:336];
    assign _150 = _18[335:332];
    assign _149 = _18[331:328];
    assign _148 = _18[327:324];
    assign _147 = _18[323:320];
    assign _146 = _18[319:316];
    assign _145 = _18[315:312];
    assign _144 = _18[311:308];
    assign _143 = _18[307:304];
    assign _142 = _18[303:300];
    assign _141 = _18[299:296];
    assign _140 = _18[295:292];
    assign _139 = _18[291:288];
    assign _138 = _18[287:284];
    assign _137 = _18[283:280];
    assign _136 = _18[279:276];
    assign _135 = _18[275:272];
    assign _134 = _18[271:268];
    assign _133 = _18[267:264];
    assign _132 = _18[263:260];
    assign _131 = _18[259:256];
    assign _130 = _18[255:252];
    assign _129 = _18[251:248];
    assign _128 = _18[247:244];
    assign _127 = _18[243:240];
    assign _126 = _18[239:236];
    assign _125 = _18[235:232];
    assign _124 = _18[231:228];
    assign _123 = _18[227:224];
    assign _122 = _18[223:220];
    assign _121 = _18[219:216];
    assign _120 = _18[215:212];
    assign _119 = _18[211:208];
    assign _118 = _18[207:204];
    assign _117 = _18[203:200];
    assign _116 = _18[199:196];
    assign _115 = _18[195:192];
    assign _114 = _18[191:188];
    assign _113 = _18[187:184];
    assign _112 = _18[183:180];
    assign _111 = _18[179:176];
    assign _110 = _18[175:172];
    assign _109 = _18[171:168];
    assign _108 = _18[167:164];
    assign _107 = _18[163:160];
    assign _106 = _18[159:156];
    assign _105 = _18[155:152];
    assign _104 = _18[151:148];
    assign _103 = _18[147:144];
    assign _102 = _18[143:140];
    assign _101 = _18[139:136];
    assign _100 = _18[135:132];
    assign _99 = _18[131:128];
    assign _98 = _18[127:124];
    assign _97 = _18[123:120];
    assign _96 = _18[119:116];
    assign _95 = _18[115:112];
    assign _94 = _18[111:108];
    assign _93 = _18[107:104];
    assign _92 = _18[103:100];
    assign _91 = _18[99:96];
    assign _90 = _18[95:92];
    assign _89 = _18[91:88];
    assign _88 = _18[87:84];
    assign _87 = _18[83:80];
    assign _86 = _18[79:76];
    assign _85 = _18[75:72];
    assign _84 = _18[71:68];
    assign _83 = _18[67:64];
    assign _82 = _18[63:60];
    assign _81 = _18[59:56];
    assign _80 = _18[55:52];
    assign _79 = _18[51:48];
    assign _78 = _18[47:44];
    assign _77 = _18[43:40];
    assign _76 = _18[39:36];
    assign _75 = _18[35:32];
    assign _74 = _18[31:28];
    assign _73 = _18[27:24];
    assign _72 = _18[23:20];
    assign _71 = _18[19:16];
    assign _70 = _18[15:12];
    assign _69 = _18[11:8];
    assign _68 = _18[7:4];
    assign _18 = data;
    assign _67 = _18[3:0];
    assign _270 = _66 + _48;
    assign _268 = _30 ? _45 : _66;
    always @* begin
        case (_37)
        0:
            _271 <= _268;
        1:
            _271 <= _66;
        2:
            _271 <= _66;
        3:
            _271 <= _270;
        4:
            _271 <= _66;
        5:
            _271 <= _66;
        6:
            _271 <= _66;
        default:
            _271 <= _66;
        endcase
    end
    assign _19 = _271;
    always @(posedge _24) begin
        if (_22)
            _66 <= _45;
        else
            _66 <= _19;
    end
    always @* begin
        case (_66)
        0:
            _195 <= _67;
        1:
            _195 <= _68;
        2:
            _195 <= _69;
        3:
            _195 <= _70;
        4:
            _195 <= _71;
        5:
            _195 <= _72;
        6:
            _195 <= _73;
        7:
            _195 <= _74;
        8:
            _195 <= _75;
        9:
            _195 <= _76;
        10:
            _195 <= _77;
        11:
            _195 <= _78;
        12:
            _195 <= _79;
        13:
            _195 <= _80;
        14:
            _195 <= _81;
        15:
            _195 <= _82;
        16:
            _195 <= _83;
        17:
            _195 <= _84;
        18:
            _195 <= _85;
        19:
            _195 <= _86;
        20:
            _195 <= _87;
        21:
            _195 <= _88;
        22:
            _195 <= _89;
        23:
            _195 <= _90;
        24:
            _195 <= _91;
        25:
            _195 <= _92;
        26:
            _195 <= _93;
        27:
            _195 <= _94;
        28:
            _195 <= _95;
        29:
            _195 <= _96;
        30:
            _195 <= _97;
        31:
            _195 <= _98;
        32:
            _195 <= _99;
        33:
            _195 <= _100;
        34:
            _195 <= _101;
        35:
            _195 <= _102;
        36:
            _195 <= _103;
        37:
            _195 <= _104;
        38:
            _195 <= _105;
        39:
            _195 <= _106;
        40:
            _195 <= _107;
        41:
            _195 <= _108;
        42:
            _195 <= _109;
        43:
            _195 <= _110;
        44:
            _195 <= _111;
        45:
            _195 <= _112;
        46:
            _195 <= _113;
        47:
            _195 <= _114;
        48:
            _195 <= _115;
        49:
            _195 <= _116;
        50:
            _195 <= _117;
        51:
            _195 <= _118;
        52:
            _195 <= _119;
        53:
            _195 <= _120;
        54:
            _195 <= _121;
        55:
            _195 <= _122;
        56:
            _195 <= _123;
        57:
            _195 <= _124;
        58:
            _195 <= _125;
        59:
            _195 <= _126;
        60:
            _195 <= _127;
        61:
            _195 <= _128;
        62:
            _195 <= _129;
        63:
            _195 <= _130;
        64:
            _195 <= _131;
        65:
            _195 <= _132;
        66:
            _195 <= _133;
        67:
            _195 <= _134;
        68:
            _195 <= _135;
        69:
            _195 <= _136;
        70:
            _195 <= _137;
        71:
            _195 <= _138;
        72:
            _195 <= _139;
        73:
            _195 <= _140;
        74:
            _195 <= _141;
        75:
            _195 <= _142;
        76:
            _195 <= _143;
        77:
            _195 <= _144;
        78:
            _195 <= _145;
        79:
            _195 <= _146;
        80:
            _195 <= _147;
        81:
            _195 <= _148;
        82:
            _195 <= _149;
        83:
            _195 <= _150;
        84:
            _195 <= _151;
        85:
            _195 <= _152;
        86:
            _195 <= _153;
        87:
            _195 <= _154;
        88:
            _195 <= _155;
        89:
            _195 <= _156;
        90:
            _195 <= _157;
        91:
            _195 <= _158;
        92:
            _195 <= _159;
        93:
            _195 <= _160;
        94:
            _195 <= _161;
        95:
            _195 <= _162;
        96:
            _195 <= _163;
        97:
            _195 <= _164;
        98:
            _195 <= _165;
        99:
            _195 <= _166;
        100:
            _195 <= _167;
        101:
            _195 <= _168;
        102:
            _195 <= _169;
        103:
            _195 <= _170;
        104:
            _195 <= _171;
        105:
            _195 <= _172;
        106:
            _195 <= _173;
        107:
            _195 <= _174;
        108:
            _195 <= _175;
        109:
            _195 <= _176;
        110:
            _195 <= _177;
        111:
            _195 <= _178;
        112:
            _195 <= _179;
        113:
            _195 <= _180;
        114:
            _195 <= _181;
        115:
            _195 <= _182;
        116:
            _195 <= _183;
        117:
            _195 <= _184;
        118:
            _195 <= _185;
        119:
            _195 <= _186;
        120:
            _195 <= _187;
        121:
            _195 <= _188;
        122:
            _195 <= _189;
        123:
            _195 <= _190;
        124:
            _195 <= _191;
        125:
            _195 <= _192;
        126:
            _195 <= _193;
        default:
            _195 <= _194;
        endcase
    end
    assign _273 = _349 == _53;
    assign _274 = _57 & _273;
    assign _278 = _274 ? _195 : _277;
    assign _20 = _278;
    always @(posedge _24) begin
        if (_22)
            _277 <= _349;
        else
            _277 <= _20;
    end
    assign _284 = _53 - _347;
    always @* begin
        case (_284)
        0:
            _285 <= _277;
        1:
            _285 <= _265;
        2:
            _285 <= _258;
        3:
            _285 <= _251;
        4:
            _285 <= _244;
        5:
            _285 <= _237;
        6:
            _285 <= _230;
        7:
            _285 <= _223;
        8:
            _285 <= _216;
        9:
            _285 <= _209;
        10:
            _285 <= _202;
        default:
            _285 <= _63;
        endcase
    end
    assign _286 = _285 < _195;
    assign _302 = _53 + _347;
    assign vdd = 1'b1;
    assign _22 = clear;
    assign _24 = clock;
    assign _26 = k;
    assign _279 = _30 ? _26 : _56;
    assign _27 = _279;
    always @(posedge _24) begin
        if (_22)
            _56 <= _349;
        else
            _56 <= _27;
    end
    assign _57 = _53 < _56;
    assign _303 = _57 ? _302 : _53;
    assign _299 = _53 - _347;
    assign _300 = _297 ? _299 : _53;
    assign _281 = _30 ? _349 : _53;
    always @* begin
        case (_37)
        0:
            _304 <= _281;
        1:
            _304 <= _300;
        2:
            _304 <= _303;
        3:
            _304 <= _53;
        4:
            _304 <= _53;
        5:
            _304 <= _53;
        6:
            _304 <= _53;
        default:
            _304 <= _53;
        endcase
    end
    assign _28 = _304;
    always @(posedge _24) begin
        if (_22)
            _53 <= _349;
        else
            _53 <= _28;
    end
    assign _282 = _349 < _53;
    assign _287 = _282 & _286;
    assign _297 = _287 & _296;
    assign _310 = _297 ? _316 : _308;
    assign _30 = start;
    assign _307 = _30 ? _312 : _35;
    always @* begin
        case (_37)
        0:
            _321 <= _307;
        1:
            _321 <= _310;
        2:
            _321 <= _313;
        3:
            _321 <= _318;
        4:
            _321 <= _35;
        5:
            _321 <= _35;
        6:
            _321 <= _35;
        default:
            _321 <= _35;
        endcase
    end
    assign _31 = _321;
    always @(posedge _24) begin
        if (_22)
            _37 <= _35;
        else
            _37 <= _31;
    end
    always @* begin
        case (_37)
        0:
            _432 <= _326;
        1:
            _432 <= _324;
        2:
            _432 <= _324;
        3:
            _432 <= _324;
        4:
            _432 <= _431;
        5:
            _432 <= _324;
        6:
            _432 <= _324;
        default:
            _432 <= _324;
        endcase
    end
    assign _32 = _432;
    always @(posedge _24) begin
        if (_22)
            _324 <= _323;
        else
            _324 <= _32;
    end
    assign result = _324;
    assign done_ = _40;

endmodule
