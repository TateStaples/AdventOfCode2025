module day7_opt_b (
    width,
    row_bits,
    clear,
    clock,
    row_last,
    row_valid,
    load,
    ready,
    done_,
    part1_result,
    part2_result,
    state
);

    input [7:0] width;
    input [255:0] row_bits;
    input clear;
    input clock;
    input row_last;
    input row_valid;
    input load;
    output ready;
    output done_;
    output [63:0] part1_result;
    output [63:0] part2_result;
    output [1:0] state;

    wire [63:0] _290;
    wire [63:0] _342;
    wire [63:0] _362;
    wire [63:0] _382;
    wire [63:0] _402;
    wire [63:0] _422;
    wire [63:0] _442;
    wire [63:0] _462;
    wire [63:0] _482;
    wire [63:0] _502;
    wire [63:0] _522;
    wire [63:0] _542;
    wire [63:0] _562;
    wire [63:0] _582;
    wire [63:0] _602;
    wire [63:0] _622;
    wire [63:0] _642;
    wire [63:0] _662;
    wire [63:0] _682;
    wire [63:0] _702;
    wire [63:0] _722;
    wire [63:0] _742;
    wire [63:0] _762;
    wire [63:0] _782;
    wire [63:0] _802;
    wire [63:0] _822;
    wire [63:0] _842;
    wire [63:0] _862;
    wire [63:0] _882;
    wire [63:0] _902;
    wire [63:0] _922;
    wire [63:0] _942;
    wire [63:0] _962;
    wire [63:0] _982;
    wire [63:0] _1002;
    wire [63:0] _1022;
    wire [63:0] _1042;
    wire [63:0] _1062;
    wire [63:0] _1082;
    wire [63:0] _1102;
    wire [63:0] _1122;
    wire [63:0] _1142;
    wire [63:0] _1162;
    wire [63:0] _1182;
    wire [63:0] _1202;
    wire [63:0] _1222;
    wire [63:0] _1242;
    wire [63:0] _1262;
    wire [63:0] _1282;
    wire [63:0] _1302;
    wire [63:0] _1322;
    wire [63:0] _1342;
    wire [63:0] _1362;
    wire [63:0] _1382;
    wire [63:0] _1402;
    wire [63:0] _1422;
    wire [63:0] _1442;
    wire [63:0] _1462;
    wire [63:0] _1482;
    wire [63:0] _1502;
    wire [63:0] _1522;
    wire [63:0] _1542;
    wire [63:0] _1562;
    wire [63:0] _1582;
    wire [63:0] _1602;
    wire [63:0] _1622;
    wire [63:0] _1642;
    wire [63:0] _1662;
    wire [63:0] _1682;
    wire [63:0] _1702;
    wire [63:0] _1722;
    wire [63:0] _1742;
    wire [63:0] _1762;
    wire [63:0] _1782;
    wire [63:0] _1802;
    wire [63:0] _1822;
    wire [63:0] _1842;
    wire [63:0] _1862;
    wire [63:0] _1882;
    wire [63:0] _1902;
    wire [63:0] _1922;
    wire [63:0] _1942;
    wire [63:0] _1962;
    wire [63:0] _1982;
    wire [63:0] _2002;
    wire [63:0] _2022;
    wire [63:0] _2042;
    wire [63:0] _2062;
    wire [63:0] _2082;
    wire [63:0] _2102;
    wire [63:0] _2122;
    wire [63:0] _2142;
    wire [63:0] _2162;
    wire [63:0] _2182;
    wire [63:0] _2202;
    wire [63:0] _2222;
    wire [63:0] _2242;
    wire [63:0] _2262;
    wire [63:0] _2282;
    wire [63:0] _2302;
    wire [63:0] _2322;
    wire [63:0] _2342;
    wire [63:0] _2362;
    wire [63:0] _2382;
    wire [63:0] _2402;
    wire [63:0] _2422;
    wire [63:0] _2442;
    wire [63:0] _2462;
    wire [63:0] _2482;
    wire [63:0] _2502;
    wire [63:0] _2522;
    wire [63:0] _2542;
    wire [63:0] _2562;
    wire [63:0] _2582;
    wire [63:0] _2602;
    wire [63:0] _2622;
    wire [63:0] _2642;
    wire [63:0] _2662;
    wire [63:0] _2682;
    wire [63:0] _2702;
    wire [63:0] _2722;
    wire [63:0] _2742;
    wire [63:0] _2762;
    wire [63:0] _2782;
    wire [63:0] _2802;
    wire [63:0] _2822;
    wire [63:0] _2842;
    wire [63:0] _2862;
    wire [63:0] _2882;
    wire [63:0] _2902;
    wire [63:0] _2922;
    wire [63:0] _2942;
    wire [63:0] _2962;
    wire [63:0] _2982;
    wire [63:0] _3002;
    wire [63:0] _3022;
    wire [63:0] _3042;
    wire [63:0] _3062;
    wire [63:0] _3082;
    wire [63:0] _3102;
    wire [63:0] _3122;
    wire [63:0] _3142;
    wire [63:0] _3162;
    wire [63:0] _3182;
    wire [63:0] _3202;
    wire [63:0] _3222;
    wire [63:0] _3242;
    wire [63:0] _3262;
    wire [63:0] _3282;
    wire [63:0] _3302;
    wire [63:0] _3322;
    wire [63:0] _3342;
    wire [63:0] _3362;
    wire [63:0] _3382;
    wire [63:0] _3402;
    wire [63:0] _3422;
    wire [63:0] _3442;
    wire [63:0] _3462;
    wire [63:0] _3482;
    wire [63:0] _3502;
    wire [63:0] _3522;
    wire [63:0] _3542;
    wire [63:0] _3562;
    wire [63:0] _3582;
    wire [63:0] _3602;
    wire [63:0] _3622;
    wire [63:0] _3642;
    wire [63:0] _3662;
    wire [63:0] _3682;
    wire [63:0] _3702;
    wire [63:0] _3722;
    wire [63:0] _3742;
    wire [63:0] _3762;
    wire [63:0] _3782;
    wire [63:0] _3802;
    wire [63:0] _3822;
    wire [63:0] _3842;
    wire [63:0] _3862;
    wire [63:0] _3882;
    wire [63:0] _3902;
    wire [63:0] _3922;
    wire [63:0] _3942;
    wire [63:0] _3962;
    wire [63:0] _3982;
    wire [63:0] _4002;
    wire [63:0] _4022;
    wire [63:0] _4042;
    wire [63:0] _4062;
    wire [63:0] _4082;
    wire [63:0] _4102;
    wire [63:0] _4122;
    wire [63:0] _4142;
    wire [63:0] _4162;
    wire [63:0] _4182;
    wire [63:0] _4202;
    wire [63:0] _4222;
    wire [63:0] _4242;
    wire [63:0] _4262;
    wire [63:0] _4282;
    wire [63:0] _4302;
    wire [63:0] _4322;
    wire [63:0] _4342;
    wire [63:0] _4362;
    wire [63:0] _4382;
    wire [63:0] _4402;
    wire [63:0] _4422;
    wire [63:0] _4442;
    wire [63:0] _4462;
    wire [63:0] _4482;
    wire [63:0] _4502;
    wire [63:0] _4522;
    wire [63:0] _4542;
    wire [63:0] _4562;
    wire [63:0] _4582;
    wire [63:0] _4602;
    wire [63:0] _4622;
    wire [63:0] _4642;
    wire [63:0] _4662;
    wire [63:0] _4682;
    wire [63:0] _4702;
    wire [63:0] _4722;
    wire [63:0] _4742;
    wire [63:0] _4762;
    wire [63:0] _4782;
    wire [63:0] _4802;
    wire [63:0] _4822;
    wire [63:0] _4842;
    wire [63:0] _4862;
    wire [63:0] _4882;
    wire [63:0] _4902;
    wire [63:0] _4922;
    wire [63:0] _4942;
    wire [63:0] _4962;
    wire [63:0] _4982;
    wire [63:0] _5002;
    wire [63:0] _5022;
    wire [63:0] _5042;
    wire [63:0] _5062;
    wire [63:0] _5082;
    wire [63:0] _5102;
    wire [63:0] _5122;
    wire [63:0] _5142;
    wire [63:0] _5162;
    wire [63:0] _5182;
    wire [63:0] _5202;
    wire [63:0] _5222;
    wire [63:0] _5242;
    wire [63:0] _5262;
    wire [63:0] _5282;
    wire [63:0] _5302;
    wire [63:0] _5322;
    wire [63:0] _5342;
    wire [63:0] _5362;
    wire [63:0] _5382;
    wire [63:0] _5402;
    wire [63:0] _5408;
    wire _288;
    wire [63:0] _5409;
    wire [63:0] _5411;
    wire [63:0] _2;
    reg [63:0] _291;
    wire _8233;
    wire [7:0] _8232;
    wire [8:0] _8234;
    wire _8230;
    wire [8:0] _8231;
    wire [8:0] _8235;
    wire _8226;
    wire [8:0] _8227;
    wire _8223;
    wire [8:0] _8224;
    wire [8:0] _8228;
    wire [8:0] _8236;
    wire _8218;
    wire [8:0] _8219;
    wire _8215;
    wire [8:0] _8216;
    wire [8:0] _8220;
    wire _8211;
    wire [8:0] _8212;
    wire _8208;
    wire [8:0] _8209;
    wire [8:0] _8213;
    wire [8:0] _8221;
    wire [8:0] _8237;
    wire _8202;
    wire [8:0] _8203;
    wire _8199;
    wire [8:0] _8200;
    wire [8:0] _8204;
    wire _8195;
    wire [8:0] _8196;
    wire _8192;
    wire [8:0] _8193;
    wire [8:0] _8197;
    wire [8:0] _8205;
    wire _8187;
    wire [8:0] _8188;
    wire _8184;
    wire [8:0] _8185;
    wire [8:0] _8189;
    wire _8180;
    wire [8:0] _8181;
    wire _8177;
    wire [8:0] _8178;
    wire [8:0] _8182;
    wire [8:0] _8190;
    wire [8:0] _8206;
    wire [8:0] _8238;
    wire _8170;
    wire [8:0] _8171;
    wire _8167;
    wire [8:0] _8168;
    wire [8:0] _8172;
    wire _8163;
    wire [8:0] _8164;
    wire _8160;
    wire [8:0] _8161;
    wire [8:0] _8165;
    wire [8:0] _8173;
    wire _8155;
    wire [8:0] _8156;
    wire _8152;
    wire [8:0] _8153;
    wire [8:0] _8157;
    wire _8148;
    wire [8:0] _8149;
    wire _8145;
    wire [8:0] _8146;
    wire [8:0] _8150;
    wire [8:0] _8158;
    wire [8:0] _8174;
    wire _8139;
    wire [8:0] _8140;
    wire _8136;
    wire [8:0] _8137;
    wire [8:0] _8141;
    wire _8132;
    wire [8:0] _8133;
    wire _8129;
    wire [8:0] _8130;
    wire [8:0] _8134;
    wire [8:0] _8142;
    wire _8124;
    wire [8:0] _8125;
    wire _8121;
    wire [8:0] _8122;
    wire [8:0] _8126;
    wire _8117;
    wire [8:0] _8118;
    wire _8114;
    wire [8:0] _8115;
    wire [8:0] _8119;
    wire [8:0] _8127;
    wire [8:0] _8143;
    wire [8:0] _8175;
    wire [8:0] _8239;
    wire _8106;
    wire [8:0] _8107;
    wire _8103;
    wire [8:0] _8104;
    wire [8:0] _8108;
    wire _8099;
    wire [8:0] _8100;
    wire _8096;
    wire [8:0] _8097;
    wire [8:0] _8101;
    wire [8:0] _8109;
    wire _8091;
    wire [8:0] _8092;
    wire _8088;
    wire [8:0] _8089;
    wire [8:0] _8093;
    wire _8084;
    wire [8:0] _8085;
    wire _8081;
    wire [8:0] _8082;
    wire [8:0] _8086;
    wire [8:0] _8094;
    wire [8:0] _8110;
    wire _8075;
    wire [8:0] _8076;
    wire _8072;
    wire [8:0] _8073;
    wire [8:0] _8077;
    wire _8068;
    wire [8:0] _8069;
    wire _8065;
    wire [8:0] _8066;
    wire [8:0] _8070;
    wire [8:0] _8078;
    wire _8060;
    wire [8:0] _8061;
    wire _8057;
    wire [8:0] _8058;
    wire [8:0] _8062;
    wire _8053;
    wire [8:0] _8054;
    wire _8050;
    wire [8:0] _8051;
    wire [8:0] _8055;
    wire [8:0] _8063;
    wire [8:0] _8079;
    wire [8:0] _8111;
    wire _8043;
    wire [8:0] _8044;
    wire _8040;
    wire [8:0] _8041;
    wire [8:0] _8045;
    wire _8036;
    wire [8:0] _8037;
    wire _8033;
    wire [8:0] _8034;
    wire [8:0] _8038;
    wire [8:0] _8046;
    wire _8028;
    wire [8:0] _8029;
    wire _8025;
    wire [8:0] _8026;
    wire [8:0] _8030;
    wire _8021;
    wire [8:0] _8022;
    wire _8018;
    wire [8:0] _8019;
    wire [8:0] _8023;
    wire [8:0] _8031;
    wire [8:0] _8047;
    wire _8012;
    wire [8:0] _8013;
    wire _8009;
    wire [8:0] _8010;
    wire [8:0] _8014;
    wire _8005;
    wire [8:0] _8006;
    wire _8002;
    wire [8:0] _8003;
    wire [8:0] _8007;
    wire [8:0] _8015;
    wire _7997;
    wire [8:0] _7998;
    wire _7994;
    wire [8:0] _7995;
    wire [8:0] _7999;
    wire _7990;
    wire [8:0] _7991;
    wire _7987;
    wire [8:0] _7988;
    wire [8:0] _7992;
    wire [8:0] _8000;
    wire [8:0] _8016;
    wire [8:0] _8048;
    wire [8:0] _8112;
    wire [8:0] _8240;
    wire _7978;
    wire [8:0] _7979;
    wire _7975;
    wire [8:0] _7976;
    wire [8:0] _7980;
    wire _7971;
    wire [8:0] _7972;
    wire _7968;
    wire [8:0] _7969;
    wire [8:0] _7973;
    wire [8:0] _7981;
    wire _7963;
    wire [8:0] _7964;
    wire _7960;
    wire [8:0] _7961;
    wire [8:0] _7965;
    wire _7956;
    wire [8:0] _7957;
    wire _7953;
    wire [8:0] _7954;
    wire [8:0] _7958;
    wire [8:0] _7966;
    wire [8:0] _7982;
    wire _7947;
    wire [8:0] _7948;
    wire _7944;
    wire [8:0] _7945;
    wire [8:0] _7949;
    wire _7940;
    wire [8:0] _7941;
    wire _7937;
    wire [8:0] _7938;
    wire [8:0] _7942;
    wire [8:0] _7950;
    wire _7932;
    wire [8:0] _7933;
    wire _7929;
    wire [8:0] _7930;
    wire [8:0] _7934;
    wire _7925;
    wire [8:0] _7926;
    wire _7922;
    wire [8:0] _7923;
    wire [8:0] _7927;
    wire [8:0] _7935;
    wire [8:0] _7951;
    wire [8:0] _7983;
    wire _7915;
    wire [8:0] _7916;
    wire _7912;
    wire [8:0] _7913;
    wire [8:0] _7917;
    wire _7908;
    wire [8:0] _7909;
    wire _7905;
    wire [8:0] _7906;
    wire [8:0] _7910;
    wire [8:0] _7918;
    wire _7900;
    wire [8:0] _7901;
    wire _7897;
    wire [8:0] _7898;
    wire [8:0] _7902;
    wire _7893;
    wire [8:0] _7894;
    wire _7890;
    wire [8:0] _7891;
    wire [8:0] _7895;
    wire [8:0] _7903;
    wire [8:0] _7919;
    wire _7884;
    wire [8:0] _7885;
    wire _7881;
    wire [8:0] _7882;
    wire [8:0] _7886;
    wire _7877;
    wire [8:0] _7878;
    wire _7874;
    wire [8:0] _7875;
    wire [8:0] _7879;
    wire [8:0] _7887;
    wire _7869;
    wire [8:0] _7870;
    wire _7866;
    wire [8:0] _7867;
    wire [8:0] _7871;
    wire _7862;
    wire [8:0] _7863;
    wire _7859;
    wire [8:0] _7860;
    wire [8:0] _7864;
    wire [8:0] _7872;
    wire [8:0] _7888;
    wire [8:0] _7920;
    wire [8:0] _7984;
    wire _7851;
    wire [8:0] _7852;
    wire _7848;
    wire [8:0] _7849;
    wire [8:0] _7853;
    wire _7844;
    wire [8:0] _7845;
    wire _7841;
    wire [8:0] _7842;
    wire [8:0] _7846;
    wire [8:0] _7854;
    wire _7836;
    wire [8:0] _7837;
    wire _7833;
    wire [8:0] _7834;
    wire [8:0] _7838;
    wire _7829;
    wire [8:0] _7830;
    wire _7826;
    wire [8:0] _7827;
    wire [8:0] _7831;
    wire [8:0] _7839;
    wire [8:0] _7855;
    wire _7820;
    wire [8:0] _7821;
    wire _7817;
    wire [8:0] _7818;
    wire [8:0] _7822;
    wire _7813;
    wire [8:0] _7814;
    wire _7810;
    wire [8:0] _7811;
    wire [8:0] _7815;
    wire [8:0] _7823;
    wire _7805;
    wire [8:0] _7806;
    wire _7802;
    wire [8:0] _7803;
    wire [8:0] _7807;
    wire _7798;
    wire [8:0] _7799;
    wire _7795;
    wire [8:0] _7796;
    wire [8:0] _7800;
    wire [8:0] _7808;
    wire [8:0] _7824;
    wire [8:0] _7856;
    wire _7788;
    wire [8:0] _7789;
    wire _7785;
    wire [8:0] _7786;
    wire [8:0] _7790;
    wire _7781;
    wire [8:0] _7782;
    wire _7778;
    wire [8:0] _7779;
    wire [8:0] _7783;
    wire [8:0] _7791;
    wire _7773;
    wire [8:0] _7774;
    wire _7770;
    wire [8:0] _7771;
    wire [8:0] _7775;
    wire _7766;
    wire [8:0] _7767;
    wire _7763;
    wire [8:0] _7764;
    wire [8:0] _7768;
    wire [8:0] _7776;
    wire [8:0] _7792;
    wire _7757;
    wire [8:0] _7758;
    wire _7754;
    wire [8:0] _7755;
    wire [8:0] _7759;
    wire _7750;
    wire [8:0] _7751;
    wire _7747;
    wire [8:0] _7748;
    wire [8:0] _7752;
    wire [8:0] _7760;
    wire _7742;
    wire [8:0] _7743;
    wire _7739;
    wire [8:0] _7740;
    wire [8:0] _7744;
    wire _7735;
    wire [8:0] _7736;
    wire _7732;
    wire [8:0] _7733;
    wire [8:0] _7737;
    wire [8:0] _7745;
    wire [8:0] _7761;
    wire [8:0] _7793;
    wire [8:0] _7857;
    wire [8:0] _7985;
    wire [8:0] _8241;
    wire _7722;
    wire [8:0] _7723;
    wire _7719;
    wire [8:0] _7720;
    wire [8:0] _7724;
    wire _7715;
    wire [8:0] _7716;
    wire _7712;
    wire [8:0] _7713;
    wire [8:0] _7717;
    wire [8:0] _7725;
    wire _7707;
    wire [8:0] _7708;
    wire _7704;
    wire [8:0] _7705;
    wire [8:0] _7709;
    wire _7700;
    wire [8:0] _7701;
    wire _7697;
    wire [8:0] _7698;
    wire [8:0] _7702;
    wire [8:0] _7710;
    wire [8:0] _7726;
    wire _7691;
    wire [8:0] _7692;
    wire _7688;
    wire [8:0] _7689;
    wire [8:0] _7693;
    wire _7684;
    wire [8:0] _7685;
    wire _7681;
    wire [8:0] _7682;
    wire [8:0] _7686;
    wire [8:0] _7694;
    wire _7676;
    wire [8:0] _7677;
    wire _7673;
    wire [8:0] _7674;
    wire [8:0] _7678;
    wire _7669;
    wire [8:0] _7670;
    wire _7666;
    wire [8:0] _7667;
    wire [8:0] _7671;
    wire [8:0] _7679;
    wire [8:0] _7695;
    wire [8:0] _7727;
    wire _7659;
    wire [8:0] _7660;
    wire _7656;
    wire [8:0] _7657;
    wire [8:0] _7661;
    wire _7652;
    wire [8:0] _7653;
    wire _7649;
    wire [8:0] _7650;
    wire [8:0] _7654;
    wire [8:0] _7662;
    wire _7644;
    wire [8:0] _7645;
    wire _7641;
    wire [8:0] _7642;
    wire [8:0] _7646;
    wire _7637;
    wire [8:0] _7638;
    wire _7634;
    wire [8:0] _7635;
    wire [8:0] _7639;
    wire [8:0] _7647;
    wire [8:0] _7663;
    wire _7628;
    wire [8:0] _7629;
    wire _7625;
    wire [8:0] _7626;
    wire [8:0] _7630;
    wire _7621;
    wire [8:0] _7622;
    wire _7618;
    wire [8:0] _7619;
    wire [8:0] _7623;
    wire [8:0] _7631;
    wire _7613;
    wire [8:0] _7614;
    wire _7610;
    wire [8:0] _7611;
    wire [8:0] _7615;
    wire _7606;
    wire [8:0] _7607;
    wire _7603;
    wire [8:0] _7604;
    wire [8:0] _7608;
    wire [8:0] _7616;
    wire [8:0] _7632;
    wire [8:0] _7664;
    wire [8:0] _7728;
    wire _7595;
    wire [8:0] _7596;
    wire _7592;
    wire [8:0] _7593;
    wire [8:0] _7597;
    wire _7588;
    wire [8:0] _7589;
    wire _7585;
    wire [8:0] _7586;
    wire [8:0] _7590;
    wire [8:0] _7598;
    wire _7580;
    wire [8:0] _7581;
    wire _7577;
    wire [8:0] _7578;
    wire [8:0] _7582;
    wire _7573;
    wire [8:0] _7574;
    wire _7570;
    wire [8:0] _7571;
    wire [8:0] _7575;
    wire [8:0] _7583;
    wire [8:0] _7599;
    wire _7564;
    wire [8:0] _7565;
    wire _7561;
    wire [8:0] _7562;
    wire [8:0] _7566;
    wire _7557;
    wire [8:0] _7558;
    wire _7554;
    wire [8:0] _7555;
    wire [8:0] _7559;
    wire [8:0] _7567;
    wire _7549;
    wire [8:0] _7550;
    wire _7546;
    wire [8:0] _7547;
    wire [8:0] _7551;
    wire _7542;
    wire [8:0] _7543;
    wire _7539;
    wire [8:0] _7540;
    wire [8:0] _7544;
    wire [8:0] _7552;
    wire [8:0] _7568;
    wire [8:0] _7600;
    wire _7532;
    wire [8:0] _7533;
    wire _7529;
    wire [8:0] _7530;
    wire [8:0] _7534;
    wire _7525;
    wire [8:0] _7526;
    wire _7522;
    wire [8:0] _7523;
    wire [8:0] _7527;
    wire [8:0] _7535;
    wire _7517;
    wire [8:0] _7518;
    wire _7514;
    wire [8:0] _7515;
    wire [8:0] _7519;
    wire _7510;
    wire [8:0] _7511;
    wire _7507;
    wire [8:0] _7508;
    wire [8:0] _7512;
    wire [8:0] _7520;
    wire [8:0] _7536;
    wire _7501;
    wire [8:0] _7502;
    wire _7498;
    wire [8:0] _7499;
    wire [8:0] _7503;
    wire _7494;
    wire [8:0] _7495;
    wire _7491;
    wire [8:0] _7492;
    wire [8:0] _7496;
    wire [8:0] _7504;
    wire _7486;
    wire [8:0] _7487;
    wire _7483;
    wire [8:0] _7484;
    wire [8:0] _7488;
    wire _7479;
    wire [8:0] _7480;
    wire _7476;
    wire [8:0] _7477;
    wire [8:0] _7481;
    wire [8:0] _7489;
    wire [8:0] _7505;
    wire [8:0] _7537;
    wire [8:0] _7601;
    wire [8:0] _7729;
    wire _7467;
    wire [8:0] _7468;
    wire _7464;
    wire [8:0] _7465;
    wire [8:0] _7469;
    wire _7460;
    wire [8:0] _7461;
    wire _7457;
    wire [8:0] _7458;
    wire [8:0] _7462;
    wire [8:0] _7470;
    wire _7452;
    wire [8:0] _7453;
    wire _7449;
    wire [8:0] _7450;
    wire [8:0] _7454;
    wire _7445;
    wire [8:0] _7446;
    wire _7442;
    wire [8:0] _7443;
    wire [8:0] _7447;
    wire [8:0] _7455;
    wire [8:0] _7471;
    wire _7436;
    wire [8:0] _7437;
    wire _7433;
    wire [8:0] _7434;
    wire [8:0] _7438;
    wire _7429;
    wire [8:0] _7430;
    wire _7426;
    wire [8:0] _7427;
    wire [8:0] _7431;
    wire [8:0] _7439;
    wire _7421;
    wire [8:0] _7422;
    wire _7418;
    wire [8:0] _7419;
    wire [8:0] _7423;
    wire _7414;
    wire [8:0] _7415;
    wire _7411;
    wire [8:0] _7412;
    wire [8:0] _7416;
    wire [8:0] _7424;
    wire [8:0] _7440;
    wire [8:0] _7472;
    wire _7404;
    wire [8:0] _7405;
    wire _7401;
    wire [8:0] _7402;
    wire [8:0] _7406;
    wire _7397;
    wire [8:0] _7398;
    wire _7394;
    wire [8:0] _7395;
    wire [8:0] _7399;
    wire [8:0] _7407;
    wire _7389;
    wire [8:0] _7390;
    wire _7386;
    wire [8:0] _7387;
    wire [8:0] _7391;
    wire _7382;
    wire [8:0] _7383;
    wire _7379;
    wire [8:0] _7380;
    wire [8:0] _7384;
    wire [8:0] _7392;
    wire [8:0] _7408;
    wire _7373;
    wire [8:0] _7374;
    wire _7370;
    wire [8:0] _7371;
    wire [8:0] _7375;
    wire _7366;
    wire [8:0] _7367;
    wire _7363;
    wire [8:0] _7364;
    wire [8:0] _7368;
    wire [8:0] _7376;
    wire _7358;
    wire [8:0] _7359;
    wire _7355;
    wire [8:0] _7356;
    wire [8:0] _7360;
    wire _7351;
    wire [8:0] _7352;
    wire _7348;
    wire [8:0] _7349;
    wire [8:0] _7353;
    wire [8:0] _7361;
    wire [8:0] _7377;
    wire [8:0] _7409;
    wire [8:0] _7473;
    wire _7340;
    wire [8:0] _7341;
    wire _7337;
    wire [8:0] _7338;
    wire [8:0] _7342;
    wire _7333;
    wire [8:0] _7334;
    wire _7330;
    wire [8:0] _7331;
    wire [8:0] _7335;
    wire [8:0] _7343;
    wire _7325;
    wire [8:0] _7326;
    wire _7322;
    wire [8:0] _7323;
    wire [8:0] _7327;
    wire _7318;
    wire [8:0] _7319;
    wire _7315;
    wire [8:0] _7316;
    wire [8:0] _7320;
    wire [8:0] _7328;
    wire [8:0] _7344;
    wire _7309;
    wire [8:0] _7310;
    wire _7306;
    wire [8:0] _7307;
    wire [8:0] _7311;
    wire _7302;
    wire [8:0] _7303;
    wire _7299;
    wire [8:0] _7300;
    wire [8:0] _7304;
    wire [8:0] _7312;
    wire _7294;
    wire [8:0] _7295;
    wire _7291;
    wire [8:0] _7292;
    wire [8:0] _7296;
    wire _7287;
    wire [8:0] _7288;
    wire _7284;
    wire [8:0] _7285;
    wire [8:0] _7289;
    wire [8:0] _7297;
    wire [8:0] _7313;
    wire [8:0] _7345;
    wire _7277;
    wire [8:0] _7278;
    wire _7274;
    wire [8:0] _7275;
    wire [8:0] _7279;
    wire _7270;
    wire [8:0] _7271;
    wire _7267;
    wire [8:0] _7268;
    wire [8:0] _7272;
    wire [8:0] _7280;
    wire _7262;
    wire [8:0] _7263;
    wire _7259;
    wire [8:0] _7260;
    wire [8:0] _7264;
    wire _7255;
    wire [8:0] _7256;
    wire _7252;
    wire [8:0] _7253;
    wire [8:0] _7257;
    wire [8:0] _7265;
    wire [8:0] _7281;
    wire _7246;
    wire [8:0] _7247;
    wire _7243;
    wire [8:0] _7244;
    wire [8:0] _7248;
    wire _7239;
    wire [8:0] _7240;
    wire _7236;
    wire [8:0] _7237;
    wire [8:0] _7241;
    wire [8:0] _7249;
    wire _7231;
    wire [8:0] _7232;
    wire _7228;
    wire [8:0] _7229;
    wire [8:0] _7233;
    wire _7224;
    wire [8:0] _7225;
    wire _5396;
    wire _5397;
    wire [63:0] _7212;
    wire [7:0] _7209;
    wire _7210;
    wire [63:0] _7213;
    wire _5376;
    wire _5377;
    wire [7:0] _7202;
    wire _7203;
    wire [63:0] _7206;
    wire [63:0] _5400;
    wire _5356;
    wire _5357;
    wire [7:0] _7195;
    wire _7196;
    wire [63:0] _7199;
    wire [63:0] _5380;
    wire _5336;
    wire _5337;
    wire [7:0] _7188;
    wire _7189;
    wire [63:0] _7192;
    wire [63:0] _5360;
    wire _5316;
    wire _5317;
    wire [7:0] _7181;
    wire _7182;
    wire [63:0] _7185;
    wire [63:0] _5340;
    wire _5296;
    wire _5297;
    wire [7:0] _7174;
    wire _7175;
    wire [63:0] _7178;
    wire [63:0] _5320;
    wire _5276;
    wire _5277;
    wire [7:0] _7167;
    wire _7168;
    wire [63:0] _7171;
    wire [63:0] _5300;
    wire _5256;
    wire _5257;
    wire [7:0] _7160;
    wire _7161;
    wire [63:0] _7164;
    wire [63:0] _5280;
    wire _5236;
    wire _5237;
    wire [7:0] _7153;
    wire _7154;
    wire [63:0] _7157;
    wire [63:0] _5260;
    wire _5216;
    wire _5217;
    wire [7:0] _7146;
    wire _7147;
    wire [63:0] _7150;
    wire [63:0] _5240;
    wire _5196;
    wire _5197;
    wire [7:0] _7139;
    wire _7140;
    wire [63:0] _7143;
    wire [63:0] _5220;
    wire _5176;
    wire _5177;
    wire [7:0] _7132;
    wire _7133;
    wire [63:0] _7136;
    wire [63:0] _5200;
    wire _5156;
    wire _5157;
    wire [7:0] _7125;
    wire _7126;
    wire [63:0] _7129;
    wire [63:0] _5180;
    wire _5136;
    wire _5137;
    wire [7:0] _7118;
    wire _7119;
    wire [63:0] _7122;
    wire [63:0] _5160;
    wire _5116;
    wire _5117;
    wire [7:0] _7111;
    wire _7112;
    wire [63:0] _7115;
    wire [63:0] _5140;
    wire _5096;
    wire _5097;
    wire [7:0] _7104;
    wire _7105;
    wire [63:0] _7108;
    wire [63:0] _5120;
    wire _5076;
    wire _5077;
    wire [7:0] _7097;
    wire _7098;
    wire [63:0] _7101;
    wire [63:0] _5100;
    wire _5056;
    wire _5057;
    wire [7:0] _7090;
    wire _7091;
    wire [63:0] _7094;
    wire [63:0] _5080;
    wire _5036;
    wire _5037;
    wire [7:0] _7083;
    wire _7084;
    wire [63:0] _7087;
    wire [63:0] _5060;
    wire _5016;
    wire _5017;
    wire [7:0] _7076;
    wire _7077;
    wire [63:0] _7080;
    wire [63:0] _5040;
    wire _4996;
    wire _4997;
    wire [7:0] _7069;
    wire _7070;
    wire [63:0] _7073;
    wire [63:0] _5020;
    wire _4976;
    wire _4977;
    wire [7:0] _7062;
    wire _7063;
    wire [63:0] _7066;
    wire [63:0] _5000;
    wire _4956;
    wire _4957;
    wire [7:0] _7055;
    wire _7056;
    wire [63:0] _7059;
    wire [63:0] _4980;
    wire _4936;
    wire _4937;
    wire [7:0] _7048;
    wire _7049;
    wire [63:0] _7052;
    wire [63:0] _4960;
    wire _4916;
    wire _4917;
    wire [7:0] _7041;
    wire _7042;
    wire [63:0] _7045;
    wire [63:0] _4940;
    wire _4896;
    wire _4897;
    wire [7:0] _7034;
    wire _7035;
    wire [63:0] _7038;
    wire [63:0] _4920;
    wire _4876;
    wire _4877;
    wire [7:0] _7027;
    wire _7028;
    wire [63:0] _7031;
    wire [63:0] _4900;
    wire _4856;
    wire _4857;
    wire [7:0] _7020;
    wire _7021;
    wire [63:0] _7024;
    wire [63:0] _4880;
    wire _4836;
    wire _4837;
    wire [7:0] _7013;
    wire _7014;
    wire [63:0] _7017;
    wire [63:0] _4860;
    wire _4816;
    wire _4817;
    wire [7:0] _7006;
    wire _7007;
    wire [63:0] _7010;
    wire [63:0] _4840;
    wire _4796;
    wire _4797;
    wire [7:0] _6999;
    wire _7000;
    wire [63:0] _7003;
    wire [63:0] _4820;
    wire _4776;
    wire _4777;
    wire [7:0] _6992;
    wire _6993;
    wire [63:0] _6996;
    wire [63:0] _4800;
    wire _4756;
    wire _4757;
    wire [7:0] _6985;
    wire _6986;
    wire [63:0] _6989;
    wire [63:0] _4780;
    wire _4736;
    wire _4737;
    wire [7:0] _6978;
    wire _6979;
    wire [63:0] _6982;
    wire [63:0] _4760;
    wire _4716;
    wire _4717;
    wire [7:0] _6971;
    wire _6972;
    wire [63:0] _6975;
    wire [63:0] _4740;
    wire _4696;
    wire _4697;
    wire [7:0] _6964;
    wire _6965;
    wire [63:0] _6968;
    wire [63:0] _4720;
    wire _4676;
    wire _4677;
    wire [7:0] _6957;
    wire _6958;
    wire [63:0] _6961;
    wire [63:0] _4700;
    wire _4656;
    wire _4657;
    wire [7:0] _6950;
    wire _6951;
    wire [63:0] _6954;
    wire [63:0] _4680;
    wire _4636;
    wire _4637;
    wire [7:0] _6943;
    wire _6944;
    wire [63:0] _6947;
    wire [63:0] _4660;
    wire _4616;
    wire _4617;
    wire [7:0] _6936;
    wire _6937;
    wire [63:0] _6940;
    wire [63:0] _4640;
    wire _4596;
    wire _4597;
    wire [7:0] _6929;
    wire _6930;
    wire [63:0] _6933;
    wire [63:0] _4620;
    wire _4576;
    wire _4577;
    wire [7:0] _6922;
    wire _6923;
    wire [63:0] _6926;
    wire [63:0] _4600;
    wire _4556;
    wire _4557;
    wire [7:0] _6915;
    wire _6916;
    wire [63:0] _6919;
    wire [63:0] _4580;
    wire _4536;
    wire _4537;
    wire [7:0] _6908;
    wire _6909;
    wire [63:0] _6912;
    wire [63:0] _4560;
    wire _4516;
    wire _4517;
    wire [7:0] _6901;
    wire _6902;
    wire [63:0] _6905;
    wire [63:0] _4540;
    wire _4496;
    wire _4497;
    wire [7:0] _6894;
    wire _6895;
    wire [63:0] _6898;
    wire [63:0] _4520;
    wire _4476;
    wire _4477;
    wire [7:0] _6887;
    wire _6888;
    wire [63:0] _6891;
    wire [63:0] _4500;
    wire _4456;
    wire _4457;
    wire [7:0] _6880;
    wire _6881;
    wire [63:0] _6884;
    wire [63:0] _4480;
    wire _4436;
    wire _4437;
    wire [7:0] _6873;
    wire _6874;
    wire [63:0] _6877;
    wire [63:0] _4460;
    wire _4416;
    wire _4417;
    wire [7:0] _6866;
    wire _6867;
    wire [63:0] _6870;
    wire [63:0] _4440;
    wire _4396;
    wire _4397;
    wire [7:0] _6859;
    wire _6860;
    wire [63:0] _6863;
    wire [63:0] _4420;
    wire _4376;
    wire _4377;
    wire [7:0] _6852;
    wire _6853;
    wire [63:0] _6856;
    wire [63:0] _4400;
    wire _4356;
    wire _4357;
    wire [7:0] _6845;
    wire _6846;
    wire [63:0] _6849;
    wire [63:0] _4380;
    wire _4336;
    wire _4337;
    wire [7:0] _6838;
    wire _6839;
    wire [63:0] _6842;
    wire [63:0] _4360;
    wire _4316;
    wire _4317;
    wire [7:0] _6831;
    wire _6832;
    wire [63:0] _6835;
    wire [63:0] _4340;
    wire _4296;
    wire _4297;
    wire [7:0] _6824;
    wire _6825;
    wire [63:0] _6828;
    wire [63:0] _4320;
    wire _4276;
    wire _4277;
    wire [7:0] _6817;
    wire _6818;
    wire [63:0] _6821;
    wire [63:0] _4300;
    wire _4256;
    wire _4257;
    wire [7:0] _6810;
    wire _6811;
    wire [63:0] _6814;
    wire [63:0] _4280;
    wire _4236;
    wire _4237;
    wire [7:0] _6803;
    wire _6804;
    wire [63:0] _6807;
    wire [63:0] _4260;
    wire _4216;
    wire _4217;
    wire [7:0] _6796;
    wire _6797;
    wire [63:0] _6800;
    wire [63:0] _4240;
    wire _4196;
    wire _4197;
    wire [7:0] _6789;
    wire _6790;
    wire [63:0] _6793;
    wire [63:0] _4220;
    wire _4176;
    wire _4177;
    wire [7:0] _6782;
    wire _6783;
    wire [63:0] _6786;
    wire [63:0] _4200;
    wire _4156;
    wire _4157;
    wire [7:0] _6775;
    wire _6776;
    wire [63:0] _6779;
    wire [63:0] _4180;
    wire _4136;
    wire _4137;
    wire [7:0] _6768;
    wire _6769;
    wire [63:0] _6772;
    wire [63:0] _4160;
    wire _4116;
    wire _4117;
    wire [7:0] _6761;
    wire _6762;
    wire [63:0] _6765;
    wire [63:0] _4140;
    wire _4096;
    wire _4097;
    wire [7:0] _6754;
    wire _6755;
    wire [63:0] _6758;
    wire [63:0] _4120;
    wire _4076;
    wire _4077;
    wire [7:0] _6747;
    wire _6748;
    wire [63:0] _6751;
    wire [63:0] _4100;
    wire _4056;
    wire _4057;
    wire [7:0] _6740;
    wire _6741;
    wire [63:0] _6744;
    wire [63:0] _4080;
    wire _4036;
    wire _4037;
    wire [7:0] _6733;
    wire _6734;
    wire [63:0] _6737;
    wire [63:0] _4060;
    wire _4016;
    wire _4017;
    wire [7:0] _6726;
    wire _6727;
    wire [63:0] _6730;
    wire [63:0] _4040;
    wire _3996;
    wire _3997;
    wire [7:0] _6719;
    wire _6720;
    wire [63:0] _6723;
    wire [63:0] _4020;
    wire _3976;
    wire _3977;
    wire [7:0] _6712;
    wire _6713;
    wire [63:0] _6716;
    wire [63:0] _4000;
    wire _3956;
    wire _3957;
    wire [7:0] _6705;
    wire _6706;
    wire [63:0] _6709;
    wire [63:0] _3980;
    wire _3936;
    wire _3937;
    wire [7:0] _6698;
    wire _6699;
    wire [63:0] _6702;
    wire [63:0] _3960;
    wire _3916;
    wire _3917;
    wire [7:0] _6691;
    wire _6692;
    wire [63:0] _6695;
    wire [63:0] _3940;
    wire _3896;
    wire _3897;
    wire [7:0] _6684;
    wire _6685;
    wire [63:0] _6688;
    wire [63:0] _3920;
    wire _3876;
    wire _3877;
    wire [7:0] _6677;
    wire _6678;
    wire [63:0] _6681;
    wire [63:0] _3900;
    wire _3856;
    wire _3857;
    wire [7:0] _6670;
    wire _6671;
    wire [63:0] _6674;
    wire [63:0] _3880;
    wire _3836;
    wire _3837;
    wire [7:0] _6663;
    wire _6664;
    wire [63:0] _6667;
    wire [63:0] _3860;
    wire _3816;
    wire _3817;
    wire [7:0] _6656;
    wire _6657;
    wire [63:0] _6660;
    wire [63:0] _3840;
    wire _3796;
    wire _3797;
    wire [7:0] _6649;
    wire _6650;
    wire [63:0] _6653;
    wire [63:0] _3820;
    wire _3776;
    wire _3777;
    wire [7:0] _6642;
    wire _6643;
    wire [63:0] _6646;
    wire [63:0] _3800;
    wire _3756;
    wire _3757;
    wire [7:0] _6635;
    wire _6636;
    wire [63:0] _6639;
    wire [63:0] _3780;
    wire _3736;
    wire _3737;
    wire [7:0] _6628;
    wire _6629;
    wire [63:0] _6632;
    wire [63:0] _3760;
    wire _3716;
    wire _3717;
    wire [7:0] _6621;
    wire _6622;
    wire [63:0] _6625;
    wire [63:0] _3740;
    wire _3696;
    wire _3697;
    wire [7:0] _6614;
    wire _6615;
    wire [63:0] _6618;
    wire [63:0] _3720;
    wire _3676;
    wire _3677;
    wire [7:0] _6607;
    wire _6608;
    wire [63:0] _6611;
    wire [63:0] _3700;
    wire _3656;
    wire _3657;
    wire [7:0] _6600;
    wire _6601;
    wire [63:0] _6604;
    wire [63:0] _3680;
    wire _3636;
    wire _3637;
    wire [7:0] _6593;
    wire _6594;
    wire [63:0] _6597;
    wire [63:0] _3660;
    wire _3616;
    wire _3617;
    wire [7:0] _6586;
    wire _6587;
    wire [63:0] _6590;
    wire [63:0] _3640;
    wire _3596;
    wire _3597;
    wire [7:0] _6579;
    wire _6580;
    wire [63:0] _6583;
    wire [63:0] _3620;
    wire _3576;
    wire _3577;
    wire [7:0] _6572;
    wire _6573;
    wire [63:0] _6576;
    wire [63:0] _3600;
    wire _3556;
    wire _3557;
    wire [7:0] _6565;
    wire _6566;
    wire [63:0] _6569;
    wire [63:0] _3580;
    wire _3536;
    wire _3537;
    wire [7:0] _6558;
    wire _6559;
    wire [63:0] _6562;
    wire [63:0] _3560;
    wire _3516;
    wire _3517;
    wire [7:0] _6551;
    wire _6552;
    wire [63:0] _6555;
    wire [63:0] _3540;
    wire _3496;
    wire _3497;
    wire [7:0] _6544;
    wire _6545;
    wire [63:0] _6548;
    wire [63:0] _3520;
    wire _3476;
    wire _3477;
    wire [7:0] _6537;
    wire _6538;
    wire [63:0] _6541;
    wire [63:0] _3500;
    wire _3456;
    wire _3457;
    wire [7:0] _6530;
    wire _6531;
    wire [63:0] _6534;
    wire [63:0] _3480;
    wire _3436;
    wire _3437;
    wire [7:0] _6523;
    wire _6524;
    wire [63:0] _6527;
    wire [63:0] _3460;
    wire _3416;
    wire _3417;
    wire [7:0] _6516;
    wire _6517;
    wire [63:0] _6520;
    wire [63:0] _3440;
    wire _3396;
    wire _3397;
    wire [7:0] _6509;
    wire _6510;
    wire [63:0] _6513;
    wire [63:0] _3420;
    wire _3376;
    wire _3377;
    wire [7:0] _6502;
    wire _6503;
    wire [63:0] _6506;
    wire [63:0] _3400;
    wire _3356;
    wire _3357;
    wire [7:0] _6495;
    wire _6496;
    wire [63:0] _6499;
    wire [63:0] _3380;
    wire _3336;
    wire _3337;
    wire [7:0] _6488;
    wire _6489;
    wire [63:0] _6492;
    wire [63:0] _3360;
    wire _3316;
    wire _3317;
    wire [7:0] _6481;
    wire _6482;
    wire [63:0] _6485;
    wire [63:0] _3340;
    wire _3296;
    wire _3297;
    wire [7:0] _6474;
    wire _6475;
    wire [63:0] _6478;
    wire [63:0] _3320;
    wire _3276;
    wire _3277;
    wire [7:0] _6467;
    wire _6468;
    wire [63:0] _6471;
    wire [63:0] _3300;
    wire _3256;
    wire _3257;
    wire [7:0] _6460;
    wire _6461;
    wire [63:0] _6464;
    wire [63:0] _3280;
    wire _3236;
    wire _3237;
    wire [7:0] _6453;
    wire _6454;
    wire [63:0] _6457;
    wire [63:0] _3260;
    wire _3216;
    wire _3217;
    wire [7:0] _6446;
    wire _6447;
    wire [63:0] _6450;
    wire [63:0] _3240;
    wire _3196;
    wire _3197;
    wire [7:0] _6439;
    wire _6440;
    wire [63:0] _6443;
    wire [63:0] _3220;
    wire _3176;
    wire _3177;
    wire [7:0] _6432;
    wire _6433;
    wire [63:0] _6436;
    wire [63:0] _3200;
    wire _3156;
    wire _3157;
    wire [7:0] _6425;
    wire _6426;
    wire [63:0] _6429;
    wire [63:0] _3180;
    wire _3136;
    wire _3137;
    wire [7:0] _6418;
    wire _6419;
    wire [63:0] _6422;
    wire [63:0] _3160;
    wire _3116;
    wire _3117;
    wire [7:0] _6411;
    wire _6412;
    wire [63:0] _6415;
    wire [63:0] _3140;
    wire _3096;
    wire _3097;
    wire [7:0] _6404;
    wire _6405;
    wire [63:0] _6408;
    wire [63:0] _3120;
    wire _3076;
    wire _3077;
    wire [7:0] _6397;
    wire _6398;
    wire [63:0] _6401;
    wire [63:0] _3100;
    wire _3056;
    wire _3057;
    wire [7:0] _6390;
    wire _6391;
    wire [63:0] _6394;
    wire [63:0] _3080;
    wire _3036;
    wire _3037;
    wire [7:0] _6383;
    wire _6384;
    wire [63:0] _6387;
    wire [63:0] _3060;
    wire _3016;
    wire _3017;
    wire [7:0] _6376;
    wire _6377;
    wire [63:0] _6380;
    wire [63:0] _3040;
    wire _2996;
    wire _2997;
    wire [7:0] _6369;
    wire _6370;
    wire [63:0] _6373;
    wire [63:0] _3020;
    wire _2976;
    wire _2977;
    wire [7:0] _6362;
    wire _6363;
    wire [63:0] _6366;
    wire [63:0] _3000;
    wire _2956;
    wire _2957;
    wire [7:0] _6355;
    wire _6356;
    wire [63:0] _6359;
    wire [63:0] _2980;
    wire _2936;
    wire _2937;
    wire [7:0] _6348;
    wire _6349;
    wire [63:0] _6352;
    wire [63:0] _2960;
    wire _2916;
    wire _2917;
    wire [7:0] _6341;
    wire _6342;
    wire [63:0] _6345;
    wire [63:0] _2940;
    wire _2896;
    wire _2897;
    wire [7:0] _6334;
    wire _6335;
    wire [63:0] _6338;
    wire [63:0] _2920;
    wire _2876;
    wire _2877;
    wire [7:0] _6327;
    wire _6328;
    wire [63:0] _6331;
    wire [63:0] _2900;
    wire _2856;
    wire _2857;
    wire [7:0] _6320;
    wire _6321;
    wire [63:0] _6324;
    wire [63:0] _2880;
    wire _2836;
    wire _2837;
    wire [7:0] _6313;
    wire _6314;
    wire [63:0] _6317;
    wire [63:0] _2860;
    wire _2816;
    wire _2817;
    wire [7:0] _6306;
    wire _6307;
    wire [63:0] _6310;
    wire [63:0] _2840;
    wire _2796;
    wire _2797;
    wire [7:0] _6299;
    wire _6300;
    wire [63:0] _6303;
    wire [63:0] _2820;
    wire _2776;
    wire _2777;
    wire [7:0] _6292;
    wire _6293;
    wire [63:0] _6296;
    wire [63:0] _2800;
    wire _2756;
    wire _2757;
    wire [7:0] _6285;
    wire _6286;
    wire [63:0] _6289;
    wire [63:0] _2780;
    wire _2736;
    wire _2737;
    wire [7:0] _6278;
    wire _6279;
    wire [63:0] _6282;
    wire [63:0] _2760;
    wire _2716;
    wire _2717;
    wire [7:0] _6271;
    wire _6272;
    wire [63:0] _6275;
    wire [63:0] _2740;
    wire _2696;
    wire _2697;
    wire [7:0] _6264;
    wire _6265;
    wire [63:0] _6268;
    wire [63:0] _2720;
    wire _2676;
    wire _2677;
    wire [7:0] _6257;
    wire _6258;
    wire [63:0] _6261;
    wire [63:0] _2700;
    wire _2656;
    wire _2657;
    wire [7:0] _6250;
    wire _6251;
    wire [63:0] _6254;
    wire [63:0] _2680;
    wire _2636;
    wire _2637;
    wire [7:0] _6243;
    wire _6244;
    wire [63:0] _6247;
    wire [63:0] _2660;
    wire _2616;
    wire _2617;
    wire [7:0] _6236;
    wire _6237;
    wire [63:0] _6240;
    wire [63:0] _2640;
    wire _2596;
    wire _2597;
    wire [7:0] _6229;
    wire _6230;
    wire [63:0] _6233;
    wire [63:0] _2620;
    wire _2576;
    wire _2577;
    wire [7:0] _6222;
    wire _6223;
    wire [63:0] _6226;
    wire [63:0] _2600;
    wire _2556;
    wire _2557;
    wire [7:0] _6215;
    wire _6216;
    wire [63:0] _6219;
    wire [63:0] _2580;
    wire _2536;
    wire _2537;
    wire [7:0] _6208;
    wire _6209;
    wire [63:0] _6212;
    wire [63:0] _2560;
    wire _2516;
    wire _2517;
    wire [7:0] _6201;
    wire _6202;
    wire [63:0] _6205;
    wire [63:0] _2540;
    wire _2496;
    wire _2497;
    wire [7:0] _6194;
    wire _6195;
    wire [63:0] _6198;
    wire [63:0] _2520;
    wire _2476;
    wire _2477;
    wire [7:0] _6187;
    wire _6188;
    wire [63:0] _6191;
    wire [63:0] _2500;
    wire _2456;
    wire _2457;
    wire [7:0] _6180;
    wire _6181;
    wire [63:0] _6184;
    wire [63:0] _2480;
    wire _2436;
    wire _2437;
    wire [7:0] _6173;
    wire _6174;
    wire [63:0] _6177;
    wire [63:0] _2460;
    wire _2416;
    wire _2417;
    wire [7:0] _6166;
    wire _6167;
    wire [63:0] _6170;
    wire [63:0] _2440;
    wire _2396;
    wire _2397;
    wire [7:0] _6159;
    wire _6160;
    wire [63:0] _6163;
    wire [63:0] _2420;
    wire _2376;
    wire _2377;
    wire [7:0] _6152;
    wire _6153;
    wire [63:0] _6156;
    wire [63:0] _2400;
    wire _2356;
    wire _2357;
    wire [7:0] _6145;
    wire _6146;
    wire [63:0] _6149;
    wire [63:0] _2380;
    wire _2336;
    wire _2337;
    wire [7:0] _6138;
    wire _6139;
    wire [63:0] _6142;
    wire [63:0] _2360;
    wire _2316;
    wire _2317;
    wire [7:0] _6131;
    wire _6132;
    wire [63:0] _6135;
    wire [63:0] _2340;
    wire _2296;
    wire _2297;
    wire [7:0] _6124;
    wire _6125;
    wire [63:0] _6128;
    wire [63:0] _2320;
    wire _2276;
    wire _2277;
    wire [7:0] _6117;
    wire _6118;
    wire [63:0] _6121;
    wire [63:0] _2300;
    wire _2256;
    wire _2257;
    wire [7:0] _6110;
    wire _6111;
    wire [63:0] _6114;
    wire [63:0] _2280;
    wire _2236;
    wire _2237;
    wire [7:0] _6103;
    wire _6104;
    wire [63:0] _6107;
    wire [63:0] _2260;
    wire _2216;
    wire _2217;
    wire [7:0] _6096;
    wire _6097;
    wire [63:0] _6100;
    wire [63:0] _2240;
    wire _2196;
    wire _2197;
    wire [7:0] _6089;
    wire _6090;
    wire [63:0] _6093;
    wire [63:0] _2220;
    wire _2176;
    wire _2177;
    wire [7:0] _6082;
    wire _6083;
    wire [63:0] _6086;
    wire [63:0] _2200;
    wire _2156;
    wire _2157;
    wire [7:0] _6075;
    wire _6076;
    wire [63:0] _6079;
    wire [63:0] _2180;
    wire _2136;
    wire _2137;
    wire [7:0] _6068;
    wire _6069;
    wire [63:0] _6072;
    wire [63:0] _2160;
    wire _2116;
    wire _2117;
    wire [7:0] _6061;
    wire _6062;
    wire [63:0] _6065;
    wire [63:0] _2140;
    wire _2096;
    wire _2097;
    wire [7:0] _6054;
    wire _6055;
    wire [63:0] _6058;
    wire [63:0] _2120;
    wire _2076;
    wire _2077;
    wire [7:0] _6047;
    wire _6048;
    wire [63:0] _6051;
    wire [63:0] _2100;
    wire _2056;
    wire _2057;
    wire [7:0] _6040;
    wire _6041;
    wire [63:0] _6044;
    wire [63:0] _2080;
    wire _2036;
    wire _2037;
    wire [7:0] _6033;
    wire _6034;
    wire [63:0] _6037;
    wire [63:0] _2060;
    wire _2016;
    wire _2017;
    wire [7:0] _6026;
    wire _6027;
    wire [63:0] _6030;
    wire [63:0] _2040;
    wire _1996;
    wire _1997;
    wire [7:0] _6019;
    wire _6020;
    wire [63:0] _6023;
    wire [63:0] _2020;
    wire _1976;
    wire _1977;
    wire [7:0] _6012;
    wire _6013;
    wire [63:0] _6016;
    wire [63:0] _2000;
    wire _1956;
    wire _1957;
    wire [7:0] _6005;
    wire _6006;
    wire [63:0] _6009;
    wire [63:0] _1980;
    wire _1936;
    wire _1937;
    wire [7:0] _5998;
    wire _5999;
    wire [63:0] _6002;
    wire [63:0] _1960;
    wire _1916;
    wire _1917;
    wire [7:0] _5991;
    wire _5992;
    wire [63:0] _5995;
    wire [63:0] _1940;
    wire _1896;
    wire _1897;
    wire [7:0] _5984;
    wire _5985;
    wire [63:0] _5988;
    wire [63:0] _1920;
    wire _1876;
    wire _1877;
    wire [7:0] _5977;
    wire _5978;
    wire [63:0] _5981;
    wire [63:0] _1900;
    wire _1856;
    wire _1857;
    wire [7:0] _5970;
    wire _5971;
    wire [63:0] _5974;
    wire [63:0] _1880;
    wire _1836;
    wire _1837;
    wire [7:0] _5963;
    wire _5964;
    wire [63:0] _5967;
    wire [63:0] _1860;
    wire _1816;
    wire _1817;
    wire [7:0] _5956;
    wire _5957;
    wire [63:0] _5960;
    wire [63:0] _1840;
    wire _1796;
    wire _1797;
    wire [7:0] _5949;
    wire _5950;
    wire [63:0] _5953;
    wire [63:0] _1820;
    wire _1776;
    wire _1777;
    wire [7:0] _5942;
    wire _5943;
    wire [63:0] _5946;
    wire [63:0] _1800;
    wire _1756;
    wire _1757;
    wire [7:0] _5935;
    wire _5936;
    wire [63:0] _5939;
    wire [63:0] _1780;
    wire _1736;
    wire _1737;
    wire [7:0] _5928;
    wire _5929;
    wire [63:0] _5932;
    wire [63:0] _1760;
    wire _1716;
    wire _1717;
    wire [7:0] _5921;
    wire _5922;
    wire [63:0] _5925;
    wire [63:0] _1740;
    wire _1696;
    wire _1697;
    wire [7:0] _5914;
    wire _5915;
    wire [63:0] _5918;
    wire [63:0] _1720;
    wire _1676;
    wire _1677;
    wire [7:0] _5907;
    wire _5908;
    wire [63:0] _5911;
    wire [63:0] _1700;
    wire _1656;
    wire _1657;
    wire [7:0] _5900;
    wire _5901;
    wire [63:0] _5904;
    wire [63:0] _1680;
    wire _1636;
    wire _1637;
    wire [7:0] _5893;
    wire _5894;
    wire [63:0] _5897;
    wire [63:0] _1660;
    wire _1616;
    wire _1617;
    wire [7:0] _5886;
    wire _5887;
    wire [63:0] _5890;
    wire [63:0] _1640;
    wire _1596;
    wire _1597;
    wire [7:0] _5879;
    wire _5880;
    wire [63:0] _5883;
    wire [63:0] _1620;
    wire _1576;
    wire _1577;
    wire [7:0] _5872;
    wire _5873;
    wire [63:0] _5876;
    wire [63:0] _1600;
    wire _1556;
    wire _1557;
    wire [7:0] _5865;
    wire _5866;
    wire [63:0] _5869;
    wire [63:0] _1580;
    wire _1536;
    wire _1537;
    wire [7:0] _5858;
    wire _5859;
    wire [63:0] _5862;
    wire [63:0] _1560;
    wire _1516;
    wire _1517;
    wire [7:0] _5851;
    wire _5852;
    wire [63:0] _5855;
    wire [63:0] _1540;
    wire _1496;
    wire _1497;
    wire [7:0] _5844;
    wire _5845;
    wire [63:0] _5848;
    wire [63:0] _1520;
    wire _1476;
    wire _1477;
    wire [7:0] _5837;
    wire _5838;
    wire [63:0] _5841;
    wire [63:0] _1500;
    wire _1456;
    wire _1457;
    wire [7:0] _5830;
    wire _5831;
    wire [63:0] _5834;
    wire [63:0] _1480;
    wire _1436;
    wire _1437;
    wire [7:0] _5823;
    wire _5824;
    wire [63:0] _5827;
    wire [63:0] _1460;
    wire _1416;
    wire _1417;
    wire [7:0] _5816;
    wire _5817;
    wire [63:0] _5820;
    wire [63:0] _1440;
    wire _1396;
    wire _1397;
    wire [7:0] _5809;
    wire _5810;
    wire [63:0] _5813;
    wire [63:0] _1420;
    wire _1376;
    wire _1377;
    wire [7:0] _5802;
    wire _5803;
    wire [63:0] _5806;
    wire [63:0] _1400;
    wire _1356;
    wire _1357;
    wire [7:0] _5795;
    wire _5796;
    wire [63:0] _5799;
    wire [63:0] _1380;
    wire _1336;
    wire _1337;
    wire [7:0] _5788;
    wire _5789;
    wire [63:0] _5792;
    wire [63:0] _1360;
    wire _1316;
    wire _1317;
    wire [7:0] _5781;
    wire _5782;
    wire [63:0] _5785;
    wire [63:0] _1340;
    wire _1296;
    wire _1297;
    wire [7:0] _5774;
    wire _5775;
    wire [63:0] _5778;
    wire [63:0] _1320;
    wire _1276;
    wire _1277;
    wire [7:0] _5767;
    wire _5768;
    wire [63:0] _5771;
    wire [63:0] _1300;
    wire _1256;
    wire _1257;
    wire [7:0] _5760;
    wire _5761;
    wire [63:0] _5764;
    wire [63:0] _1280;
    wire _1236;
    wire _1237;
    wire [7:0] _5753;
    wire _5754;
    wire [63:0] _5757;
    wire [63:0] _1260;
    wire _1216;
    wire _1217;
    wire [7:0] _5746;
    wire _5747;
    wire [63:0] _5750;
    wire [63:0] _1240;
    wire _1196;
    wire _1197;
    wire [7:0] _5739;
    wire _5740;
    wire [63:0] _5743;
    wire [63:0] _1220;
    wire _1176;
    wire _1177;
    wire [7:0] _5732;
    wire _5733;
    wire [63:0] _5736;
    wire [63:0] _1200;
    wire _1156;
    wire _1157;
    wire [7:0] _5725;
    wire _5726;
    wire [63:0] _5729;
    wire [63:0] _1180;
    wire _1136;
    wire _1137;
    wire [7:0] _5718;
    wire _5719;
    wire [63:0] _5722;
    wire [63:0] _1160;
    wire _1116;
    wire _1117;
    wire [7:0] _5711;
    wire _5712;
    wire [63:0] _5715;
    wire [63:0] _1140;
    wire _1096;
    wire _1097;
    wire [7:0] _5704;
    wire _5705;
    wire [63:0] _5708;
    wire [63:0] _1120;
    wire _1076;
    wire _1077;
    wire [7:0] _5697;
    wire _5698;
    wire [63:0] _5701;
    wire [63:0] _1100;
    wire _1056;
    wire _1057;
    wire [7:0] _5690;
    wire _5691;
    wire [63:0] _5694;
    wire [63:0] _1080;
    wire _1036;
    wire _1037;
    wire [7:0] _5683;
    wire _5684;
    wire [63:0] _5687;
    wire [63:0] _1060;
    wire _1016;
    wire _1017;
    wire [7:0] _5676;
    wire _5677;
    wire [63:0] _5680;
    wire [63:0] _1040;
    wire _996;
    wire _997;
    wire [7:0] _5669;
    wire _5670;
    wire [63:0] _5673;
    wire [63:0] _1020;
    wire _976;
    wire _977;
    wire [7:0] _5662;
    wire _5663;
    wire [63:0] _5666;
    wire [63:0] _1000;
    wire _956;
    wire _957;
    wire [7:0] _5655;
    wire _5656;
    wire [63:0] _5659;
    wire [63:0] _980;
    wire _936;
    wire _937;
    wire [7:0] _5648;
    wire _5649;
    wire [63:0] _5652;
    wire [63:0] _960;
    wire _916;
    wire _917;
    wire [7:0] _5641;
    wire _5642;
    wire [63:0] _5645;
    wire [63:0] _940;
    wire _896;
    wire _897;
    wire [7:0] _5634;
    wire _5635;
    wire [63:0] _5638;
    wire [63:0] _920;
    wire _876;
    wire _877;
    wire [7:0] _5627;
    wire _5628;
    wire [63:0] _5631;
    wire [63:0] _900;
    wire _856;
    wire _857;
    wire [7:0] _5620;
    wire _5621;
    wire [63:0] _5624;
    wire [63:0] _880;
    wire _836;
    wire _837;
    wire [7:0] _5613;
    wire _5614;
    wire [63:0] _5617;
    wire [63:0] _860;
    wire _816;
    wire _817;
    wire [7:0] _5606;
    wire _5607;
    wire [63:0] _5610;
    wire [63:0] _840;
    wire _796;
    wire _797;
    wire [7:0] _5599;
    wire _5600;
    wire [63:0] _5603;
    wire [63:0] _820;
    wire _776;
    wire _777;
    wire [7:0] _5592;
    wire _5593;
    wire [63:0] _5596;
    wire [63:0] _800;
    wire _756;
    wire _757;
    wire [7:0] _5585;
    wire _5586;
    wire [63:0] _5589;
    wire [63:0] _780;
    wire _736;
    wire _737;
    wire [7:0] _5578;
    wire _5579;
    wire [63:0] _5582;
    wire [63:0] _760;
    wire _716;
    wire _717;
    wire [7:0] _5571;
    wire _5572;
    wire [63:0] _5575;
    wire [63:0] _740;
    wire _696;
    wire _697;
    wire [7:0] _5564;
    wire _5565;
    wire [63:0] _5568;
    wire [63:0] _720;
    wire _676;
    wire _677;
    wire [7:0] _5557;
    wire _5558;
    wire [63:0] _5561;
    wire [63:0] _700;
    wire _656;
    wire _657;
    wire [7:0] _5550;
    wire _5551;
    wire [63:0] _5554;
    wire [63:0] _680;
    wire _636;
    wire _637;
    wire [7:0] _5543;
    wire _5544;
    wire [63:0] _5547;
    wire [63:0] _660;
    wire _616;
    wire _617;
    wire [7:0] _5536;
    wire _5537;
    wire [63:0] _5540;
    wire [63:0] _640;
    wire _596;
    wire _597;
    wire [7:0] _5529;
    wire _5530;
    wire [63:0] _5533;
    wire [63:0] _620;
    wire _576;
    wire _577;
    wire [7:0] _5522;
    wire _5523;
    wire [63:0] _5526;
    wire [63:0] _600;
    wire _556;
    wire _557;
    wire [7:0] _5515;
    wire _5516;
    wire [63:0] _5519;
    wire [63:0] _580;
    wire _536;
    wire _537;
    wire [7:0] _5508;
    wire _5509;
    wire [63:0] _5512;
    wire [63:0] _560;
    wire _516;
    wire _517;
    wire [7:0] _5501;
    wire _5502;
    wire [63:0] _5505;
    wire [63:0] _540;
    wire _496;
    wire _497;
    wire [7:0] _5494;
    wire _5495;
    wire [63:0] _5498;
    wire [63:0] _520;
    wire _476;
    wire _477;
    wire [7:0] _5487;
    wire _5488;
    wire [63:0] _5491;
    wire [63:0] _500;
    wire _456;
    wire _457;
    wire [7:0] _5480;
    wire _5481;
    wire [63:0] _5484;
    wire [63:0] _480;
    wire _436;
    wire _437;
    wire [7:0] _5473;
    wire _5474;
    wire [63:0] _5477;
    wire [63:0] _460;
    wire _416;
    wire _417;
    wire [7:0] _5466;
    wire _5467;
    wire [63:0] _5470;
    wire [63:0] _440;
    wire _396;
    wire _397;
    wire [7:0] _5459;
    wire _5460;
    wire [63:0] _5463;
    wire [63:0] _420;
    wire _376;
    wire _377;
    wire [7:0] _5452;
    wire _5453;
    wire [63:0] _5456;
    wire [63:0] _400;
    wire _356;
    wire _357;
    wire [7:0] _5445;
    wire _5446;
    wire [63:0] _5449;
    wire [63:0] _380;
    wire _336;
    wire _337;
    wire [7:0] _5438;
    wire _5439;
    wire [63:0] _5442;
    wire [63:0] _360;
    wire _317;
    wire _318;
    wire [7:0] _5431;
    wire _5432;
    wire [63:0] _5435;
    wire [63:0] _340;
    wire _302;
    wire _5414;
    wire _5412;
    wire _5413;
    wire _5415;
    wire _4;
    reg _303;
    wire gnd;
    wire _304;
    wire _305;
    wire [7:0] _6;
    wire [6:0] _5420;
    wire [7:0] _5421;
    reg [7:0] _5418;
    wire [7:0] _5422;
    wire [7:0] _7;
    wire _5425;
    wire [63:0] _5428;
    wire [63:0] _321;
    wire [63:0] _308;
    wire [63:0] _322;
    wire [63:0] _5423;
    wire [63:0] _5429;
    wire [63:0] _8;
    reg [63:0] _295;
    wire _297;
    wire _298;
    wire _292;
    wire _299;
    wire _306;
    wire [63:0] _326;
    wire [63:0] _324;
    wire [63:0] _327;
    wire [63:0] _341;
    wire [63:0] _5430;
    wire [63:0] _5436;
    wire [63:0] _9;
    reg [63:0] _312;
    wire _314;
    wire _315;
    wire _309;
    wire _316;
    wire _319;
    wire [63:0] _346;
    wire [63:0] _344;
    wire [63:0] _347;
    wire [63:0] _361;
    wire [63:0] _5437;
    wire [63:0] _5443;
    wire [63:0] _10;
    reg [63:0] _331;
    wire _333;
    wire _334;
    wire _328;
    wire _335;
    wire _338;
    wire [63:0] _366;
    wire [63:0] _364;
    wire [63:0] _367;
    wire [63:0] _381;
    wire [63:0] _5444;
    wire [63:0] _5450;
    wire [63:0] _11;
    reg [63:0] _351;
    wire _353;
    wire _354;
    wire _348;
    wire _355;
    wire _358;
    wire [63:0] _386;
    wire [63:0] _384;
    wire [63:0] _387;
    wire [63:0] _401;
    wire [63:0] _5451;
    wire [63:0] _5457;
    wire [63:0] _12;
    reg [63:0] _371;
    wire _373;
    wire _374;
    wire _368;
    wire _375;
    wire _378;
    wire [63:0] _406;
    wire [63:0] _404;
    wire [63:0] _407;
    wire [63:0] _421;
    wire [63:0] _5458;
    wire [63:0] _5464;
    wire [63:0] _13;
    reg [63:0] _391;
    wire _393;
    wire _394;
    wire _388;
    wire _395;
    wire _398;
    wire [63:0] _426;
    wire [63:0] _424;
    wire [63:0] _427;
    wire [63:0] _441;
    wire [63:0] _5465;
    wire [63:0] _5471;
    wire [63:0] _14;
    reg [63:0] _411;
    wire _413;
    wire _414;
    wire _408;
    wire _415;
    wire _418;
    wire [63:0] _446;
    wire [63:0] _444;
    wire [63:0] _447;
    wire [63:0] _461;
    wire [63:0] _5472;
    wire [63:0] _5478;
    wire [63:0] _15;
    reg [63:0] _431;
    wire _433;
    wire _434;
    wire _428;
    wire _435;
    wire _438;
    wire [63:0] _466;
    wire [63:0] _464;
    wire [63:0] _467;
    wire [63:0] _481;
    wire [63:0] _5479;
    wire [63:0] _5485;
    wire [63:0] _16;
    reg [63:0] _451;
    wire _453;
    wire _454;
    wire _448;
    wire _455;
    wire _458;
    wire [63:0] _486;
    wire [63:0] _484;
    wire [63:0] _487;
    wire [63:0] _501;
    wire [63:0] _5486;
    wire [63:0] _5492;
    wire [63:0] _17;
    reg [63:0] _471;
    wire _473;
    wire _474;
    wire _468;
    wire _475;
    wire _478;
    wire [63:0] _506;
    wire [63:0] _504;
    wire [63:0] _507;
    wire [63:0] _521;
    wire [63:0] _5493;
    wire [63:0] _5499;
    wire [63:0] _18;
    reg [63:0] _491;
    wire _493;
    wire _494;
    wire _488;
    wire _495;
    wire _498;
    wire [63:0] _526;
    wire [63:0] _524;
    wire [63:0] _527;
    wire [63:0] _541;
    wire [63:0] _5500;
    wire [63:0] _5506;
    wire [63:0] _19;
    reg [63:0] _511;
    wire _513;
    wire _514;
    wire _508;
    wire _515;
    wire _518;
    wire [63:0] _546;
    wire [63:0] _544;
    wire [63:0] _547;
    wire [63:0] _561;
    wire [63:0] _5507;
    wire [63:0] _5513;
    wire [63:0] _20;
    reg [63:0] _531;
    wire _533;
    wire _534;
    wire _528;
    wire _535;
    wire _538;
    wire [63:0] _566;
    wire [63:0] _564;
    wire [63:0] _567;
    wire [63:0] _581;
    wire [63:0] _5514;
    wire [63:0] _5520;
    wire [63:0] _21;
    reg [63:0] _551;
    wire _553;
    wire _554;
    wire _548;
    wire _555;
    wire _558;
    wire [63:0] _586;
    wire [63:0] _584;
    wire [63:0] _587;
    wire [63:0] _601;
    wire [63:0] _5521;
    wire [63:0] _5527;
    wire [63:0] _22;
    reg [63:0] _571;
    wire _573;
    wire _574;
    wire _568;
    wire _575;
    wire _578;
    wire [63:0] _606;
    wire [63:0] _604;
    wire [63:0] _607;
    wire [63:0] _621;
    wire [63:0] _5528;
    wire [63:0] _5534;
    wire [63:0] _23;
    reg [63:0] _591;
    wire _593;
    wire _594;
    wire _588;
    wire _595;
    wire _598;
    wire [63:0] _626;
    wire [63:0] _624;
    wire [63:0] _627;
    wire [63:0] _641;
    wire [63:0] _5535;
    wire [63:0] _5541;
    wire [63:0] _24;
    reg [63:0] _611;
    wire _613;
    wire _614;
    wire _608;
    wire _615;
    wire _618;
    wire [63:0] _646;
    wire [63:0] _644;
    wire [63:0] _647;
    wire [63:0] _661;
    wire [63:0] _5542;
    wire [63:0] _5548;
    wire [63:0] _25;
    reg [63:0] _631;
    wire _633;
    wire _634;
    wire _628;
    wire _635;
    wire _638;
    wire [63:0] _666;
    wire [63:0] _664;
    wire [63:0] _667;
    wire [63:0] _681;
    wire [63:0] _5549;
    wire [63:0] _5555;
    wire [63:0] _26;
    reg [63:0] _651;
    wire _653;
    wire _654;
    wire _648;
    wire _655;
    wire _658;
    wire [63:0] _686;
    wire [63:0] _684;
    wire [63:0] _687;
    wire [63:0] _701;
    wire [63:0] _5556;
    wire [63:0] _5562;
    wire [63:0] _27;
    reg [63:0] _671;
    wire _673;
    wire _674;
    wire _668;
    wire _675;
    wire _678;
    wire [63:0] _706;
    wire [63:0] _704;
    wire [63:0] _707;
    wire [63:0] _721;
    wire [63:0] _5563;
    wire [63:0] _5569;
    wire [63:0] _28;
    reg [63:0] _691;
    wire _693;
    wire _694;
    wire _688;
    wire _695;
    wire _698;
    wire [63:0] _726;
    wire [63:0] _724;
    wire [63:0] _727;
    wire [63:0] _741;
    wire [63:0] _5570;
    wire [63:0] _5576;
    wire [63:0] _29;
    reg [63:0] _711;
    wire _713;
    wire _714;
    wire _708;
    wire _715;
    wire _718;
    wire [63:0] _746;
    wire [63:0] _744;
    wire [63:0] _747;
    wire [63:0] _761;
    wire [63:0] _5577;
    wire [63:0] _5583;
    wire [63:0] _30;
    reg [63:0] _731;
    wire _733;
    wire _734;
    wire _728;
    wire _735;
    wire _738;
    wire [63:0] _766;
    wire [63:0] _764;
    wire [63:0] _767;
    wire [63:0] _781;
    wire [63:0] _5584;
    wire [63:0] _5590;
    wire [63:0] _31;
    reg [63:0] _751;
    wire _753;
    wire _754;
    wire _748;
    wire _755;
    wire _758;
    wire [63:0] _786;
    wire [63:0] _784;
    wire [63:0] _787;
    wire [63:0] _801;
    wire [63:0] _5591;
    wire [63:0] _5597;
    wire [63:0] _32;
    reg [63:0] _771;
    wire _773;
    wire _774;
    wire _768;
    wire _775;
    wire _778;
    wire [63:0] _806;
    wire [63:0] _804;
    wire [63:0] _807;
    wire [63:0] _821;
    wire [63:0] _5598;
    wire [63:0] _5604;
    wire [63:0] _33;
    reg [63:0] _791;
    wire _793;
    wire _794;
    wire _788;
    wire _795;
    wire _798;
    wire [63:0] _826;
    wire [63:0] _824;
    wire [63:0] _827;
    wire [63:0] _841;
    wire [63:0] _5605;
    wire [63:0] _5611;
    wire [63:0] _34;
    reg [63:0] _811;
    wire _813;
    wire _814;
    wire _808;
    wire _815;
    wire _818;
    wire [63:0] _846;
    wire [63:0] _844;
    wire [63:0] _847;
    wire [63:0] _861;
    wire [63:0] _5612;
    wire [63:0] _5618;
    wire [63:0] _35;
    reg [63:0] _831;
    wire _833;
    wire _834;
    wire _828;
    wire _835;
    wire _838;
    wire [63:0] _866;
    wire [63:0] _864;
    wire [63:0] _867;
    wire [63:0] _881;
    wire [63:0] _5619;
    wire [63:0] _5625;
    wire [63:0] _36;
    reg [63:0] _851;
    wire _853;
    wire _854;
    wire _848;
    wire _855;
    wire _858;
    wire [63:0] _886;
    wire [63:0] _884;
    wire [63:0] _887;
    wire [63:0] _901;
    wire [63:0] _5626;
    wire [63:0] _5632;
    wire [63:0] _37;
    reg [63:0] _871;
    wire _873;
    wire _874;
    wire _868;
    wire _875;
    wire _878;
    wire [63:0] _906;
    wire [63:0] _904;
    wire [63:0] _907;
    wire [63:0] _921;
    wire [63:0] _5633;
    wire [63:0] _5639;
    wire [63:0] _38;
    reg [63:0] _891;
    wire _893;
    wire _894;
    wire _888;
    wire _895;
    wire _898;
    wire [63:0] _926;
    wire [63:0] _924;
    wire [63:0] _927;
    wire [63:0] _941;
    wire [63:0] _5640;
    wire [63:0] _5646;
    wire [63:0] _39;
    reg [63:0] _911;
    wire _913;
    wire _914;
    wire _908;
    wire _915;
    wire _918;
    wire [63:0] _946;
    wire [63:0] _944;
    wire [63:0] _947;
    wire [63:0] _961;
    wire [63:0] _5647;
    wire [63:0] _5653;
    wire [63:0] _40;
    reg [63:0] _931;
    wire _933;
    wire _934;
    wire _928;
    wire _935;
    wire _938;
    wire [63:0] _966;
    wire [63:0] _964;
    wire [63:0] _967;
    wire [63:0] _981;
    wire [63:0] _5654;
    wire [63:0] _5660;
    wire [63:0] _41;
    reg [63:0] _951;
    wire _953;
    wire _954;
    wire _948;
    wire _955;
    wire _958;
    wire [63:0] _986;
    wire [63:0] _984;
    wire [63:0] _987;
    wire [63:0] _1001;
    wire [63:0] _5661;
    wire [63:0] _5667;
    wire [63:0] _42;
    reg [63:0] _971;
    wire _973;
    wire _974;
    wire _968;
    wire _975;
    wire _978;
    wire [63:0] _1006;
    wire [63:0] _1004;
    wire [63:0] _1007;
    wire [63:0] _1021;
    wire [63:0] _5668;
    wire [63:0] _5674;
    wire [63:0] _43;
    reg [63:0] _991;
    wire _993;
    wire _994;
    wire _988;
    wire _995;
    wire _998;
    wire [63:0] _1026;
    wire [63:0] _1024;
    wire [63:0] _1027;
    wire [63:0] _1041;
    wire [63:0] _5675;
    wire [63:0] _5681;
    wire [63:0] _44;
    reg [63:0] _1011;
    wire _1013;
    wire _1014;
    wire _1008;
    wire _1015;
    wire _1018;
    wire [63:0] _1046;
    wire [63:0] _1044;
    wire [63:0] _1047;
    wire [63:0] _1061;
    wire [63:0] _5682;
    wire [63:0] _5688;
    wire [63:0] _45;
    reg [63:0] _1031;
    wire _1033;
    wire _1034;
    wire _1028;
    wire _1035;
    wire _1038;
    wire [63:0] _1066;
    wire [63:0] _1064;
    wire [63:0] _1067;
    wire [63:0] _1081;
    wire [63:0] _5689;
    wire [63:0] _5695;
    wire [63:0] _46;
    reg [63:0] _1051;
    wire _1053;
    wire _1054;
    wire _1048;
    wire _1055;
    wire _1058;
    wire [63:0] _1086;
    wire [63:0] _1084;
    wire [63:0] _1087;
    wire [63:0] _1101;
    wire [63:0] _5696;
    wire [63:0] _5702;
    wire [63:0] _47;
    reg [63:0] _1071;
    wire _1073;
    wire _1074;
    wire _1068;
    wire _1075;
    wire _1078;
    wire [63:0] _1106;
    wire [63:0] _1104;
    wire [63:0] _1107;
    wire [63:0] _1121;
    wire [63:0] _5703;
    wire [63:0] _5709;
    wire [63:0] _48;
    reg [63:0] _1091;
    wire _1093;
    wire _1094;
    wire _1088;
    wire _1095;
    wire _1098;
    wire [63:0] _1126;
    wire [63:0] _1124;
    wire [63:0] _1127;
    wire [63:0] _1141;
    wire [63:0] _5710;
    wire [63:0] _5716;
    wire [63:0] _49;
    reg [63:0] _1111;
    wire _1113;
    wire _1114;
    wire _1108;
    wire _1115;
    wire _1118;
    wire [63:0] _1146;
    wire [63:0] _1144;
    wire [63:0] _1147;
    wire [63:0] _1161;
    wire [63:0] _5717;
    wire [63:0] _5723;
    wire [63:0] _50;
    reg [63:0] _1131;
    wire _1133;
    wire _1134;
    wire _1128;
    wire _1135;
    wire _1138;
    wire [63:0] _1166;
    wire [63:0] _1164;
    wire [63:0] _1167;
    wire [63:0] _1181;
    wire [63:0] _5724;
    wire [63:0] _5730;
    wire [63:0] _51;
    reg [63:0] _1151;
    wire _1153;
    wire _1154;
    wire _1148;
    wire _1155;
    wire _1158;
    wire [63:0] _1186;
    wire [63:0] _1184;
    wire [63:0] _1187;
    wire [63:0] _1201;
    wire [63:0] _5731;
    wire [63:0] _5737;
    wire [63:0] _52;
    reg [63:0] _1171;
    wire _1173;
    wire _1174;
    wire _1168;
    wire _1175;
    wire _1178;
    wire [63:0] _1206;
    wire [63:0] _1204;
    wire [63:0] _1207;
    wire [63:0] _1221;
    wire [63:0] _5738;
    wire [63:0] _5744;
    wire [63:0] _53;
    reg [63:0] _1191;
    wire _1193;
    wire _1194;
    wire _1188;
    wire _1195;
    wire _1198;
    wire [63:0] _1226;
    wire [63:0] _1224;
    wire [63:0] _1227;
    wire [63:0] _1241;
    wire [63:0] _5745;
    wire [63:0] _5751;
    wire [63:0] _54;
    reg [63:0] _1211;
    wire _1213;
    wire _1214;
    wire _1208;
    wire _1215;
    wire _1218;
    wire [63:0] _1246;
    wire [63:0] _1244;
    wire [63:0] _1247;
    wire [63:0] _1261;
    wire [63:0] _5752;
    wire [63:0] _5758;
    wire [63:0] _55;
    reg [63:0] _1231;
    wire _1233;
    wire _1234;
    wire _1228;
    wire _1235;
    wire _1238;
    wire [63:0] _1266;
    wire [63:0] _1264;
    wire [63:0] _1267;
    wire [63:0] _1281;
    wire [63:0] _5759;
    wire [63:0] _5765;
    wire [63:0] _56;
    reg [63:0] _1251;
    wire _1253;
    wire _1254;
    wire _1248;
    wire _1255;
    wire _1258;
    wire [63:0] _1286;
    wire [63:0] _1284;
    wire [63:0] _1287;
    wire [63:0] _1301;
    wire [63:0] _5766;
    wire [63:0] _5772;
    wire [63:0] _57;
    reg [63:0] _1271;
    wire _1273;
    wire _1274;
    wire _1268;
    wire _1275;
    wire _1278;
    wire [63:0] _1306;
    wire [63:0] _1304;
    wire [63:0] _1307;
    wire [63:0] _1321;
    wire [63:0] _5773;
    wire [63:0] _5779;
    wire [63:0] _58;
    reg [63:0] _1291;
    wire _1293;
    wire _1294;
    wire _1288;
    wire _1295;
    wire _1298;
    wire [63:0] _1326;
    wire [63:0] _1324;
    wire [63:0] _1327;
    wire [63:0] _1341;
    wire [63:0] _5780;
    wire [63:0] _5786;
    wire [63:0] _59;
    reg [63:0] _1311;
    wire _1313;
    wire _1314;
    wire _1308;
    wire _1315;
    wire _1318;
    wire [63:0] _1346;
    wire [63:0] _1344;
    wire [63:0] _1347;
    wire [63:0] _1361;
    wire [63:0] _5787;
    wire [63:0] _5793;
    wire [63:0] _60;
    reg [63:0] _1331;
    wire _1333;
    wire _1334;
    wire _1328;
    wire _1335;
    wire _1338;
    wire [63:0] _1366;
    wire [63:0] _1364;
    wire [63:0] _1367;
    wire [63:0] _1381;
    wire [63:0] _5794;
    wire [63:0] _5800;
    wire [63:0] _61;
    reg [63:0] _1351;
    wire _1353;
    wire _1354;
    wire _1348;
    wire _1355;
    wire _1358;
    wire [63:0] _1386;
    wire [63:0] _1384;
    wire [63:0] _1387;
    wire [63:0] _1401;
    wire [63:0] _5801;
    wire [63:0] _5807;
    wire [63:0] _62;
    reg [63:0] _1371;
    wire _1373;
    wire _1374;
    wire _1368;
    wire _1375;
    wire _1378;
    wire [63:0] _1406;
    wire [63:0] _1404;
    wire [63:0] _1407;
    wire [63:0] _1421;
    wire [63:0] _5808;
    wire [63:0] _5814;
    wire [63:0] _63;
    reg [63:0] _1391;
    wire _1393;
    wire _1394;
    wire _1388;
    wire _1395;
    wire _1398;
    wire [63:0] _1426;
    wire [63:0] _1424;
    wire [63:0] _1427;
    wire [63:0] _1441;
    wire [63:0] _5815;
    wire [63:0] _5821;
    wire [63:0] _64;
    reg [63:0] _1411;
    wire _1413;
    wire _1414;
    wire _1408;
    wire _1415;
    wire _1418;
    wire [63:0] _1446;
    wire [63:0] _1444;
    wire [63:0] _1447;
    wire [63:0] _1461;
    wire [63:0] _5822;
    wire [63:0] _5828;
    wire [63:0] _65;
    reg [63:0] _1431;
    wire _1433;
    wire _1434;
    wire _1428;
    wire _1435;
    wire _1438;
    wire [63:0] _1466;
    wire [63:0] _1464;
    wire [63:0] _1467;
    wire [63:0] _1481;
    wire [63:0] _5829;
    wire [63:0] _5835;
    wire [63:0] _66;
    reg [63:0] _1451;
    wire _1453;
    wire _1454;
    wire _1448;
    wire _1455;
    wire _1458;
    wire [63:0] _1486;
    wire [63:0] _1484;
    wire [63:0] _1487;
    wire [63:0] _1501;
    wire [63:0] _5836;
    wire [63:0] _5842;
    wire [63:0] _67;
    reg [63:0] _1471;
    wire _1473;
    wire _1474;
    wire _1468;
    wire _1475;
    wire _1478;
    wire [63:0] _1506;
    wire [63:0] _1504;
    wire [63:0] _1507;
    wire [63:0] _1521;
    wire [63:0] _5843;
    wire [63:0] _5849;
    wire [63:0] _68;
    reg [63:0] _1491;
    wire _1493;
    wire _1494;
    wire _1488;
    wire _1495;
    wire _1498;
    wire [63:0] _1526;
    wire [63:0] _1524;
    wire [63:0] _1527;
    wire [63:0] _1541;
    wire [63:0] _5850;
    wire [63:0] _5856;
    wire [63:0] _69;
    reg [63:0] _1511;
    wire _1513;
    wire _1514;
    wire _1508;
    wire _1515;
    wire _1518;
    wire [63:0] _1546;
    wire [63:0] _1544;
    wire [63:0] _1547;
    wire [63:0] _1561;
    wire [63:0] _5857;
    wire [63:0] _5863;
    wire [63:0] _70;
    reg [63:0] _1531;
    wire _1533;
    wire _1534;
    wire _1528;
    wire _1535;
    wire _1538;
    wire [63:0] _1566;
    wire [63:0] _1564;
    wire [63:0] _1567;
    wire [63:0] _1581;
    wire [63:0] _5864;
    wire [63:0] _5870;
    wire [63:0] _71;
    reg [63:0] _1551;
    wire _1553;
    wire _1554;
    wire _1548;
    wire _1555;
    wire _1558;
    wire [63:0] _1586;
    wire [63:0] _1584;
    wire [63:0] _1587;
    wire [63:0] _1601;
    wire [63:0] _5871;
    wire [63:0] _5877;
    wire [63:0] _72;
    reg [63:0] _1571;
    wire _1573;
    wire _1574;
    wire _1568;
    wire _1575;
    wire _1578;
    wire [63:0] _1606;
    wire [63:0] _1604;
    wire [63:0] _1607;
    wire [63:0] _1621;
    wire [63:0] _5878;
    wire [63:0] _5884;
    wire [63:0] _73;
    reg [63:0] _1591;
    wire _1593;
    wire _1594;
    wire _1588;
    wire _1595;
    wire _1598;
    wire [63:0] _1626;
    wire [63:0] _1624;
    wire [63:0] _1627;
    wire [63:0] _1641;
    wire [63:0] _5885;
    wire [63:0] _5891;
    wire [63:0] _74;
    reg [63:0] _1611;
    wire _1613;
    wire _1614;
    wire _1608;
    wire _1615;
    wire _1618;
    wire [63:0] _1646;
    wire [63:0] _1644;
    wire [63:0] _1647;
    wire [63:0] _1661;
    wire [63:0] _5892;
    wire [63:0] _5898;
    wire [63:0] _75;
    reg [63:0] _1631;
    wire _1633;
    wire _1634;
    wire _1628;
    wire _1635;
    wire _1638;
    wire [63:0] _1666;
    wire [63:0] _1664;
    wire [63:0] _1667;
    wire [63:0] _1681;
    wire [63:0] _5899;
    wire [63:0] _5905;
    wire [63:0] _76;
    reg [63:0] _1651;
    wire _1653;
    wire _1654;
    wire _1648;
    wire _1655;
    wire _1658;
    wire [63:0] _1686;
    wire [63:0] _1684;
    wire [63:0] _1687;
    wire [63:0] _1701;
    wire [63:0] _5906;
    wire [63:0] _5912;
    wire [63:0] _77;
    reg [63:0] _1671;
    wire _1673;
    wire _1674;
    wire _1668;
    wire _1675;
    wire _1678;
    wire [63:0] _1706;
    wire [63:0] _1704;
    wire [63:0] _1707;
    wire [63:0] _1721;
    wire [63:0] _5913;
    wire [63:0] _5919;
    wire [63:0] _78;
    reg [63:0] _1691;
    wire _1693;
    wire _1694;
    wire _1688;
    wire _1695;
    wire _1698;
    wire [63:0] _1726;
    wire [63:0] _1724;
    wire [63:0] _1727;
    wire [63:0] _1741;
    wire [63:0] _5920;
    wire [63:0] _5926;
    wire [63:0] _79;
    reg [63:0] _1711;
    wire _1713;
    wire _1714;
    wire _1708;
    wire _1715;
    wire _1718;
    wire [63:0] _1746;
    wire [63:0] _1744;
    wire [63:0] _1747;
    wire [63:0] _1761;
    wire [63:0] _5927;
    wire [63:0] _5933;
    wire [63:0] _80;
    reg [63:0] _1731;
    wire _1733;
    wire _1734;
    wire _1728;
    wire _1735;
    wire _1738;
    wire [63:0] _1766;
    wire [63:0] _1764;
    wire [63:0] _1767;
    wire [63:0] _1781;
    wire [63:0] _5934;
    wire [63:0] _5940;
    wire [63:0] _81;
    reg [63:0] _1751;
    wire _1753;
    wire _1754;
    wire _1748;
    wire _1755;
    wire _1758;
    wire [63:0] _1786;
    wire [63:0] _1784;
    wire [63:0] _1787;
    wire [63:0] _1801;
    wire [63:0] _5941;
    wire [63:0] _5947;
    wire [63:0] _82;
    reg [63:0] _1771;
    wire _1773;
    wire _1774;
    wire _1768;
    wire _1775;
    wire _1778;
    wire [63:0] _1806;
    wire [63:0] _1804;
    wire [63:0] _1807;
    wire [63:0] _1821;
    wire [63:0] _5948;
    wire [63:0] _5954;
    wire [63:0] _83;
    reg [63:0] _1791;
    wire _1793;
    wire _1794;
    wire _1788;
    wire _1795;
    wire _1798;
    wire [63:0] _1826;
    wire [63:0] _1824;
    wire [63:0] _1827;
    wire [63:0] _1841;
    wire [63:0] _5955;
    wire [63:0] _5961;
    wire [63:0] _84;
    reg [63:0] _1811;
    wire _1813;
    wire _1814;
    wire _1808;
    wire _1815;
    wire _1818;
    wire [63:0] _1846;
    wire [63:0] _1844;
    wire [63:0] _1847;
    wire [63:0] _1861;
    wire [63:0] _5962;
    wire [63:0] _5968;
    wire [63:0] _85;
    reg [63:0] _1831;
    wire _1833;
    wire _1834;
    wire _1828;
    wire _1835;
    wire _1838;
    wire [63:0] _1866;
    wire [63:0] _1864;
    wire [63:0] _1867;
    wire [63:0] _1881;
    wire [63:0] _5969;
    wire [63:0] _5975;
    wire [63:0] _86;
    reg [63:0] _1851;
    wire _1853;
    wire _1854;
    wire _1848;
    wire _1855;
    wire _1858;
    wire [63:0] _1886;
    wire [63:0] _1884;
    wire [63:0] _1887;
    wire [63:0] _1901;
    wire [63:0] _5976;
    wire [63:0] _5982;
    wire [63:0] _87;
    reg [63:0] _1871;
    wire _1873;
    wire _1874;
    wire _1868;
    wire _1875;
    wire _1878;
    wire [63:0] _1906;
    wire [63:0] _1904;
    wire [63:0] _1907;
    wire [63:0] _1921;
    wire [63:0] _5983;
    wire [63:0] _5989;
    wire [63:0] _88;
    reg [63:0] _1891;
    wire _1893;
    wire _1894;
    wire _1888;
    wire _1895;
    wire _1898;
    wire [63:0] _1926;
    wire [63:0] _1924;
    wire [63:0] _1927;
    wire [63:0] _1941;
    wire [63:0] _5990;
    wire [63:0] _5996;
    wire [63:0] _89;
    reg [63:0] _1911;
    wire _1913;
    wire _1914;
    wire _1908;
    wire _1915;
    wire _1918;
    wire [63:0] _1946;
    wire [63:0] _1944;
    wire [63:0] _1947;
    wire [63:0] _1961;
    wire [63:0] _5997;
    wire [63:0] _6003;
    wire [63:0] _90;
    reg [63:0] _1931;
    wire _1933;
    wire _1934;
    wire _1928;
    wire _1935;
    wire _1938;
    wire [63:0] _1966;
    wire [63:0] _1964;
    wire [63:0] _1967;
    wire [63:0] _1981;
    wire [63:0] _6004;
    wire [63:0] _6010;
    wire [63:0] _91;
    reg [63:0] _1951;
    wire _1953;
    wire _1954;
    wire _1948;
    wire _1955;
    wire _1958;
    wire [63:0] _1986;
    wire [63:0] _1984;
    wire [63:0] _1987;
    wire [63:0] _2001;
    wire [63:0] _6011;
    wire [63:0] _6017;
    wire [63:0] _92;
    reg [63:0] _1971;
    wire _1973;
    wire _1974;
    wire _1968;
    wire _1975;
    wire _1978;
    wire [63:0] _2006;
    wire [63:0] _2004;
    wire [63:0] _2007;
    wire [63:0] _2021;
    wire [63:0] _6018;
    wire [63:0] _6024;
    wire [63:0] _93;
    reg [63:0] _1991;
    wire _1993;
    wire _1994;
    wire _1988;
    wire _1995;
    wire _1998;
    wire [63:0] _2026;
    wire [63:0] _2024;
    wire [63:0] _2027;
    wire [63:0] _2041;
    wire [63:0] _6025;
    wire [63:0] _6031;
    wire [63:0] _94;
    reg [63:0] _2011;
    wire _2013;
    wire _2014;
    wire _2008;
    wire _2015;
    wire _2018;
    wire [63:0] _2046;
    wire [63:0] _2044;
    wire [63:0] _2047;
    wire [63:0] _2061;
    wire [63:0] _6032;
    wire [63:0] _6038;
    wire [63:0] _95;
    reg [63:0] _2031;
    wire _2033;
    wire _2034;
    wire _2028;
    wire _2035;
    wire _2038;
    wire [63:0] _2066;
    wire [63:0] _2064;
    wire [63:0] _2067;
    wire [63:0] _2081;
    wire [63:0] _6039;
    wire [63:0] _6045;
    wire [63:0] _96;
    reg [63:0] _2051;
    wire _2053;
    wire _2054;
    wire _2048;
    wire _2055;
    wire _2058;
    wire [63:0] _2086;
    wire [63:0] _2084;
    wire [63:0] _2087;
    wire [63:0] _2101;
    wire [63:0] _6046;
    wire [63:0] _6052;
    wire [63:0] _97;
    reg [63:0] _2071;
    wire _2073;
    wire _2074;
    wire _2068;
    wire _2075;
    wire _2078;
    wire [63:0] _2106;
    wire [63:0] _2104;
    wire [63:0] _2107;
    wire [63:0] _2121;
    wire [63:0] _6053;
    wire [63:0] _6059;
    wire [63:0] _98;
    reg [63:0] _2091;
    wire _2093;
    wire _2094;
    wire _2088;
    wire _2095;
    wire _2098;
    wire [63:0] _2126;
    wire [63:0] _2124;
    wire [63:0] _2127;
    wire [63:0] _2141;
    wire [63:0] _6060;
    wire [63:0] _6066;
    wire [63:0] _99;
    reg [63:0] _2111;
    wire _2113;
    wire _2114;
    wire _2108;
    wire _2115;
    wire _2118;
    wire [63:0] _2146;
    wire [63:0] _2144;
    wire [63:0] _2147;
    wire [63:0] _2161;
    wire [63:0] _6067;
    wire [63:0] _6073;
    wire [63:0] _100;
    reg [63:0] _2131;
    wire _2133;
    wire _2134;
    wire _2128;
    wire _2135;
    wire _2138;
    wire [63:0] _2166;
    wire [63:0] _2164;
    wire [63:0] _2167;
    wire [63:0] _2181;
    wire [63:0] _6074;
    wire [63:0] _6080;
    wire [63:0] _101;
    reg [63:0] _2151;
    wire _2153;
    wire _2154;
    wire _2148;
    wire _2155;
    wire _2158;
    wire [63:0] _2186;
    wire [63:0] _2184;
    wire [63:0] _2187;
    wire [63:0] _2201;
    wire [63:0] _6081;
    wire [63:0] _6087;
    wire [63:0] _102;
    reg [63:0] _2171;
    wire _2173;
    wire _2174;
    wire _2168;
    wire _2175;
    wire _2178;
    wire [63:0] _2206;
    wire [63:0] _2204;
    wire [63:0] _2207;
    wire [63:0] _2221;
    wire [63:0] _6088;
    wire [63:0] _6094;
    wire [63:0] _103;
    reg [63:0] _2191;
    wire _2193;
    wire _2194;
    wire _2188;
    wire _2195;
    wire _2198;
    wire [63:0] _2226;
    wire [63:0] _2224;
    wire [63:0] _2227;
    wire [63:0] _2241;
    wire [63:0] _6095;
    wire [63:0] _6101;
    wire [63:0] _104;
    reg [63:0] _2211;
    wire _2213;
    wire _2214;
    wire _2208;
    wire _2215;
    wire _2218;
    wire [63:0] _2246;
    wire [63:0] _2244;
    wire [63:0] _2247;
    wire [63:0] _2261;
    wire [63:0] _6102;
    wire [63:0] _6108;
    wire [63:0] _105;
    reg [63:0] _2231;
    wire _2233;
    wire _2234;
    wire _2228;
    wire _2235;
    wire _2238;
    wire [63:0] _2266;
    wire [63:0] _2264;
    wire [63:0] _2267;
    wire [63:0] _2281;
    wire [63:0] _6109;
    wire [63:0] _6115;
    wire [63:0] _106;
    reg [63:0] _2251;
    wire _2253;
    wire _2254;
    wire _2248;
    wire _2255;
    wire _2258;
    wire [63:0] _2286;
    wire [63:0] _2284;
    wire [63:0] _2287;
    wire [63:0] _2301;
    wire [63:0] _6116;
    wire [63:0] _6122;
    wire [63:0] _107;
    reg [63:0] _2271;
    wire _2273;
    wire _2274;
    wire _2268;
    wire _2275;
    wire _2278;
    wire [63:0] _2306;
    wire [63:0] _2304;
    wire [63:0] _2307;
    wire [63:0] _2321;
    wire [63:0] _6123;
    wire [63:0] _6129;
    wire [63:0] _108;
    reg [63:0] _2291;
    wire _2293;
    wire _2294;
    wire _2288;
    wire _2295;
    wire _2298;
    wire [63:0] _2326;
    wire [63:0] _2324;
    wire [63:0] _2327;
    wire [63:0] _2341;
    wire [63:0] _6130;
    wire [63:0] _6136;
    wire [63:0] _109;
    reg [63:0] _2311;
    wire _2313;
    wire _2314;
    wire _2308;
    wire _2315;
    wire _2318;
    wire [63:0] _2346;
    wire [63:0] _2344;
    wire [63:0] _2347;
    wire [63:0] _2361;
    wire [63:0] _6137;
    wire [63:0] _6143;
    wire [63:0] _110;
    reg [63:0] _2331;
    wire _2333;
    wire _2334;
    wire _2328;
    wire _2335;
    wire _2338;
    wire [63:0] _2366;
    wire [63:0] _2364;
    wire [63:0] _2367;
    wire [63:0] _2381;
    wire [63:0] _6144;
    wire [63:0] _6150;
    wire [63:0] _111;
    reg [63:0] _2351;
    wire _2353;
    wire _2354;
    wire _2348;
    wire _2355;
    wire _2358;
    wire [63:0] _2386;
    wire [63:0] _2384;
    wire [63:0] _2387;
    wire [63:0] _2401;
    wire [63:0] _6151;
    wire [63:0] _6157;
    wire [63:0] _112;
    reg [63:0] _2371;
    wire _2373;
    wire _2374;
    wire _2368;
    wire _2375;
    wire _2378;
    wire [63:0] _2406;
    wire [63:0] _2404;
    wire [63:0] _2407;
    wire [63:0] _2421;
    wire [63:0] _6158;
    wire [63:0] _6164;
    wire [63:0] _113;
    reg [63:0] _2391;
    wire _2393;
    wire _2394;
    wire _2388;
    wire _2395;
    wire _2398;
    wire [63:0] _2426;
    wire [63:0] _2424;
    wire [63:0] _2427;
    wire [63:0] _2441;
    wire [63:0] _6165;
    wire [63:0] _6171;
    wire [63:0] _114;
    reg [63:0] _2411;
    wire _2413;
    wire _2414;
    wire _2408;
    wire _2415;
    wire _2418;
    wire [63:0] _2446;
    wire [63:0] _2444;
    wire [63:0] _2447;
    wire [63:0] _2461;
    wire [63:0] _6172;
    wire [63:0] _6178;
    wire [63:0] _115;
    reg [63:0] _2431;
    wire _2433;
    wire _2434;
    wire _2428;
    wire _2435;
    wire _2438;
    wire [63:0] _2466;
    wire [63:0] _2464;
    wire [63:0] _2467;
    wire [63:0] _2481;
    wire [63:0] _6179;
    wire [63:0] _6185;
    wire [63:0] _116;
    reg [63:0] _2451;
    wire _2453;
    wire _2454;
    wire _2448;
    wire _2455;
    wire _2458;
    wire [63:0] _2486;
    wire [63:0] _2484;
    wire [63:0] _2487;
    wire [63:0] _2501;
    wire [63:0] _6186;
    wire [63:0] _6192;
    wire [63:0] _117;
    reg [63:0] _2471;
    wire _2473;
    wire _2474;
    wire _2468;
    wire _2475;
    wire _2478;
    wire [63:0] _2506;
    wire [63:0] _2504;
    wire [63:0] _2507;
    wire [63:0] _2521;
    wire [63:0] _6193;
    wire [63:0] _6199;
    wire [63:0] _118;
    reg [63:0] _2491;
    wire _2493;
    wire _2494;
    wire _2488;
    wire _2495;
    wire _2498;
    wire [63:0] _2526;
    wire [63:0] _2524;
    wire [63:0] _2527;
    wire [63:0] _2541;
    wire [63:0] _6200;
    wire [63:0] _6206;
    wire [63:0] _119;
    reg [63:0] _2511;
    wire _2513;
    wire _2514;
    wire _2508;
    wire _2515;
    wire _2518;
    wire [63:0] _2546;
    wire [63:0] _2544;
    wire [63:0] _2547;
    wire [63:0] _2561;
    wire [63:0] _6207;
    wire [63:0] _6213;
    wire [63:0] _120;
    reg [63:0] _2531;
    wire _2533;
    wire _2534;
    wire _2528;
    wire _2535;
    wire _2538;
    wire [63:0] _2566;
    wire [63:0] _2564;
    wire [63:0] _2567;
    wire [63:0] _2581;
    wire [63:0] _6214;
    wire [63:0] _6220;
    wire [63:0] _121;
    reg [63:0] _2551;
    wire _2553;
    wire _2554;
    wire _2548;
    wire _2555;
    wire _2558;
    wire [63:0] _2586;
    wire [63:0] _2584;
    wire [63:0] _2587;
    wire [63:0] _2601;
    wire [63:0] _6221;
    wire [63:0] _6227;
    wire [63:0] _122;
    reg [63:0] _2571;
    wire _2573;
    wire _2574;
    wire _2568;
    wire _2575;
    wire _2578;
    wire [63:0] _2606;
    wire [63:0] _2604;
    wire [63:0] _2607;
    wire [63:0] _2621;
    wire [63:0] _6228;
    wire [63:0] _6234;
    wire [63:0] _123;
    reg [63:0] _2591;
    wire _2593;
    wire _2594;
    wire _2588;
    wire _2595;
    wire _2598;
    wire [63:0] _2626;
    wire [63:0] _2624;
    wire [63:0] _2627;
    wire [63:0] _2641;
    wire [63:0] _6235;
    wire [63:0] _6241;
    wire [63:0] _124;
    reg [63:0] _2611;
    wire _2613;
    wire _2614;
    wire _2608;
    wire _2615;
    wire _2618;
    wire [63:0] _2646;
    wire [63:0] _2644;
    wire [63:0] _2647;
    wire [63:0] _2661;
    wire [63:0] _6242;
    wire [63:0] _6248;
    wire [63:0] _125;
    reg [63:0] _2631;
    wire _2633;
    wire _2634;
    wire _2628;
    wire _2635;
    wire _2638;
    wire [63:0] _2666;
    wire [63:0] _2664;
    wire [63:0] _2667;
    wire [63:0] _2681;
    wire [63:0] _6249;
    wire [63:0] _6255;
    wire [63:0] _126;
    reg [63:0] _2651;
    wire _2653;
    wire _2654;
    wire _2648;
    wire _2655;
    wire _2658;
    wire [63:0] _2686;
    wire [63:0] _2684;
    wire [63:0] _2687;
    wire [63:0] _2701;
    wire [63:0] _6256;
    wire [63:0] _6262;
    wire [63:0] _127;
    reg [63:0] _2671;
    wire _2673;
    wire _2674;
    wire _2668;
    wire _2675;
    wire _2678;
    wire [63:0] _2706;
    wire [63:0] _2704;
    wire [63:0] _2707;
    wire [63:0] _2721;
    wire [63:0] _6263;
    wire [63:0] _6269;
    wire [63:0] _128;
    reg [63:0] _2691;
    wire _2693;
    wire _2694;
    wire _2688;
    wire _2695;
    wire _2698;
    wire [63:0] _2726;
    wire [63:0] _2724;
    wire [63:0] _2727;
    wire [63:0] _2741;
    wire [63:0] _6270;
    wire [63:0] _6276;
    wire [63:0] _129;
    reg [63:0] _2711;
    wire _2713;
    wire _2714;
    wire _2708;
    wire _2715;
    wire _2718;
    wire [63:0] _2746;
    wire [63:0] _2744;
    wire [63:0] _2747;
    wire [63:0] _2761;
    wire [63:0] _6277;
    wire [63:0] _6283;
    wire [63:0] _130;
    reg [63:0] _2731;
    wire _2733;
    wire _2734;
    wire _2728;
    wire _2735;
    wire _2738;
    wire [63:0] _2766;
    wire [63:0] _2764;
    wire [63:0] _2767;
    wire [63:0] _2781;
    wire [63:0] _6284;
    wire [63:0] _6290;
    wire [63:0] _131;
    reg [63:0] _2751;
    wire _2753;
    wire _2754;
    wire _2748;
    wire _2755;
    wire _2758;
    wire [63:0] _2786;
    wire [63:0] _2784;
    wire [63:0] _2787;
    wire [63:0] _2801;
    wire [63:0] _6291;
    wire [63:0] _6297;
    wire [63:0] _132;
    reg [63:0] _2771;
    wire _2773;
    wire _2774;
    wire _2768;
    wire _2775;
    wire _2778;
    wire [63:0] _2806;
    wire [63:0] _2804;
    wire [63:0] _2807;
    wire [63:0] _2821;
    wire [63:0] _6298;
    wire [63:0] _6304;
    wire [63:0] _133;
    reg [63:0] _2791;
    wire _2793;
    wire _2794;
    wire _2788;
    wire _2795;
    wire _2798;
    wire [63:0] _2826;
    wire [63:0] _2824;
    wire [63:0] _2827;
    wire [63:0] _2841;
    wire [63:0] _6305;
    wire [63:0] _6311;
    wire [63:0] _134;
    reg [63:0] _2811;
    wire _2813;
    wire _2814;
    wire _2808;
    wire _2815;
    wire _2818;
    wire [63:0] _2846;
    wire [63:0] _2844;
    wire [63:0] _2847;
    wire [63:0] _2861;
    wire [63:0] _6312;
    wire [63:0] _6318;
    wire [63:0] _135;
    reg [63:0] _2831;
    wire _2833;
    wire _2834;
    wire _2828;
    wire _2835;
    wire _2838;
    wire [63:0] _2866;
    wire [63:0] _2864;
    wire [63:0] _2867;
    wire [63:0] _2881;
    wire [63:0] _6319;
    wire [63:0] _6325;
    wire [63:0] _136;
    reg [63:0] _2851;
    wire _2853;
    wire _2854;
    wire _2848;
    wire _2855;
    wire _2858;
    wire [63:0] _2886;
    wire [63:0] _2884;
    wire [63:0] _2887;
    wire [63:0] _2901;
    wire [63:0] _6326;
    wire [63:0] _6332;
    wire [63:0] _137;
    reg [63:0] _2871;
    wire _2873;
    wire _2874;
    wire _2868;
    wire _2875;
    wire _2878;
    wire [63:0] _2906;
    wire [63:0] _2904;
    wire [63:0] _2907;
    wire [63:0] _2921;
    wire [63:0] _6333;
    wire [63:0] _6339;
    wire [63:0] _138;
    reg [63:0] _2891;
    wire _2893;
    wire _2894;
    wire _2888;
    wire _2895;
    wire _2898;
    wire [63:0] _2926;
    wire [63:0] _2924;
    wire [63:0] _2927;
    wire [63:0] _2941;
    wire [63:0] _6340;
    wire [63:0] _6346;
    wire [63:0] _139;
    reg [63:0] _2911;
    wire _2913;
    wire _2914;
    wire _2908;
    wire _2915;
    wire _2918;
    wire [63:0] _2946;
    wire [63:0] _2944;
    wire [63:0] _2947;
    wire [63:0] _2961;
    wire [63:0] _6347;
    wire [63:0] _6353;
    wire [63:0] _140;
    reg [63:0] _2931;
    wire _2933;
    wire _2934;
    wire _2928;
    wire _2935;
    wire _2938;
    wire [63:0] _2966;
    wire [63:0] _2964;
    wire [63:0] _2967;
    wire [63:0] _2981;
    wire [63:0] _6354;
    wire [63:0] _6360;
    wire [63:0] _141;
    reg [63:0] _2951;
    wire _2953;
    wire _2954;
    wire _2948;
    wire _2955;
    wire _2958;
    wire [63:0] _2986;
    wire [63:0] _2984;
    wire [63:0] _2987;
    wire [63:0] _3001;
    wire [63:0] _6361;
    wire [63:0] _6367;
    wire [63:0] _142;
    reg [63:0] _2971;
    wire _2973;
    wire _2974;
    wire _2968;
    wire _2975;
    wire _2978;
    wire [63:0] _3006;
    wire [63:0] _3004;
    wire [63:0] _3007;
    wire [63:0] _3021;
    wire [63:0] _6368;
    wire [63:0] _6374;
    wire [63:0] _143;
    reg [63:0] _2991;
    wire _2993;
    wire _2994;
    wire _2988;
    wire _2995;
    wire _2998;
    wire [63:0] _3026;
    wire [63:0] _3024;
    wire [63:0] _3027;
    wire [63:0] _3041;
    wire [63:0] _6375;
    wire [63:0] _6381;
    wire [63:0] _144;
    reg [63:0] _3011;
    wire _3013;
    wire _3014;
    wire _3008;
    wire _3015;
    wire _3018;
    wire [63:0] _3046;
    wire [63:0] _3044;
    wire [63:0] _3047;
    wire [63:0] _3061;
    wire [63:0] _6382;
    wire [63:0] _6388;
    wire [63:0] _145;
    reg [63:0] _3031;
    wire _3033;
    wire _3034;
    wire _3028;
    wire _3035;
    wire _3038;
    wire [63:0] _3066;
    wire [63:0] _3064;
    wire [63:0] _3067;
    wire [63:0] _3081;
    wire [63:0] _6389;
    wire [63:0] _6395;
    wire [63:0] _146;
    reg [63:0] _3051;
    wire _3053;
    wire _3054;
    wire _3048;
    wire _3055;
    wire _3058;
    wire [63:0] _3086;
    wire [63:0] _3084;
    wire [63:0] _3087;
    wire [63:0] _3101;
    wire [63:0] _6396;
    wire [63:0] _6402;
    wire [63:0] _147;
    reg [63:0] _3071;
    wire _3073;
    wire _3074;
    wire _3068;
    wire _3075;
    wire _3078;
    wire [63:0] _3106;
    wire [63:0] _3104;
    wire [63:0] _3107;
    wire [63:0] _3121;
    wire [63:0] _6403;
    wire [63:0] _6409;
    wire [63:0] _148;
    reg [63:0] _3091;
    wire _3093;
    wire _3094;
    wire _3088;
    wire _3095;
    wire _3098;
    wire [63:0] _3126;
    wire [63:0] _3124;
    wire [63:0] _3127;
    wire [63:0] _3141;
    wire [63:0] _6410;
    wire [63:0] _6416;
    wire [63:0] _149;
    reg [63:0] _3111;
    wire _3113;
    wire _3114;
    wire _3108;
    wire _3115;
    wire _3118;
    wire [63:0] _3146;
    wire [63:0] _3144;
    wire [63:0] _3147;
    wire [63:0] _3161;
    wire [63:0] _6417;
    wire [63:0] _6423;
    wire [63:0] _150;
    reg [63:0] _3131;
    wire _3133;
    wire _3134;
    wire _3128;
    wire _3135;
    wire _3138;
    wire [63:0] _3166;
    wire [63:0] _3164;
    wire [63:0] _3167;
    wire [63:0] _3181;
    wire [63:0] _6424;
    wire [63:0] _6430;
    wire [63:0] _151;
    reg [63:0] _3151;
    wire _3153;
    wire _3154;
    wire _3148;
    wire _3155;
    wire _3158;
    wire [63:0] _3186;
    wire [63:0] _3184;
    wire [63:0] _3187;
    wire [63:0] _3201;
    wire [63:0] _6431;
    wire [63:0] _6437;
    wire [63:0] _152;
    reg [63:0] _3171;
    wire _3173;
    wire _3174;
    wire _3168;
    wire _3175;
    wire _3178;
    wire [63:0] _3206;
    wire [63:0] _3204;
    wire [63:0] _3207;
    wire [63:0] _3221;
    wire [63:0] _6438;
    wire [63:0] _6444;
    wire [63:0] _153;
    reg [63:0] _3191;
    wire _3193;
    wire _3194;
    wire _3188;
    wire _3195;
    wire _3198;
    wire [63:0] _3226;
    wire [63:0] _3224;
    wire [63:0] _3227;
    wire [63:0] _3241;
    wire [63:0] _6445;
    wire [63:0] _6451;
    wire [63:0] _154;
    reg [63:0] _3211;
    wire _3213;
    wire _3214;
    wire _3208;
    wire _3215;
    wire _3218;
    wire [63:0] _3246;
    wire [63:0] _3244;
    wire [63:0] _3247;
    wire [63:0] _3261;
    wire [63:0] _6452;
    wire [63:0] _6458;
    wire [63:0] _155;
    reg [63:0] _3231;
    wire _3233;
    wire _3234;
    wire _3228;
    wire _3235;
    wire _3238;
    wire [63:0] _3266;
    wire [63:0] _3264;
    wire [63:0] _3267;
    wire [63:0] _3281;
    wire [63:0] _6459;
    wire [63:0] _6465;
    wire [63:0] _156;
    reg [63:0] _3251;
    wire _3253;
    wire _3254;
    wire _3248;
    wire _3255;
    wire _3258;
    wire [63:0] _3286;
    wire [63:0] _3284;
    wire [63:0] _3287;
    wire [63:0] _3301;
    wire [63:0] _6466;
    wire [63:0] _6472;
    wire [63:0] _157;
    reg [63:0] _3271;
    wire _3273;
    wire _3274;
    wire _3268;
    wire _3275;
    wire _3278;
    wire [63:0] _3306;
    wire [63:0] _3304;
    wire [63:0] _3307;
    wire [63:0] _3321;
    wire [63:0] _6473;
    wire [63:0] _6479;
    wire [63:0] _158;
    reg [63:0] _3291;
    wire _3293;
    wire _3294;
    wire _3288;
    wire _3295;
    wire _3298;
    wire [63:0] _3326;
    wire [63:0] _3324;
    wire [63:0] _3327;
    wire [63:0] _3341;
    wire [63:0] _6480;
    wire [63:0] _6486;
    wire [63:0] _159;
    reg [63:0] _3311;
    wire _3313;
    wire _3314;
    wire _3308;
    wire _3315;
    wire _3318;
    wire [63:0] _3346;
    wire [63:0] _3344;
    wire [63:0] _3347;
    wire [63:0] _3361;
    wire [63:0] _6487;
    wire [63:0] _6493;
    wire [63:0] _160;
    reg [63:0] _3331;
    wire _3333;
    wire _3334;
    wire _3328;
    wire _3335;
    wire _3338;
    wire [63:0] _3366;
    wire [63:0] _3364;
    wire [63:0] _3367;
    wire [63:0] _3381;
    wire [63:0] _6494;
    wire [63:0] _6500;
    wire [63:0] _161;
    reg [63:0] _3351;
    wire _3353;
    wire _3354;
    wire _3348;
    wire _3355;
    wire _3358;
    wire [63:0] _3386;
    wire [63:0] _3384;
    wire [63:0] _3387;
    wire [63:0] _3401;
    wire [63:0] _6501;
    wire [63:0] _6507;
    wire [63:0] _162;
    reg [63:0] _3371;
    wire _3373;
    wire _3374;
    wire _3368;
    wire _3375;
    wire _3378;
    wire [63:0] _3406;
    wire [63:0] _3404;
    wire [63:0] _3407;
    wire [63:0] _3421;
    wire [63:0] _6508;
    wire [63:0] _6514;
    wire [63:0] _163;
    reg [63:0] _3391;
    wire _3393;
    wire _3394;
    wire _3388;
    wire _3395;
    wire _3398;
    wire [63:0] _3426;
    wire [63:0] _3424;
    wire [63:0] _3427;
    wire [63:0] _3441;
    wire [63:0] _6515;
    wire [63:0] _6521;
    wire [63:0] _164;
    reg [63:0] _3411;
    wire _3413;
    wire _3414;
    wire _3408;
    wire _3415;
    wire _3418;
    wire [63:0] _3446;
    wire [63:0] _3444;
    wire [63:0] _3447;
    wire [63:0] _3461;
    wire [63:0] _6522;
    wire [63:0] _6528;
    wire [63:0] _165;
    reg [63:0] _3431;
    wire _3433;
    wire _3434;
    wire _3428;
    wire _3435;
    wire _3438;
    wire [63:0] _3466;
    wire [63:0] _3464;
    wire [63:0] _3467;
    wire [63:0] _3481;
    wire [63:0] _6529;
    wire [63:0] _6535;
    wire [63:0] _166;
    reg [63:0] _3451;
    wire _3453;
    wire _3454;
    wire _3448;
    wire _3455;
    wire _3458;
    wire [63:0] _3486;
    wire [63:0] _3484;
    wire [63:0] _3487;
    wire [63:0] _3501;
    wire [63:0] _6536;
    wire [63:0] _6542;
    wire [63:0] _167;
    reg [63:0] _3471;
    wire _3473;
    wire _3474;
    wire _3468;
    wire _3475;
    wire _3478;
    wire [63:0] _3506;
    wire [63:0] _3504;
    wire [63:0] _3507;
    wire [63:0] _3521;
    wire [63:0] _6543;
    wire [63:0] _6549;
    wire [63:0] _168;
    reg [63:0] _3491;
    wire _3493;
    wire _3494;
    wire _3488;
    wire _3495;
    wire _3498;
    wire [63:0] _3526;
    wire [63:0] _3524;
    wire [63:0] _3527;
    wire [63:0] _3541;
    wire [63:0] _6550;
    wire [63:0] _6556;
    wire [63:0] _169;
    reg [63:0] _3511;
    wire _3513;
    wire _3514;
    wire _3508;
    wire _3515;
    wire _3518;
    wire [63:0] _3546;
    wire [63:0] _3544;
    wire [63:0] _3547;
    wire [63:0] _3561;
    wire [63:0] _6557;
    wire [63:0] _6563;
    wire [63:0] _170;
    reg [63:0] _3531;
    wire _3533;
    wire _3534;
    wire _3528;
    wire _3535;
    wire _3538;
    wire [63:0] _3566;
    wire [63:0] _3564;
    wire [63:0] _3567;
    wire [63:0] _3581;
    wire [63:0] _6564;
    wire [63:0] _6570;
    wire [63:0] _171;
    reg [63:0] _3551;
    wire _3553;
    wire _3554;
    wire _3548;
    wire _3555;
    wire _3558;
    wire [63:0] _3586;
    wire [63:0] _3584;
    wire [63:0] _3587;
    wire [63:0] _3601;
    wire [63:0] _6571;
    wire [63:0] _6577;
    wire [63:0] _172;
    reg [63:0] _3571;
    wire _3573;
    wire _3574;
    wire _3568;
    wire _3575;
    wire _3578;
    wire [63:0] _3606;
    wire [63:0] _3604;
    wire [63:0] _3607;
    wire [63:0] _3621;
    wire [63:0] _6578;
    wire [63:0] _6584;
    wire [63:0] _173;
    reg [63:0] _3591;
    wire _3593;
    wire _3594;
    wire _3588;
    wire _3595;
    wire _3598;
    wire [63:0] _3626;
    wire [63:0] _3624;
    wire [63:0] _3627;
    wire [63:0] _3641;
    wire [63:0] _6585;
    wire [63:0] _6591;
    wire [63:0] _174;
    reg [63:0] _3611;
    wire _3613;
    wire _3614;
    wire _3608;
    wire _3615;
    wire _3618;
    wire [63:0] _3646;
    wire [63:0] _3644;
    wire [63:0] _3647;
    wire [63:0] _3661;
    wire [63:0] _6592;
    wire [63:0] _6598;
    wire [63:0] _175;
    reg [63:0] _3631;
    wire _3633;
    wire _3634;
    wire _3628;
    wire _3635;
    wire _3638;
    wire [63:0] _3666;
    wire [63:0] _3664;
    wire [63:0] _3667;
    wire [63:0] _3681;
    wire [63:0] _6599;
    wire [63:0] _6605;
    wire [63:0] _176;
    reg [63:0] _3651;
    wire _3653;
    wire _3654;
    wire _3648;
    wire _3655;
    wire _3658;
    wire [63:0] _3686;
    wire [63:0] _3684;
    wire [63:0] _3687;
    wire [63:0] _3701;
    wire [63:0] _6606;
    wire [63:0] _6612;
    wire [63:0] _177;
    reg [63:0] _3671;
    wire _3673;
    wire _3674;
    wire _3668;
    wire _3675;
    wire _3678;
    wire [63:0] _3706;
    wire [63:0] _3704;
    wire [63:0] _3707;
    wire [63:0] _3721;
    wire [63:0] _6613;
    wire [63:0] _6619;
    wire [63:0] _178;
    reg [63:0] _3691;
    wire _3693;
    wire _3694;
    wire _3688;
    wire _3695;
    wire _3698;
    wire [63:0] _3726;
    wire [63:0] _3724;
    wire [63:0] _3727;
    wire [63:0] _3741;
    wire [63:0] _6620;
    wire [63:0] _6626;
    wire [63:0] _179;
    reg [63:0] _3711;
    wire _3713;
    wire _3714;
    wire _3708;
    wire _3715;
    wire _3718;
    wire [63:0] _3746;
    wire [63:0] _3744;
    wire [63:0] _3747;
    wire [63:0] _3761;
    wire [63:0] _6627;
    wire [63:0] _6633;
    wire [63:0] _180;
    reg [63:0] _3731;
    wire _3733;
    wire _3734;
    wire _3728;
    wire _3735;
    wire _3738;
    wire [63:0] _3766;
    wire [63:0] _3764;
    wire [63:0] _3767;
    wire [63:0] _3781;
    wire [63:0] _6634;
    wire [63:0] _6640;
    wire [63:0] _181;
    reg [63:0] _3751;
    wire _3753;
    wire _3754;
    wire _3748;
    wire _3755;
    wire _3758;
    wire [63:0] _3786;
    wire [63:0] _3784;
    wire [63:0] _3787;
    wire [63:0] _3801;
    wire [63:0] _6641;
    wire [63:0] _6647;
    wire [63:0] _182;
    reg [63:0] _3771;
    wire _3773;
    wire _3774;
    wire _3768;
    wire _3775;
    wire _3778;
    wire [63:0] _3806;
    wire [63:0] _3804;
    wire [63:0] _3807;
    wire [63:0] _3821;
    wire [63:0] _6648;
    wire [63:0] _6654;
    wire [63:0] _183;
    reg [63:0] _3791;
    wire _3793;
    wire _3794;
    wire _3788;
    wire _3795;
    wire _3798;
    wire [63:0] _3826;
    wire [63:0] _3824;
    wire [63:0] _3827;
    wire [63:0] _3841;
    wire [63:0] _6655;
    wire [63:0] _6661;
    wire [63:0] _184;
    reg [63:0] _3811;
    wire _3813;
    wire _3814;
    wire _3808;
    wire _3815;
    wire _3818;
    wire [63:0] _3846;
    wire [63:0] _3844;
    wire [63:0] _3847;
    wire [63:0] _3861;
    wire [63:0] _6662;
    wire [63:0] _6668;
    wire [63:0] _185;
    reg [63:0] _3831;
    wire _3833;
    wire _3834;
    wire _3828;
    wire _3835;
    wire _3838;
    wire [63:0] _3866;
    wire [63:0] _3864;
    wire [63:0] _3867;
    wire [63:0] _3881;
    wire [63:0] _6669;
    wire [63:0] _6675;
    wire [63:0] _186;
    reg [63:0] _3851;
    wire _3853;
    wire _3854;
    wire _3848;
    wire _3855;
    wire _3858;
    wire [63:0] _3886;
    wire [63:0] _3884;
    wire [63:0] _3887;
    wire [63:0] _3901;
    wire [63:0] _6676;
    wire [63:0] _6682;
    wire [63:0] _187;
    reg [63:0] _3871;
    wire _3873;
    wire _3874;
    wire _3868;
    wire _3875;
    wire _3878;
    wire [63:0] _3906;
    wire [63:0] _3904;
    wire [63:0] _3907;
    wire [63:0] _3921;
    wire [63:0] _6683;
    wire [63:0] _6689;
    wire [63:0] _188;
    reg [63:0] _3891;
    wire _3893;
    wire _3894;
    wire _3888;
    wire _3895;
    wire _3898;
    wire [63:0] _3926;
    wire [63:0] _3924;
    wire [63:0] _3927;
    wire [63:0] _3941;
    wire [63:0] _6690;
    wire [63:0] _6696;
    wire [63:0] _189;
    reg [63:0] _3911;
    wire _3913;
    wire _3914;
    wire _3908;
    wire _3915;
    wire _3918;
    wire [63:0] _3946;
    wire [63:0] _3944;
    wire [63:0] _3947;
    wire [63:0] _3961;
    wire [63:0] _6697;
    wire [63:0] _6703;
    wire [63:0] _190;
    reg [63:0] _3931;
    wire _3933;
    wire _3934;
    wire _3928;
    wire _3935;
    wire _3938;
    wire [63:0] _3966;
    wire [63:0] _3964;
    wire [63:0] _3967;
    wire [63:0] _3981;
    wire [63:0] _6704;
    wire [63:0] _6710;
    wire [63:0] _191;
    reg [63:0] _3951;
    wire _3953;
    wire _3954;
    wire _3948;
    wire _3955;
    wire _3958;
    wire [63:0] _3986;
    wire [63:0] _3984;
    wire [63:0] _3987;
    wire [63:0] _4001;
    wire [63:0] _6711;
    wire [63:0] _6717;
    wire [63:0] _192;
    reg [63:0] _3971;
    wire _3973;
    wire _3974;
    wire _3968;
    wire _3975;
    wire _3978;
    wire [63:0] _4006;
    wire [63:0] _4004;
    wire [63:0] _4007;
    wire [63:0] _4021;
    wire [63:0] _6718;
    wire [63:0] _6724;
    wire [63:0] _193;
    reg [63:0] _3991;
    wire _3993;
    wire _3994;
    wire _3988;
    wire _3995;
    wire _3998;
    wire [63:0] _4026;
    wire [63:0] _4024;
    wire [63:0] _4027;
    wire [63:0] _4041;
    wire [63:0] _6725;
    wire [63:0] _6731;
    wire [63:0] _194;
    reg [63:0] _4011;
    wire _4013;
    wire _4014;
    wire _4008;
    wire _4015;
    wire _4018;
    wire [63:0] _4046;
    wire [63:0] _4044;
    wire [63:0] _4047;
    wire [63:0] _4061;
    wire [63:0] _6732;
    wire [63:0] _6738;
    wire [63:0] _195;
    reg [63:0] _4031;
    wire _4033;
    wire _4034;
    wire _4028;
    wire _4035;
    wire _4038;
    wire [63:0] _4066;
    wire [63:0] _4064;
    wire [63:0] _4067;
    wire [63:0] _4081;
    wire [63:0] _6739;
    wire [63:0] _6745;
    wire [63:0] _196;
    reg [63:0] _4051;
    wire _4053;
    wire _4054;
    wire _4048;
    wire _4055;
    wire _4058;
    wire [63:0] _4086;
    wire [63:0] _4084;
    wire [63:0] _4087;
    wire [63:0] _4101;
    wire [63:0] _6746;
    wire [63:0] _6752;
    wire [63:0] _197;
    reg [63:0] _4071;
    wire _4073;
    wire _4074;
    wire _4068;
    wire _4075;
    wire _4078;
    wire [63:0] _4106;
    wire [63:0] _4104;
    wire [63:0] _4107;
    wire [63:0] _4121;
    wire [63:0] _6753;
    wire [63:0] _6759;
    wire [63:0] _198;
    reg [63:0] _4091;
    wire _4093;
    wire _4094;
    wire _4088;
    wire _4095;
    wire _4098;
    wire [63:0] _4126;
    wire [63:0] _4124;
    wire [63:0] _4127;
    wire [63:0] _4141;
    wire [63:0] _6760;
    wire [63:0] _6766;
    wire [63:0] _199;
    reg [63:0] _4111;
    wire _4113;
    wire _4114;
    wire _4108;
    wire _4115;
    wire _4118;
    wire [63:0] _4146;
    wire [63:0] _4144;
    wire [63:0] _4147;
    wire [63:0] _4161;
    wire [63:0] _6767;
    wire [63:0] _6773;
    wire [63:0] _200;
    reg [63:0] _4131;
    wire _4133;
    wire _4134;
    wire _4128;
    wire _4135;
    wire _4138;
    wire [63:0] _4166;
    wire [63:0] _4164;
    wire [63:0] _4167;
    wire [63:0] _4181;
    wire [63:0] _6774;
    wire [63:0] _6780;
    wire [63:0] _201;
    reg [63:0] _4151;
    wire _4153;
    wire _4154;
    wire _4148;
    wire _4155;
    wire _4158;
    wire [63:0] _4186;
    wire [63:0] _4184;
    wire [63:0] _4187;
    wire [63:0] _4201;
    wire [63:0] _6781;
    wire [63:0] _6787;
    wire [63:0] _202;
    reg [63:0] _4171;
    wire _4173;
    wire _4174;
    wire _4168;
    wire _4175;
    wire _4178;
    wire [63:0] _4206;
    wire [63:0] _4204;
    wire [63:0] _4207;
    wire [63:0] _4221;
    wire [63:0] _6788;
    wire [63:0] _6794;
    wire [63:0] _203;
    reg [63:0] _4191;
    wire _4193;
    wire _4194;
    wire _4188;
    wire _4195;
    wire _4198;
    wire [63:0] _4226;
    wire [63:0] _4224;
    wire [63:0] _4227;
    wire [63:0] _4241;
    wire [63:0] _6795;
    wire [63:0] _6801;
    wire [63:0] _204;
    reg [63:0] _4211;
    wire _4213;
    wire _4214;
    wire _4208;
    wire _4215;
    wire _4218;
    wire [63:0] _4246;
    wire [63:0] _4244;
    wire [63:0] _4247;
    wire [63:0] _4261;
    wire [63:0] _6802;
    wire [63:0] _6808;
    wire [63:0] _205;
    reg [63:0] _4231;
    wire _4233;
    wire _4234;
    wire _4228;
    wire _4235;
    wire _4238;
    wire [63:0] _4266;
    wire [63:0] _4264;
    wire [63:0] _4267;
    wire [63:0] _4281;
    wire [63:0] _6809;
    wire [63:0] _6815;
    wire [63:0] _206;
    reg [63:0] _4251;
    wire _4253;
    wire _4254;
    wire _4248;
    wire _4255;
    wire _4258;
    wire [63:0] _4286;
    wire [63:0] _4284;
    wire [63:0] _4287;
    wire [63:0] _4301;
    wire [63:0] _6816;
    wire [63:0] _6822;
    wire [63:0] _207;
    reg [63:0] _4271;
    wire _4273;
    wire _4274;
    wire _4268;
    wire _4275;
    wire _4278;
    wire [63:0] _4306;
    wire [63:0] _4304;
    wire [63:0] _4307;
    wire [63:0] _4321;
    wire [63:0] _6823;
    wire [63:0] _6829;
    wire [63:0] _208;
    reg [63:0] _4291;
    wire _4293;
    wire _4294;
    wire _4288;
    wire _4295;
    wire _4298;
    wire [63:0] _4326;
    wire [63:0] _4324;
    wire [63:0] _4327;
    wire [63:0] _4341;
    wire [63:0] _6830;
    wire [63:0] _6836;
    wire [63:0] _209;
    reg [63:0] _4311;
    wire _4313;
    wire _4314;
    wire _4308;
    wire _4315;
    wire _4318;
    wire [63:0] _4346;
    wire [63:0] _4344;
    wire [63:0] _4347;
    wire [63:0] _4361;
    wire [63:0] _6837;
    wire [63:0] _6843;
    wire [63:0] _210;
    reg [63:0] _4331;
    wire _4333;
    wire _4334;
    wire _4328;
    wire _4335;
    wire _4338;
    wire [63:0] _4366;
    wire [63:0] _4364;
    wire [63:0] _4367;
    wire [63:0] _4381;
    wire [63:0] _6844;
    wire [63:0] _6850;
    wire [63:0] _211;
    reg [63:0] _4351;
    wire _4353;
    wire _4354;
    wire _4348;
    wire _4355;
    wire _4358;
    wire [63:0] _4386;
    wire [63:0] _4384;
    wire [63:0] _4387;
    wire [63:0] _4401;
    wire [63:0] _6851;
    wire [63:0] _6857;
    wire [63:0] _212;
    reg [63:0] _4371;
    wire _4373;
    wire _4374;
    wire _4368;
    wire _4375;
    wire _4378;
    wire [63:0] _4406;
    wire [63:0] _4404;
    wire [63:0] _4407;
    wire [63:0] _4421;
    wire [63:0] _6858;
    wire [63:0] _6864;
    wire [63:0] _213;
    reg [63:0] _4391;
    wire _4393;
    wire _4394;
    wire _4388;
    wire _4395;
    wire _4398;
    wire [63:0] _4426;
    wire [63:0] _4424;
    wire [63:0] _4427;
    wire [63:0] _4441;
    wire [63:0] _6865;
    wire [63:0] _6871;
    wire [63:0] _214;
    reg [63:0] _4411;
    wire _4413;
    wire _4414;
    wire _4408;
    wire _4415;
    wire _4418;
    wire [63:0] _4446;
    wire [63:0] _4444;
    wire [63:0] _4447;
    wire [63:0] _4461;
    wire [63:0] _6872;
    wire [63:0] _6878;
    wire [63:0] _215;
    reg [63:0] _4431;
    wire _4433;
    wire _4434;
    wire _4428;
    wire _4435;
    wire _4438;
    wire [63:0] _4466;
    wire [63:0] _4464;
    wire [63:0] _4467;
    wire [63:0] _4481;
    wire [63:0] _6879;
    wire [63:0] _6885;
    wire [63:0] _216;
    reg [63:0] _4451;
    wire _4453;
    wire _4454;
    wire _4448;
    wire _4455;
    wire _4458;
    wire [63:0] _4486;
    wire [63:0] _4484;
    wire [63:0] _4487;
    wire [63:0] _4501;
    wire [63:0] _6886;
    wire [63:0] _6892;
    wire [63:0] _217;
    reg [63:0] _4471;
    wire _4473;
    wire _4474;
    wire _4468;
    wire _4475;
    wire _4478;
    wire [63:0] _4506;
    wire [63:0] _4504;
    wire [63:0] _4507;
    wire [63:0] _4521;
    wire [63:0] _6893;
    wire [63:0] _6899;
    wire [63:0] _218;
    reg [63:0] _4491;
    wire _4493;
    wire _4494;
    wire _4488;
    wire _4495;
    wire _4498;
    wire [63:0] _4526;
    wire [63:0] _4524;
    wire [63:0] _4527;
    wire [63:0] _4541;
    wire [63:0] _6900;
    wire [63:0] _6906;
    wire [63:0] _219;
    reg [63:0] _4511;
    wire _4513;
    wire _4514;
    wire _4508;
    wire _4515;
    wire _4518;
    wire [63:0] _4546;
    wire [63:0] _4544;
    wire [63:0] _4547;
    wire [63:0] _4561;
    wire [63:0] _6907;
    wire [63:0] _6913;
    wire [63:0] _220;
    reg [63:0] _4531;
    wire _4533;
    wire _4534;
    wire _4528;
    wire _4535;
    wire _4538;
    wire [63:0] _4566;
    wire [63:0] _4564;
    wire [63:0] _4567;
    wire [63:0] _4581;
    wire [63:0] _6914;
    wire [63:0] _6920;
    wire [63:0] _221;
    reg [63:0] _4551;
    wire _4553;
    wire _4554;
    wire _4548;
    wire _4555;
    wire _4558;
    wire [63:0] _4586;
    wire [63:0] _4584;
    wire [63:0] _4587;
    wire [63:0] _4601;
    wire [63:0] _6921;
    wire [63:0] _6927;
    wire [63:0] _222;
    reg [63:0] _4571;
    wire _4573;
    wire _4574;
    wire _4568;
    wire _4575;
    wire _4578;
    wire [63:0] _4606;
    wire [63:0] _4604;
    wire [63:0] _4607;
    wire [63:0] _4621;
    wire [63:0] _6928;
    wire [63:0] _6934;
    wire [63:0] _223;
    reg [63:0] _4591;
    wire _4593;
    wire _4594;
    wire _4588;
    wire _4595;
    wire _4598;
    wire [63:0] _4626;
    wire [63:0] _4624;
    wire [63:0] _4627;
    wire [63:0] _4641;
    wire [63:0] _6935;
    wire [63:0] _6941;
    wire [63:0] _224;
    reg [63:0] _4611;
    wire _4613;
    wire _4614;
    wire _4608;
    wire _4615;
    wire _4618;
    wire [63:0] _4646;
    wire [63:0] _4644;
    wire [63:0] _4647;
    wire [63:0] _4661;
    wire [63:0] _6942;
    wire [63:0] _6948;
    wire [63:0] _225;
    reg [63:0] _4631;
    wire _4633;
    wire _4634;
    wire _4628;
    wire _4635;
    wire _4638;
    wire [63:0] _4666;
    wire [63:0] _4664;
    wire [63:0] _4667;
    wire [63:0] _4681;
    wire [63:0] _6949;
    wire [63:0] _6955;
    wire [63:0] _226;
    reg [63:0] _4651;
    wire _4653;
    wire _4654;
    wire _4648;
    wire _4655;
    wire _4658;
    wire [63:0] _4686;
    wire [63:0] _4684;
    wire [63:0] _4687;
    wire [63:0] _4701;
    wire [63:0] _6956;
    wire [63:0] _6962;
    wire [63:0] _227;
    reg [63:0] _4671;
    wire _4673;
    wire _4674;
    wire _4668;
    wire _4675;
    wire _4678;
    wire [63:0] _4706;
    wire [63:0] _4704;
    wire [63:0] _4707;
    wire [63:0] _4721;
    wire [63:0] _6963;
    wire [63:0] _6969;
    wire [63:0] _228;
    reg [63:0] _4691;
    wire _4693;
    wire _4694;
    wire _4688;
    wire _4695;
    wire _4698;
    wire [63:0] _4726;
    wire [63:0] _4724;
    wire [63:0] _4727;
    wire [63:0] _4741;
    wire [63:0] _6970;
    wire [63:0] _6976;
    wire [63:0] _229;
    reg [63:0] _4711;
    wire _4713;
    wire _4714;
    wire _4708;
    wire _4715;
    wire _4718;
    wire [63:0] _4746;
    wire [63:0] _4744;
    wire [63:0] _4747;
    wire [63:0] _4761;
    wire [63:0] _6977;
    wire [63:0] _6983;
    wire [63:0] _230;
    reg [63:0] _4731;
    wire _4733;
    wire _4734;
    wire _4728;
    wire _4735;
    wire _4738;
    wire [63:0] _4766;
    wire [63:0] _4764;
    wire [63:0] _4767;
    wire [63:0] _4781;
    wire [63:0] _6984;
    wire [63:0] _6990;
    wire [63:0] _231;
    reg [63:0] _4751;
    wire _4753;
    wire _4754;
    wire _4748;
    wire _4755;
    wire _4758;
    wire [63:0] _4786;
    wire [63:0] _4784;
    wire [63:0] _4787;
    wire [63:0] _4801;
    wire [63:0] _6991;
    wire [63:0] _6997;
    wire [63:0] _232;
    reg [63:0] _4771;
    wire _4773;
    wire _4774;
    wire _4768;
    wire _4775;
    wire _4778;
    wire [63:0] _4806;
    wire [63:0] _4804;
    wire [63:0] _4807;
    wire [63:0] _4821;
    wire [63:0] _6998;
    wire [63:0] _7004;
    wire [63:0] _233;
    reg [63:0] _4791;
    wire _4793;
    wire _4794;
    wire _4788;
    wire _4795;
    wire _4798;
    wire [63:0] _4826;
    wire [63:0] _4824;
    wire [63:0] _4827;
    wire [63:0] _4841;
    wire [63:0] _7005;
    wire [63:0] _7011;
    wire [63:0] _234;
    reg [63:0] _4811;
    wire _4813;
    wire _4814;
    wire _4808;
    wire _4815;
    wire _4818;
    wire [63:0] _4846;
    wire [63:0] _4844;
    wire [63:0] _4847;
    wire [63:0] _4861;
    wire [63:0] _7012;
    wire [63:0] _7018;
    wire [63:0] _235;
    reg [63:0] _4831;
    wire _4833;
    wire _4834;
    wire _4828;
    wire _4835;
    wire _4838;
    wire [63:0] _4866;
    wire [63:0] _4864;
    wire [63:0] _4867;
    wire [63:0] _4881;
    wire [63:0] _7019;
    wire [63:0] _7025;
    wire [63:0] _236;
    reg [63:0] _4851;
    wire _4853;
    wire _4854;
    wire _4848;
    wire _4855;
    wire _4858;
    wire [63:0] _4886;
    wire [63:0] _4884;
    wire [63:0] _4887;
    wire [63:0] _4901;
    wire [63:0] _7026;
    wire [63:0] _7032;
    wire [63:0] _237;
    reg [63:0] _4871;
    wire _4873;
    wire _4874;
    wire _4868;
    wire _4875;
    wire _4878;
    wire [63:0] _4906;
    wire [63:0] _4904;
    wire [63:0] _4907;
    wire [63:0] _4921;
    wire [63:0] _7033;
    wire [63:0] _7039;
    wire [63:0] _238;
    reg [63:0] _4891;
    wire _4893;
    wire _4894;
    wire _4888;
    wire _4895;
    wire _4898;
    wire [63:0] _4926;
    wire [63:0] _4924;
    wire [63:0] _4927;
    wire [63:0] _4941;
    wire [63:0] _7040;
    wire [63:0] _7046;
    wire [63:0] _239;
    reg [63:0] _4911;
    wire _4913;
    wire _4914;
    wire _4908;
    wire _4915;
    wire _4918;
    wire [63:0] _4946;
    wire [63:0] _4944;
    wire [63:0] _4947;
    wire [63:0] _4961;
    wire [63:0] _7047;
    wire [63:0] _7053;
    wire [63:0] _240;
    reg [63:0] _4931;
    wire _4933;
    wire _4934;
    wire _4928;
    wire _4935;
    wire _4938;
    wire [63:0] _4966;
    wire [63:0] _4964;
    wire [63:0] _4967;
    wire [63:0] _4981;
    wire [63:0] _7054;
    wire [63:0] _7060;
    wire [63:0] _241;
    reg [63:0] _4951;
    wire _4953;
    wire _4954;
    wire _4948;
    wire _4955;
    wire _4958;
    wire [63:0] _4986;
    wire [63:0] _4984;
    wire [63:0] _4987;
    wire [63:0] _5001;
    wire [63:0] _7061;
    wire [63:0] _7067;
    wire [63:0] _242;
    reg [63:0] _4971;
    wire _4973;
    wire _4974;
    wire _4968;
    wire _4975;
    wire _4978;
    wire [63:0] _5006;
    wire [63:0] _5004;
    wire [63:0] _5007;
    wire [63:0] _5021;
    wire [63:0] _7068;
    wire [63:0] _7074;
    wire [63:0] _243;
    reg [63:0] _4991;
    wire _4993;
    wire _4994;
    wire _4988;
    wire _4995;
    wire _4998;
    wire [63:0] _5026;
    wire [63:0] _5024;
    wire [63:0] _5027;
    wire [63:0] _5041;
    wire [63:0] _7075;
    wire [63:0] _7081;
    wire [63:0] _244;
    reg [63:0] _5011;
    wire _5013;
    wire _5014;
    wire _5008;
    wire _5015;
    wire _5018;
    wire [63:0] _5046;
    wire [63:0] _5044;
    wire [63:0] _5047;
    wire [63:0] _5061;
    wire [63:0] _7082;
    wire [63:0] _7088;
    wire [63:0] _245;
    reg [63:0] _5031;
    wire _5033;
    wire _5034;
    wire _5028;
    wire _5035;
    wire _5038;
    wire [63:0] _5066;
    wire [63:0] _5064;
    wire [63:0] _5067;
    wire [63:0] _5081;
    wire [63:0] _7089;
    wire [63:0] _7095;
    wire [63:0] _246;
    reg [63:0] _5051;
    wire _5053;
    wire _5054;
    wire _5048;
    wire _5055;
    wire _5058;
    wire [63:0] _5086;
    wire [63:0] _5084;
    wire [63:0] _5087;
    wire [63:0] _5101;
    wire [63:0] _7096;
    wire [63:0] _7102;
    wire [63:0] _247;
    reg [63:0] _5071;
    wire _5073;
    wire _5074;
    wire _5068;
    wire _5075;
    wire _5078;
    wire [63:0] _5106;
    wire [63:0] _5104;
    wire [63:0] _5107;
    wire [63:0] _5121;
    wire [63:0] _7103;
    wire [63:0] _7109;
    wire [63:0] _248;
    reg [63:0] _5091;
    wire _5093;
    wire _5094;
    wire _5088;
    wire _5095;
    wire _5098;
    wire [63:0] _5126;
    wire [63:0] _5124;
    wire [63:0] _5127;
    wire [63:0] _5141;
    wire [63:0] _7110;
    wire [63:0] _7116;
    wire [63:0] _249;
    reg [63:0] _5111;
    wire _5113;
    wire _5114;
    wire _5108;
    wire _5115;
    wire _5118;
    wire [63:0] _5146;
    wire [63:0] _5144;
    wire [63:0] _5147;
    wire [63:0] _5161;
    wire [63:0] _7117;
    wire [63:0] _7123;
    wire [63:0] _250;
    reg [63:0] _5131;
    wire _5133;
    wire _5134;
    wire _5128;
    wire _5135;
    wire _5138;
    wire [63:0] _5166;
    wire [63:0] _5164;
    wire [63:0] _5167;
    wire [63:0] _5181;
    wire [63:0] _7124;
    wire [63:0] _7130;
    wire [63:0] _251;
    reg [63:0] _5151;
    wire _5153;
    wire _5154;
    wire _5148;
    wire _5155;
    wire _5158;
    wire [63:0] _5186;
    wire [63:0] _5184;
    wire [63:0] _5187;
    wire [63:0] _5201;
    wire [63:0] _7131;
    wire [63:0] _7137;
    wire [63:0] _252;
    reg [63:0] _5171;
    wire _5173;
    wire _5174;
    wire _5168;
    wire _5175;
    wire _5178;
    wire [63:0] _5206;
    wire [63:0] _5204;
    wire [63:0] _5207;
    wire [63:0] _5221;
    wire [63:0] _7138;
    wire [63:0] _7144;
    wire [63:0] _253;
    reg [63:0] _5191;
    wire _5193;
    wire _5194;
    wire _5188;
    wire _5195;
    wire _5198;
    wire [63:0] _5226;
    wire [63:0] _5224;
    wire [63:0] _5227;
    wire [63:0] _5241;
    wire [63:0] _7145;
    wire [63:0] _7151;
    wire [63:0] _254;
    reg [63:0] _5211;
    wire _5213;
    wire _5214;
    wire _5208;
    wire _5215;
    wire _5218;
    wire [63:0] _5246;
    wire [63:0] _5244;
    wire [63:0] _5247;
    wire [63:0] _5261;
    wire [63:0] _7152;
    wire [63:0] _7158;
    wire [63:0] _255;
    reg [63:0] _5231;
    wire _5233;
    wire _5234;
    wire _5228;
    wire _5235;
    wire _5238;
    wire [63:0] _5266;
    wire [63:0] _5264;
    wire [63:0] _5267;
    wire [63:0] _5281;
    wire [63:0] _7159;
    wire [63:0] _7165;
    wire [63:0] _256;
    reg [63:0] _5251;
    wire _5253;
    wire _5254;
    wire _5248;
    wire _5255;
    wire _5258;
    wire [63:0] _5286;
    wire [63:0] _5284;
    wire [63:0] _5287;
    wire [63:0] _5301;
    wire [63:0] _7166;
    wire [63:0] _7172;
    wire [63:0] _257;
    reg [63:0] _5271;
    wire _5273;
    wire _5274;
    wire _5268;
    wire _5275;
    wire _5278;
    wire [63:0] _5306;
    wire [63:0] _5304;
    wire [63:0] _5307;
    wire [63:0] _5321;
    wire [63:0] _7173;
    wire [63:0] _7179;
    wire [63:0] _258;
    reg [63:0] _5291;
    wire _5293;
    wire _5294;
    wire _5288;
    wire _5295;
    wire _5298;
    wire [63:0] _5326;
    wire [63:0] _5324;
    wire [63:0] _5327;
    wire [63:0] _5341;
    wire [63:0] _7180;
    wire [63:0] _7186;
    wire [63:0] _259;
    reg [63:0] _5311;
    wire _5313;
    wire _5314;
    wire _5308;
    wire _5315;
    wire _5318;
    wire [63:0] _5346;
    wire [63:0] _5344;
    wire [63:0] _5347;
    wire [63:0] _5361;
    wire [63:0] _7187;
    wire [63:0] _7193;
    wire [63:0] _260;
    reg [63:0] _5331;
    wire _5333;
    wire _5334;
    wire _5328;
    wire _5335;
    wire _5338;
    wire [63:0] _5366;
    wire [63:0] _5364;
    wire [63:0] _5367;
    wire [63:0] _5381;
    wire [63:0] _7194;
    wire [63:0] _7200;
    wire [63:0] _261;
    reg [63:0] _5351;
    wire _5353;
    wire _5354;
    wire _5348;
    wire _5355;
    wire _5358;
    wire [63:0] _5386;
    wire [63:0] _5384;
    wire [63:0] _5387;
    wire [63:0] _5401;
    wire [63:0] _7201;
    wire [63:0] _7207;
    wire [63:0] _262;
    reg [63:0] _5371;
    wire _5373;
    wire _5374;
    wire _5368;
    wire _5375;
    wire _5378;
    wire [63:0] _5406;
    wire [63:0] _5404;
    wire [63:0] _5407;
    wire [63:0] _7208;
    wire [63:0] _7214;
    wire [63:0] _263;
    reg [63:0] _5391;
    wire _5393;
    wire _5394;
    wire [255:0] _265;
    wire _5388;
    wire _5395;
    wire _5398;
    wire [255:0] _7220;
    wire _7221;
    wire [8:0] _7222;
    wire [8:0] _7226;
    wire [8:0] _7234;
    wire [8:0] _7250;
    wire [8:0] _7282;
    wire [8:0] _7346;
    wire [8:0] _7474;
    wire [8:0] _7730;
    wire [8:0] _8242;
    wire [54:0] _7218;
    wire [63:0] _8243;
    wire [63:0] _8244;
    wire [63:0] _8245;
    wire [63:0] _8247;
    wire [63:0] _266;
    reg [63:0] _7217;
    wire _8249;
    wire vdd;
    wire [1:0] _282;
    wire _270;
    wire _272;
    wire [1:0] _8248;
    wire _274;
    wire _276;
    wire _287;
    wire _8250;
    wire [1:0] _8251;
    wire _278;
    wire [1:0] _8252;
    wire [1:0] _279;
    reg [1:0] _284;
    wire _286;
    assign _290 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign _342 = _322 + _341;
    assign _362 = _342 + _361;
    assign _382 = _362 + _381;
    assign _402 = _382 + _401;
    assign _422 = _402 + _421;
    assign _442 = _422 + _441;
    assign _462 = _442 + _461;
    assign _482 = _462 + _481;
    assign _502 = _482 + _501;
    assign _522 = _502 + _521;
    assign _542 = _522 + _541;
    assign _562 = _542 + _561;
    assign _582 = _562 + _581;
    assign _602 = _582 + _601;
    assign _622 = _602 + _621;
    assign _642 = _622 + _641;
    assign _662 = _642 + _661;
    assign _682 = _662 + _681;
    assign _702 = _682 + _701;
    assign _722 = _702 + _721;
    assign _742 = _722 + _741;
    assign _762 = _742 + _761;
    assign _782 = _762 + _781;
    assign _802 = _782 + _801;
    assign _822 = _802 + _821;
    assign _842 = _822 + _841;
    assign _862 = _842 + _861;
    assign _882 = _862 + _881;
    assign _902 = _882 + _901;
    assign _922 = _902 + _921;
    assign _942 = _922 + _941;
    assign _962 = _942 + _961;
    assign _982 = _962 + _981;
    assign _1002 = _982 + _1001;
    assign _1022 = _1002 + _1021;
    assign _1042 = _1022 + _1041;
    assign _1062 = _1042 + _1061;
    assign _1082 = _1062 + _1081;
    assign _1102 = _1082 + _1101;
    assign _1122 = _1102 + _1121;
    assign _1142 = _1122 + _1141;
    assign _1162 = _1142 + _1161;
    assign _1182 = _1162 + _1181;
    assign _1202 = _1182 + _1201;
    assign _1222 = _1202 + _1221;
    assign _1242 = _1222 + _1241;
    assign _1262 = _1242 + _1261;
    assign _1282 = _1262 + _1281;
    assign _1302 = _1282 + _1301;
    assign _1322 = _1302 + _1321;
    assign _1342 = _1322 + _1341;
    assign _1362 = _1342 + _1361;
    assign _1382 = _1362 + _1381;
    assign _1402 = _1382 + _1401;
    assign _1422 = _1402 + _1421;
    assign _1442 = _1422 + _1441;
    assign _1462 = _1442 + _1461;
    assign _1482 = _1462 + _1481;
    assign _1502 = _1482 + _1501;
    assign _1522 = _1502 + _1521;
    assign _1542 = _1522 + _1541;
    assign _1562 = _1542 + _1561;
    assign _1582 = _1562 + _1581;
    assign _1602 = _1582 + _1601;
    assign _1622 = _1602 + _1621;
    assign _1642 = _1622 + _1641;
    assign _1662 = _1642 + _1661;
    assign _1682 = _1662 + _1681;
    assign _1702 = _1682 + _1701;
    assign _1722 = _1702 + _1721;
    assign _1742 = _1722 + _1741;
    assign _1762 = _1742 + _1761;
    assign _1782 = _1762 + _1781;
    assign _1802 = _1782 + _1801;
    assign _1822 = _1802 + _1821;
    assign _1842 = _1822 + _1841;
    assign _1862 = _1842 + _1861;
    assign _1882 = _1862 + _1881;
    assign _1902 = _1882 + _1901;
    assign _1922 = _1902 + _1921;
    assign _1942 = _1922 + _1941;
    assign _1962 = _1942 + _1961;
    assign _1982 = _1962 + _1981;
    assign _2002 = _1982 + _2001;
    assign _2022 = _2002 + _2021;
    assign _2042 = _2022 + _2041;
    assign _2062 = _2042 + _2061;
    assign _2082 = _2062 + _2081;
    assign _2102 = _2082 + _2101;
    assign _2122 = _2102 + _2121;
    assign _2142 = _2122 + _2141;
    assign _2162 = _2142 + _2161;
    assign _2182 = _2162 + _2181;
    assign _2202 = _2182 + _2201;
    assign _2222 = _2202 + _2221;
    assign _2242 = _2222 + _2241;
    assign _2262 = _2242 + _2261;
    assign _2282 = _2262 + _2281;
    assign _2302 = _2282 + _2301;
    assign _2322 = _2302 + _2321;
    assign _2342 = _2322 + _2341;
    assign _2362 = _2342 + _2361;
    assign _2382 = _2362 + _2381;
    assign _2402 = _2382 + _2401;
    assign _2422 = _2402 + _2421;
    assign _2442 = _2422 + _2441;
    assign _2462 = _2442 + _2461;
    assign _2482 = _2462 + _2481;
    assign _2502 = _2482 + _2501;
    assign _2522 = _2502 + _2521;
    assign _2542 = _2522 + _2541;
    assign _2562 = _2542 + _2561;
    assign _2582 = _2562 + _2581;
    assign _2602 = _2582 + _2601;
    assign _2622 = _2602 + _2621;
    assign _2642 = _2622 + _2641;
    assign _2662 = _2642 + _2661;
    assign _2682 = _2662 + _2681;
    assign _2702 = _2682 + _2701;
    assign _2722 = _2702 + _2721;
    assign _2742 = _2722 + _2741;
    assign _2762 = _2742 + _2761;
    assign _2782 = _2762 + _2781;
    assign _2802 = _2782 + _2801;
    assign _2822 = _2802 + _2821;
    assign _2842 = _2822 + _2841;
    assign _2862 = _2842 + _2861;
    assign _2882 = _2862 + _2881;
    assign _2902 = _2882 + _2901;
    assign _2922 = _2902 + _2921;
    assign _2942 = _2922 + _2941;
    assign _2962 = _2942 + _2961;
    assign _2982 = _2962 + _2981;
    assign _3002 = _2982 + _3001;
    assign _3022 = _3002 + _3021;
    assign _3042 = _3022 + _3041;
    assign _3062 = _3042 + _3061;
    assign _3082 = _3062 + _3081;
    assign _3102 = _3082 + _3101;
    assign _3122 = _3102 + _3121;
    assign _3142 = _3122 + _3141;
    assign _3162 = _3142 + _3161;
    assign _3182 = _3162 + _3181;
    assign _3202 = _3182 + _3201;
    assign _3222 = _3202 + _3221;
    assign _3242 = _3222 + _3241;
    assign _3262 = _3242 + _3261;
    assign _3282 = _3262 + _3281;
    assign _3302 = _3282 + _3301;
    assign _3322 = _3302 + _3321;
    assign _3342 = _3322 + _3341;
    assign _3362 = _3342 + _3361;
    assign _3382 = _3362 + _3381;
    assign _3402 = _3382 + _3401;
    assign _3422 = _3402 + _3421;
    assign _3442 = _3422 + _3441;
    assign _3462 = _3442 + _3461;
    assign _3482 = _3462 + _3481;
    assign _3502 = _3482 + _3501;
    assign _3522 = _3502 + _3521;
    assign _3542 = _3522 + _3541;
    assign _3562 = _3542 + _3561;
    assign _3582 = _3562 + _3581;
    assign _3602 = _3582 + _3601;
    assign _3622 = _3602 + _3621;
    assign _3642 = _3622 + _3641;
    assign _3662 = _3642 + _3661;
    assign _3682 = _3662 + _3681;
    assign _3702 = _3682 + _3701;
    assign _3722 = _3702 + _3721;
    assign _3742 = _3722 + _3741;
    assign _3762 = _3742 + _3761;
    assign _3782 = _3762 + _3781;
    assign _3802 = _3782 + _3801;
    assign _3822 = _3802 + _3821;
    assign _3842 = _3822 + _3841;
    assign _3862 = _3842 + _3861;
    assign _3882 = _3862 + _3881;
    assign _3902 = _3882 + _3901;
    assign _3922 = _3902 + _3921;
    assign _3942 = _3922 + _3941;
    assign _3962 = _3942 + _3961;
    assign _3982 = _3962 + _3981;
    assign _4002 = _3982 + _4001;
    assign _4022 = _4002 + _4021;
    assign _4042 = _4022 + _4041;
    assign _4062 = _4042 + _4061;
    assign _4082 = _4062 + _4081;
    assign _4102 = _4082 + _4101;
    assign _4122 = _4102 + _4121;
    assign _4142 = _4122 + _4141;
    assign _4162 = _4142 + _4161;
    assign _4182 = _4162 + _4181;
    assign _4202 = _4182 + _4201;
    assign _4222 = _4202 + _4221;
    assign _4242 = _4222 + _4241;
    assign _4262 = _4242 + _4261;
    assign _4282 = _4262 + _4281;
    assign _4302 = _4282 + _4301;
    assign _4322 = _4302 + _4321;
    assign _4342 = _4322 + _4341;
    assign _4362 = _4342 + _4361;
    assign _4382 = _4362 + _4381;
    assign _4402 = _4382 + _4401;
    assign _4422 = _4402 + _4421;
    assign _4442 = _4422 + _4441;
    assign _4462 = _4442 + _4461;
    assign _4482 = _4462 + _4481;
    assign _4502 = _4482 + _4501;
    assign _4522 = _4502 + _4521;
    assign _4542 = _4522 + _4541;
    assign _4562 = _4542 + _4561;
    assign _4582 = _4562 + _4581;
    assign _4602 = _4582 + _4601;
    assign _4622 = _4602 + _4621;
    assign _4642 = _4622 + _4641;
    assign _4662 = _4642 + _4661;
    assign _4682 = _4662 + _4681;
    assign _4702 = _4682 + _4701;
    assign _4722 = _4702 + _4721;
    assign _4742 = _4722 + _4741;
    assign _4762 = _4742 + _4761;
    assign _4782 = _4762 + _4781;
    assign _4802 = _4782 + _4801;
    assign _4822 = _4802 + _4821;
    assign _4842 = _4822 + _4841;
    assign _4862 = _4842 + _4861;
    assign _4882 = _4862 + _4881;
    assign _4902 = _4882 + _4901;
    assign _4922 = _4902 + _4921;
    assign _4942 = _4922 + _4941;
    assign _4962 = _4942 + _4961;
    assign _4982 = _4962 + _4981;
    assign _5002 = _4982 + _5001;
    assign _5022 = _5002 + _5021;
    assign _5042 = _5022 + _5041;
    assign _5062 = _5042 + _5061;
    assign _5082 = _5062 + _5081;
    assign _5102 = _5082 + _5101;
    assign _5122 = _5102 + _5121;
    assign _5142 = _5122 + _5141;
    assign _5162 = _5142 + _5161;
    assign _5182 = _5162 + _5181;
    assign _5202 = _5182 + _5201;
    assign _5222 = _5202 + _5221;
    assign _5242 = _5222 + _5241;
    assign _5262 = _5242 + _5261;
    assign _5282 = _5262 + _5281;
    assign _5302 = _5282 + _5301;
    assign _5322 = _5302 + _5321;
    assign _5342 = _5322 + _5341;
    assign _5362 = _5342 + _5361;
    assign _5382 = _5362 + _5381;
    assign _5402 = _5382 + _5401;
    assign _5408 = _5402 + _5407;
    assign _288 = _287 & _274;
    assign _5409 = _288 ? _5408 : _291;
    assign _5411 = _278 ? _290 : _5409;
    assign _2 = _5411;
    always @(posedge _272) begin
        if (_270)
            _291 <= _290;
        else
            _291 <= _2;
    end
    assign _8233 = _7220[0:0];
    assign _8232 = 8'b00000000;
    assign _8234 = { _8232,
                     _8233 };
    assign _8230 = _7220[1:1];
    assign _8231 = { _8232,
                     _8230 };
    assign _8235 = _8231 + _8234;
    assign _8226 = _7220[2:2];
    assign _8227 = { _8232,
                     _8226 };
    assign _8223 = _7220[3:3];
    assign _8224 = { _8232,
                     _8223 };
    assign _8228 = _8224 + _8227;
    assign _8236 = _8228 + _8235;
    assign _8218 = _7220[4:4];
    assign _8219 = { _8232,
                     _8218 };
    assign _8215 = _7220[5:5];
    assign _8216 = { _8232,
                     _8215 };
    assign _8220 = _8216 + _8219;
    assign _8211 = _7220[6:6];
    assign _8212 = { _8232,
                     _8211 };
    assign _8208 = _7220[7:7];
    assign _8209 = { _8232,
                     _8208 };
    assign _8213 = _8209 + _8212;
    assign _8221 = _8213 + _8220;
    assign _8237 = _8221 + _8236;
    assign _8202 = _7220[8:8];
    assign _8203 = { _8232,
                     _8202 };
    assign _8199 = _7220[9:9];
    assign _8200 = { _8232,
                     _8199 };
    assign _8204 = _8200 + _8203;
    assign _8195 = _7220[10:10];
    assign _8196 = { _8232,
                     _8195 };
    assign _8192 = _7220[11:11];
    assign _8193 = { _8232,
                     _8192 };
    assign _8197 = _8193 + _8196;
    assign _8205 = _8197 + _8204;
    assign _8187 = _7220[12:12];
    assign _8188 = { _8232,
                     _8187 };
    assign _8184 = _7220[13:13];
    assign _8185 = { _8232,
                     _8184 };
    assign _8189 = _8185 + _8188;
    assign _8180 = _7220[14:14];
    assign _8181 = { _8232,
                     _8180 };
    assign _8177 = _7220[15:15];
    assign _8178 = { _8232,
                     _8177 };
    assign _8182 = _8178 + _8181;
    assign _8190 = _8182 + _8189;
    assign _8206 = _8190 + _8205;
    assign _8238 = _8206 + _8237;
    assign _8170 = _7220[16:16];
    assign _8171 = { _8232,
                     _8170 };
    assign _8167 = _7220[17:17];
    assign _8168 = { _8232,
                     _8167 };
    assign _8172 = _8168 + _8171;
    assign _8163 = _7220[18:18];
    assign _8164 = { _8232,
                     _8163 };
    assign _8160 = _7220[19:19];
    assign _8161 = { _8232,
                     _8160 };
    assign _8165 = _8161 + _8164;
    assign _8173 = _8165 + _8172;
    assign _8155 = _7220[20:20];
    assign _8156 = { _8232,
                     _8155 };
    assign _8152 = _7220[21:21];
    assign _8153 = { _8232,
                     _8152 };
    assign _8157 = _8153 + _8156;
    assign _8148 = _7220[22:22];
    assign _8149 = { _8232,
                     _8148 };
    assign _8145 = _7220[23:23];
    assign _8146 = { _8232,
                     _8145 };
    assign _8150 = _8146 + _8149;
    assign _8158 = _8150 + _8157;
    assign _8174 = _8158 + _8173;
    assign _8139 = _7220[24:24];
    assign _8140 = { _8232,
                     _8139 };
    assign _8136 = _7220[25:25];
    assign _8137 = { _8232,
                     _8136 };
    assign _8141 = _8137 + _8140;
    assign _8132 = _7220[26:26];
    assign _8133 = { _8232,
                     _8132 };
    assign _8129 = _7220[27:27];
    assign _8130 = { _8232,
                     _8129 };
    assign _8134 = _8130 + _8133;
    assign _8142 = _8134 + _8141;
    assign _8124 = _7220[28:28];
    assign _8125 = { _8232,
                     _8124 };
    assign _8121 = _7220[29:29];
    assign _8122 = { _8232,
                     _8121 };
    assign _8126 = _8122 + _8125;
    assign _8117 = _7220[30:30];
    assign _8118 = { _8232,
                     _8117 };
    assign _8114 = _7220[31:31];
    assign _8115 = { _8232,
                     _8114 };
    assign _8119 = _8115 + _8118;
    assign _8127 = _8119 + _8126;
    assign _8143 = _8127 + _8142;
    assign _8175 = _8143 + _8174;
    assign _8239 = _8175 + _8238;
    assign _8106 = _7220[32:32];
    assign _8107 = { _8232,
                     _8106 };
    assign _8103 = _7220[33:33];
    assign _8104 = { _8232,
                     _8103 };
    assign _8108 = _8104 + _8107;
    assign _8099 = _7220[34:34];
    assign _8100 = { _8232,
                     _8099 };
    assign _8096 = _7220[35:35];
    assign _8097 = { _8232,
                     _8096 };
    assign _8101 = _8097 + _8100;
    assign _8109 = _8101 + _8108;
    assign _8091 = _7220[36:36];
    assign _8092 = { _8232,
                     _8091 };
    assign _8088 = _7220[37:37];
    assign _8089 = { _8232,
                     _8088 };
    assign _8093 = _8089 + _8092;
    assign _8084 = _7220[38:38];
    assign _8085 = { _8232,
                     _8084 };
    assign _8081 = _7220[39:39];
    assign _8082 = { _8232,
                     _8081 };
    assign _8086 = _8082 + _8085;
    assign _8094 = _8086 + _8093;
    assign _8110 = _8094 + _8109;
    assign _8075 = _7220[40:40];
    assign _8076 = { _8232,
                     _8075 };
    assign _8072 = _7220[41:41];
    assign _8073 = { _8232,
                     _8072 };
    assign _8077 = _8073 + _8076;
    assign _8068 = _7220[42:42];
    assign _8069 = { _8232,
                     _8068 };
    assign _8065 = _7220[43:43];
    assign _8066 = { _8232,
                     _8065 };
    assign _8070 = _8066 + _8069;
    assign _8078 = _8070 + _8077;
    assign _8060 = _7220[44:44];
    assign _8061 = { _8232,
                     _8060 };
    assign _8057 = _7220[45:45];
    assign _8058 = { _8232,
                     _8057 };
    assign _8062 = _8058 + _8061;
    assign _8053 = _7220[46:46];
    assign _8054 = { _8232,
                     _8053 };
    assign _8050 = _7220[47:47];
    assign _8051 = { _8232,
                     _8050 };
    assign _8055 = _8051 + _8054;
    assign _8063 = _8055 + _8062;
    assign _8079 = _8063 + _8078;
    assign _8111 = _8079 + _8110;
    assign _8043 = _7220[48:48];
    assign _8044 = { _8232,
                     _8043 };
    assign _8040 = _7220[49:49];
    assign _8041 = { _8232,
                     _8040 };
    assign _8045 = _8041 + _8044;
    assign _8036 = _7220[50:50];
    assign _8037 = { _8232,
                     _8036 };
    assign _8033 = _7220[51:51];
    assign _8034 = { _8232,
                     _8033 };
    assign _8038 = _8034 + _8037;
    assign _8046 = _8038 + _8045;
    assign _8028 = _7220[52:52];
    assign _8029 = { _8232,
                     _8028 };
    assign _8025 = _7220[53:53];
    assign _8026 = { _8232,
                     _8025 };
    assign _8030 = _8026 + _8029;
    assign _8021 = _7220[54:54];
    assign _8022 = { _8232,
                     _8021 };
    assign _8018 = _7220[55:55];
    assign _8019 = { _8232,
                     _8018 };
    assign _8023 = _8019 + _8022;
    assign _8031 = _8023 + _8030;
    assign _8047 = _8031 + _8046;
    assign _8012 = _7220[56:56];
    assign _8013 = { _8232,
                     _8012 };
    assign _8009 = _7220[57:57];
    assign _8010 = { _8232,
                     _8009 };
    assign _8014 = _8010 + _8013;
    assign _8005 = _7220[58:58];
    assign _8006 = { _8232,
                     _8005 };
    assign _8002 = _7220[59:59];
    assign _8003 = { _8232,
                     _8002 };
    assign _8007 = _8003 + _8006;
    assign _8015 = _8007 + _8014;
    assign _7997 = _7220[60:60];
    assign _7998 = { _8232,
                     _7997 };
    assign _7994 = _7220[61:61];
    assign _7995 = { _8232,
                     _7994 };
    assign _7999 = _7995 + _7998;
    assign _7990 = _7220[62:62];
    assign _7991 = { _8232,
                     _7990 };
    assign _7987 = _7220[63:63];
    assign _7988 = { _8232,
                     _7987 };
    assign _7992 = _7988 + _7991;
    assign _8000 = _7992 + _7999;
    assign _8016 = _8000 + _8015;
    assign _8048 = _8016 + _8047;
    assign _8112 = _8048 + _8111;
    assign _8240 = _8112 + _8239;
    assign _7978 = _7220[64:64];
    assign _7979 = { _8232,
                     _7978 };
    assign _7975 = _7220[65:65];
    assign _7976 = { _8232,
                     _7975 };
    assign _7980 = _7976 + _7979;
    assign _7971 = _7220[66:66];
    assign _7972 = { _8232,
                     _7971 };
    assign _7968 = _7220[67:67];
    assign _7969 = { _8232,
                     _7968 };
    assign _7973 = _7969 + _7972;
    assign _7981 = _7973 + _7980;
    assign _7963 = _7220[68:68];
    assign _7964 = { _8232,
                     _7963 };
    assign _7960 = _7220[69:69];
    assign _7961 = { _8232,
                     _7960 };
    assign _7965 = _7961 + _7964;
    assign _7956 = _7220[70:70];
    assign _7957 = { _8232,
                     _7956 };
    assign _7953 = _7220[71:71];
    assign _7954 = { _8232,
                     _7953 };
    assign _7958 = _7954 + _7957;
    assign _7966 = _7958 + _7965;
    assign _7982 = _7966 + _7981;
    assign _7947 = _7220[72:72];
    assign _7948 = { _8232,
                     _7947 };
    assign _7944 = _7220[73:73];
    assign _7945 = { _8232,
                     _7944 };
    assign _7949 = _7945 + _7948;
    assign _7940 = _7220[74:74];
    assign _7941 = { _8232,
                     _7940 };
    assign _7937 = _7220[75:75];
    assign _7938 = { _8232,
                     _7937 };
    assign _7942 = _7938 + _7941;
    assign _7950 = _7942 + _7949;
    assign _7932 = _7220[76:76];
    assign _7933 = { _8232,
                     _7932 };
    assign _7929 = _7220[77:77];
    assign _7930 = { _8232,
                     _7929 };
    assign _7934 = _7930 + _7933;
    assign _7925 = _7220[78:78];
    assign _7926 = { _8232,
                     _7925 };
    assign _7922 = _7220[79:79];
    assign _7923 = { _8232,
                     _7922 };
    assign _7927 = _7923 + _7926;
    assign _7935 = _7927 + _7934;
    assign _7951 = _7935 + _7950;
    assign _7983 = _7951 + _7982;
    assign _7915 = _7220[80:80];
    assign _7916 = { _8232,
                     _7915 };
    assign _7912 = _7220[81:81];
    assign _7913 = { _8232,
                     _7912 };
    assign _7917 = _7913 + _7916;
    assign _7908 = _7220[82:82];
    assign _7909 = { _8232,
                     _7908 };
    assign _7905 = _7220[83:83];
    assign _7906 = { _8232,
                     _7905 };
    assign _7910 = _7906 + _7909;
    assign _7918 = _7910 + _7917;
    assign _7900 = _7220[84:84];
    assign _7901 = { _8232,
                     _7900 };
    assign _7897 = _7220[85:85];
    assign _7898 = { _8232,
                     _7897 };
    assign _7902 = _7898 + _7901;
    assign _7893 = _7220[86:86];
    assign _7894 = { _8232,
                     _7893 };
    assign _7890 = _7220[87:87];
    assign _7891 = { _8232,
                     _7890 };
    assign _7895 = _7891 + _7894;
    assign _7903 = _7895 + _7902;
    assign _7919 = _7903 + _7918;
    assign _7884 = _7220[88:88];
    assign _7885 = { _8232,
                     _7884 };
    assign _7881 = _7220[89:89];
    assign _7882 = { _8232,
                     _7881 };
    assign _7886 = _7882 + _7885;
    assign _7877 = _7220[90:90];
    assign _7878 = { _8232,
                     _7877 };
    assign _7874 = _7220[91:91];
    assign _7875 = { _8232,
                     _7874 };
    assign _7879 = _7875 + _7878;
    assign _7887 = _7879 + _7886;
    assign _7869 = _7220[92:92];
    assign _7870 = { _8232,
                     _7869 };
    assign _7866 = _7220[93:93];
    assign _7867 = { _8232,
                     _7866 };
    assign _7871 = _7867 + _7870;
    assign _7862 = _7220[94:94];
    assign _7863 = { _8232,
                     _7862 };
    assign _7859 = _7220[95:95];
    assign _7860 = { _8232,
                     _7859 };
    assign _7864 = _7860 + _7863;
    assign _7872 = _7864 + _7871;
    assign _7888 = _7872 + _7887;
    assign _7920 = _7888 + _7919;
    assign _7984 = _7920 + _7983;
    assign _7851 = _7220[96:96];
    assign _7852 = { _8232,
                     _7851 };
    assign _7848 = _7220[97:97];
    assign _7849 = { _8232,
                     _7848 };
    assign _7853 = _7849 + _7852;
    assign _7844 = _7220[98:98];
    assign _7845 = { _8232,
                     _7844 };
    assign _7841 = _7220[99:99];
    assign _7842 = { _8232,
                     _7841 };
    assign _7846 = _7842 + _7845;
    assign _7854 = _7846 + _7853;
    assign _7836 = _7220[100:100];
    assign _7837 = { _8232,
                     _7836 };
    assign _7833 = _7220[101:101];
    assign _7834 = { _8232,
                     _7833 };
    assign _7838 = _7834 + _7837;
    assign _7829 = _7220[102:102];
    assign _7830 = { _8232,
                     _7829 };
    assign _7826 = _7220[103:103];
    assign _7827 = { _8232,
                     _7826 };
    assign _7831 = _7827 + _7830;
    assign _7839 = _7831 + _7838;
    assign _7855 = _7839 + _7854;
    assign _7820 = _7220[104:104];
    assign _7821 = { _8232,
                     _7820 };
    assign _7817 = _7220[105:105];
    assign _7818 = { _8232,
                     _7817 };
    assign _7822 = _7818 + _7821;
    assign _7813 = _7220[106:106];
    assign _7814 = { _8232,
                     _7813 };
    assign _7810 = _7220[107:107];
    assign _7811 = { _8232,
                     _7810 };
    assign _7815 = _7811 + _7814;
    assign _7823 = _7815 + _7822;
    assign _7805 = _7220[108:108];
    assign _7806 = { _8232,
                     _7805 };
    assign _7802 = _7220[109:109];
    assign _7803 = { _8232,
                     _7802 };
    assign _7807 = _7803 + _7806;
    assign _7798 = _7220[110:110];
    assign _7799 = { _8232,
                     _7798 };
    assign _7795 = _7220[111:111];
    assign _7796 = { _8232,
                     _7795 };
    assign _7800 = _7796 + _7799;
    assign _7808 = _7800 + _7807;
    assign _7824 = _7808 + _7823;
    assign _7856 = _7824 + _7855;
    assign _7788 = _7220[112:112];
    assign _7789 = { _8232,
                     _7788 };
    assign _7785 = _7220[113:113];
    assign _7786 = { _8232,
                     _7785 };
    assign _7790 = _7786 + _7789;
    assign _7781 = _7220[114:114];
    assign _7782 = { _8232,
                     _7781 };
    assign _7778 = _7220[115:115];
    assign _7779 = { _8232,
                     _7778 };
    assign _7783 = _7779 + _7782;
    assign _7791 = _7783 + _7790;
    assign _7773 = _7220[116:116];
    assign _7774 = { _8232,
                     _7773 };
    assign _7770 = _7220[117:117];
    assign _7771 = { _8232,
                     _7770 };
    assign _7775 = _7771 + _7774;
    assign _7766 = _7220[118:118];
    assign _7767 = { _8232,
                     _7766 };
    assign _7763 = _7220[119:119];
    assign _7764 = { _8232,
                     _7763 };
    assign _7768 = _7764 + _7767;
    assign _7776 = _7768 + _7775;
    assign _7792 = _7776 + _7791;
    assign _7757 = _7220[120:120];
    assign _7758 = { _8232,
                     _7757 };
    assign _7754 = _7220[121:121];
    assign _7755 = { _8232,
                     _7754 };
    assign _7759 = _7755 + _7758;
    assign _7750 = _7220[122:122];
    assign _7751 = { _8232,
                     _7750 };
    assign _7747 = _7220[123:123];
    assign _7748 = { _8232,
                     _7747 };
    assign _7752 = _7748 + _7751;
    assign _7760 = _7752 + _7759;
    assign _7742 = _7220[124:124];
    assign _7743 = { _8232,
                     _7742 };
    assign _7739 = _7220[125:125];
    assign _7740 = { _8232,
                     _7739 };
    assign _7744 = _7740 + _7743;
    assign _7735 = _7220[126:126];
    assign _7736 = { _8232,
                     _7735 };
    assign _7732 = _7220[127:127];
    assign _7733 = { _8232,
                     _7732 };
    assign _7737 = _7733 + _7736;
    assign _7745 = _7737 + _7744;
    assign _7761 = _7745 + _7760;
    assign _7793 = _7761 + _7792;
    assign _7857 = _7793 + _7856;
    assign _7985 = _7857 + _7984;
    assign _8241 = _7985 + _8240;
    assign _7722 = _7220[128:128];
    assign _7723 = { _8232,
                     _7722 };
    assign _7719 = _7220[129:129];
    assign _7720 = { _8232,
                     _7719 };
    assign _7724 = _7720 + _7723;
    assign _7715 = _7220[130:130];
    assign _7716 = { _8232,
                     _7715 };
    assign _7712 = _7220[131:131];
    assign _7713 = { _8232,
                     _7712 };
    assign _7717 = _7713 + _7716;
    assign _7725 = _7717 + _7724;
    assign _7707 = _7220[132:132];
    assign _7708 = { _8232,
                     _7707 };
    assign _7704 = _7220[133:133];
    assign _7705 = { _8232,
                     _7704 };
    assign _7709 = _7705 + _7708;
    assign _7700 = _7220[134:134];
    assign _7701 = { _8232,
                     _7700 };
    assign _7697 = _7220[135:135];
    assign _7698 = { _8232,
                     _7697 };
    assign _7702 = _7698 + _7701;
    assign _7710 = _7702 + _7709;
    assign _7726 = _7710 + _7725;
    assign _7691 = _7220[136:136];
    assign _7692 = { _8232,
                     _7691 };
    assign _7688 = _7220[137:137];
    assign _7689 = { _8232,
                     _7688 };
    assign _7693 = _7689 + _7692;
    assign _7684 = _7220[138:138];
    assign _7685 = { _8232,
                     _7684 };
    assign _7681 = _7220[139:139];
    assign _7682 = { _8232,
                     _7681 };
    assign _7686 = _7682 + _7685;
    assign _7694 = _7686 + _7693;
    assign _7676 = _7220[140:140];
    assign _7677 = { _8232,
                     _7676 };
    assign _7673 = _7220[141:141];
    assign _7674 = { _8232,
                     _7673 };
    assign _7678 = _7674 + _7677;
    assign _7669 = _7220[142:142];
    assign _7670 = { _8232,
                     _7669 };
    assign _7666 = _7220[143:143];
    assign _7667 = { _8232,
                     _7666 };
    assign _7671 = _7667 + _7670;
    assign _7679 = _7671 + _7678;
    assign _7695 = _7679 + _7694;
    assign _7727 = _7695 + _7726;
    assign _7659 = _7220[144:144];
    assign _7660 = { _8232,
                     _7659 };
    assign _7656 = _7220[145:145];
    assign _7657 = { _8232,
                     _7656 };
    assign _7661 = _7657 + _7660;
    assign _7652 = _7220[146:146];
    assign _7653 = { _8232,
                     _7652 };
    assign _7649 = _7220[147:147];
    assign _7650 = { _8232,
                     _7649 };
    assign _7654 = _7650 + _7653;
    assign _7662 = _7654 + _7661;
    assign _7644 = _7220[148:148];
    assign _7645 = { _8232,
                     _7644 };
    assign _7641 = _7220[149:149];
    assign _7642 = { _8232,
                     _7641 };
    assign _7646 = _7642 + _7645;
    assign _7637 = _7220[150:150];
    assign _7638 = { _8232,
                     _7637 };
    assign _7634 = _7220[151:151];
    assign _7635 = { _8232,
                     _7634 };
    assign _7639 = _7635 + _7638;
    assign _7647 = _7639 + _7646;
    assign _7663 = _7647 + _7662;
    assign _7628 = _7220[152:152];
    assign _7629 = { _8232,
                     _7628 };
    assign _7625 = _7220[153:153];
    assign _7626 = { _8232,
                     _7625 };
    assign _7630 = _7626 + _7629;
    assign _7621 = _7220[154:154];
    assign _7622 = { _8232,
                     _7621 };
    assign _7618 = _7220[155:155];
    assign _7619 = { _8232,
                     _7618 };
    assign _7623 = _7619 + _7622;
    assign _7631 = _7623 + _7630;
    assign _7613 = _7220[156:156];
    assign _7614 = { _8232,
                     _7613 };
    assign _7610 = _7220[157:157];
    assign _7611 = { _8232,
                     _7610 };
    assign _7615 = _7611 + _7614;
    assign _7606 = _7220[158:158];
    assign _7607 = { _8232,
                     _7606 };
    assign _7603 = _7220[159:159];
    assign _7604 = { _8232,
                     _7603 };
    assign _7608 = _7604 + _7607;
    assign _7616 = _7608 + _7615;
    assign _7632 = _7616 + _7631;
    assign _7664 = _7632 + _7663;
    assign _7728 = _7664 + _7727;
    assign _7595 = _7220[160:160];
    assign _7596 = { _8232,
                     _7595 };
    assign _7592 = _7220[161:161];
    assign _7593 = { _8232,
                     _7592 };
    assign _7597 = _7593 + _7596;
    assign _7588 = _7220[162:162];
    assign _7589 = { _8232,
                     _7588 };
    assign _7585 = _7220[163:163];
    assign _7586 = { _8232,
                     _7585 };
    assign _7590 = _7586 + _7589;
    assign _7598 = _7590 + _7597;
    assign _7580 = _7220[164:164];
    assign _7581 = { _8232,
                     _7580 };
    assign _7577 = _7220[165:165];
    assign _7578 = { _8232,
                     _7577 };
    assign _7582 = _7578 + _7581;
    assign _7573 = _7220[166:166];
    assign _7574 = { _8232,
                     _7573 };
    assign _7570 = _7220[167:167];
    assign _7571 = { _8232,
                     _7570 };
    assign _7575 = _7571 + _7574;
    assign _7583 = _7575 + _7582;
    assign _7599 = _7583 + _7598;
    assign _7564 = _7220[168:168];
    assign _7565 = { _8232,
                     _7564 };
    assign _7561 = _7220[169:169];
    assign _7562 = { _8232,
                     _7561 };
    assign _7566 = _7562 + _7565;
    assign _7557 = _7220[170:170];
    assign _7558 = { _8232,
                     _7557 };
    assign _7554 = _7220[171:171];
    assign _7555 = { _8232,
                     _7554 };
    assign _7559 = _7555 + _7558;
    assign _7567 = _7559 + _7566;
    assign _7549 = _7220[172:172];
    assign _7550 = { _8232,
                     _7549 };
    assign _7546 = _7220[173:173];
    assign _7547 = { _8232,
                     _7546 };
    assign _7551 = _7547 + _7550;
    assign _7542 = _7220[174:174];
    assign _7543 = { _8232,
                     _7542 };
    assign _7539 = _7220[175:175];
    assign _7540 = { _8232,
                     _7539 };
    assign _7544 = _7540 + _7543;
    assign _7552 = _7544 + _7551;
    assign _7568 = _7552 + _7567;
    assign _7600 = _7568 + _7599;
    assign _7532 = _7220[176:176];
    assign _7533 = { _8232,
                     _7532 };
    assign _7529 = _7220[177:177];
    assign _7530 = { _8232,
                     _7529 };
    assign _7534 = _7530 + _7533;
    assign _7525 = _7220[178:178];
    assign _7526 = { _8232,
                     _7525 };
    assign _7522 = _7220[179:179];
    assign _7523 = { _8232,
                     _7522 };
    assign _7527 = _7523 + _7526;
    assign _7535 = _7527 + _7534;
    assign _7517 = _7220[180:180];
    assign _7518 = { _8232,
                     _7517 };
    assign _7514 = _7220[181:181];
    assign _7515 = { _8232,
                     _7514 };
    assign _7519 = _7515 + _7518;
    assign _7510 = _7220[182:182];
    assign _7511 = { _8232,
                     _7510 };
    assign _7507 = _7220[183:183];
    assign _7508 = { _8232,
                     _7507 };
    assign _7512 = _7508 + _7511;
    assign _7520 = _7512 + _7519;
    assign _7536 = _7520 + _7535;
    assign _7501 = _7220[184:184];
    assign _7502 = { _8232,
                     _7501 };
    assign _7498 = _7220[185:185];
    assign _7499 = { _8232,
                     _7498 };
    assign _7503 = _7499 + _7502;
    assign _7494 = _7220[186:186];
    assign _7495 = { _8232,
                     _7494 };
    assign _7491 = _7220[187:187];
    assign _7492 = { _8232,
                     _7491 };
    assign _7496 = _7492 + _7495;
    assign _7504 = _7496 + _7503;
    assign _7486 = _7220[188:188];
    assign _7487 = { _8232,
                     _7486 };
    assign _7483 = _7220[189:189];
    assign _7484 = { _8232,
                     _7483 };
    assign _7488 = _7484 + _7487;
    assign _7479 = _7220[190:190];
    assign _7480 = { _8232,
                     _7479 };
    assign _7476 = _7220[191:191];
    assign _7477 = { _8232,
                     _7476 };
    assign _7481 = _7477 + _7480;
    assign _7489 = _7481 + _7488;
    assign _7505 = _7489 + _7504;
    assign _7537 = _7505 + _7536;
    assign _7601 = _7537 + _7600;
    assign _7729 = _7601 + _7728;
    assign _7467 = _7220[192:192];
    assign _7468 = { _8232,
                     _7467 };
    assign _7464 = _7220[193:193];
    assign _7465 = { _8232,
                     _7464 };
    assign _7469 = _7465 + _7468;
    assign _7460 = _7220[194:194];
    assign _7461 = { _8232,
                     _7460 };
    assign _7457 = _7220[195:195];
    assign _7458 = { _8232,
                     _7457 };
    assign _7462 = _7458 + _7461;
    assign _7470 = _7462 + _7469;
    assign _7452 = _7220[196:196];
    assign _7453 = { _8232,
                     _7452 };
    assign _7449 = _7220[197:197];
    assign _7450 = { _8232,
                     _7449 };
    assign _7454 = _7450 + _7453;
    assign _7445 = _7220[198:198];
    assign _7446 = { _8232,
                     _7445 };
    assign _7442 = _7220[199:199];
    assign _7443 = { _8232,
                     _7442 };
    assign _7447 = _7443 + _7446;
    assign _7455 = _7447 + _7454;
    assign _7471 = _7455 + _7470;
    assign _7436 = _7220[200:200];
    assign _7437 = { _8232,
                     _7436 };
    assign _7433 = _7220[201:201];
    assign _7434 = { _8232,
                     _7433 };
    assign _7438 = _7434 + _7437;
    assign _7429 = _7220[202:202];
    assign _7430 = { _8232,
                     _7429 };
    assign _7426 = _7220[203:203];
    assign _7427 = { _8232,
                     _7426 };
    assign _7431 = _7427 + _7430;
    assign _7439 = _7431 + _7438;
    assign _7421 = _7220[204:204];
    assign _7422 = { _8232,
                     _7421 };
    assign _7418 = _7220[205:205];
    assign _7419 = { _8232,
                     _7418 };
    assign _7423 = _7419 + _7422;
    assign _7414 = _7220[206:206];
    assign _7415 = { _8232,
                     _7414 };
    assign _7411 = _7220[207:207];
    assign _7412 = { _8232,
                     _7411 };
    assign _7416 = _7412 + _7415;
    assign _7424 = _7416 + _7423;
    assign _7440 = _7424 + _7439;
    assign _7472 = _7440 + _7471;
    assign _7404 = _7220[208:208];
    assign _7405 = { _8232,
                     _7404 };
    assign _7401 = _7220[209:209];
    assign _7402 = { _8232,
                     _7401 };
    assign _7406 = _7402 + _7405;
    assign _7397 = _7220[210:210];
    assign _7398 = { _8232,
                     _7397 };
    assign _7394 = _7220[211:211];
    assign _7395 = { _8232,
                     _7394 };
    assign _7399 = _7395 + _7398;
    assign _7407 = _7399 + _7406;
    assign _7389 = _7220[212:212];
    assign _7390 = { _8232,
                     _7389 };
    assign _7386 = _7220[213:213];
    assign _7387 = { _8232,
                     _7386 };
    assign _7391 = _7387 + _7390;
    assign _7382 = _7220[214:214];
    assign _7383 = { _8232,
                     _7382 };
    assign _7379 = _7220[215:215];
    assign _7380 = { _8232,
                     _7379 };
    assign _7384 = _7380 + _7383;
    assign _7392 = _7384 + _7391;
    assign _7408 = _7392 + _7407;
    assign _7373 = _7220[216:216];
    assign _7374 = { _8232,
                     _7373 };
    assign _7370 = _7220[217:217];
    assign _7371 = { _8232,
                     _7370 };
    assign _7375 = _7371 + _7374;
    assign _7366 = _7220[218:218];
    assign _7367 = { _8232,
                     _7366 };
    assign _7363 = _7220[219:219];
    assign _7364 = { _8232,
                     _7363 };
    assign _7368 = _7364 + _7367;
    assign _7376 = _7368 + _7375;
    assign _7358 = _7220[220:220];
    assign _7359 = { _8232,
                     _7358 };
    assign _7355 = _7220[221:221];
    assign _7356 = { _8232,
                     _7355 };
    assign _7360 = _7356 + _7359;
    assign _7351 = _7220[222:222];
    assign _7352 = { _8232,
                     _7351 };
    assign _7348 = _7220[223:223];
    assign _7349 = { _8232,
                     _7348 };
    assign _7353 = _7349 + _7352;
    assign _7361 = _7353 + _7360;
    assign _7377 = _7361 + _7376;
    assign _7409 = _7377 + _7408;
    assign _7473 = _7409 + _7472;
    assign _7340 = _7220[224:224];
    assign _7341 = { _8232,
                     _7340 };
    assign _7337 = _7220[225:225];
    assign _7338 = { _8232,
                     _7337 };
    assign _7342 = _7338 + _7341;
    assign _7333 = _7220[226:226];
    assign _7334 = { _8232,
                     _7333 };
    assign _7330 = _7220[227:227];
    assign _7331 = { _8232,
                     _7330 };
    assign _7335 = _7331 + _7334;
    assign _7343 = _7335 + _7342;
    assign _7325 = _7220[228:228];
    assign _7326 = { _8232,
                     _7325 };
    assign _7322 = _7220[229:229];
    assign _7323 = { _8232,
                     _7322 };
    assign _7327 = _7323 + _7326;
    assign _7318 = _7220[230:230];
    assign _7319 = { _8232,
                     _7318 };
    assign _7315 = _7220[231:231];
    assign _7316 = { _8232,
                     _7315 };
    assign _7320 = _7316 + _7319;
    assign _7328 = _7320 + _7327;
    assign _7344 = _7328 + _7343;
    assign _7309 = _7220[232:232];
    assign _7310 = { _8232,
                     _7309 };
    assign _7306 = _7220[233:233];
    assign _7307 = { _8232,
                     _7306 };
    assign _7311 = _7307 + _7310;
    assign _7302 = _7220[234:234];
    assign _7303 = { _8232,
                     _7302 };
    assign _7299 = _7220[235:235];
    assign _7300 = { _8232,
                     _7299 };
    assign _7304 = _7300 + _7303;
    assign _7312 = _7304 + _7311;
    assign _7294 = _7220[236:236];
    assign _7295 = { _8232,
                     _7294 };
    assign _7291 = _7220[237:237];
    assign _7292 = { _8232,
                     _7291 };
    assign _7296 = _7292 + _7295;
    assign _7287 = _7220[238:238];
    assign _7288 = { _8232,
                     _7287 };
    assign _7284 = _7220[239:239];
    assign _7285 = { _8232,
                     _7284 };
    assign _7289 = _7285 + _7288;
    assign _7297 = _7289 + _7296;
    assign _7313 = _7297 + _7312;
    assign _7345 = _7313 + _7344;
    assign _7277 = _7220[240:240];
    assign _7278 = { _8232,
                     _7277 };
    assign _7274 = _7220[241:241];
    assign _7275 = { _8232,
                     _7274 };
    assign _7279 = _7275 + _7278;
    assign _7270 = _7220[242:242];
    assign _7271 = { _8232,
                     _7270 };
    assign _7267 = _7220[243:243];
    assign _7268 = { _8232,
                     _7267 };
    assign _7272 = _7268 + _7271;
    assign _7280 = _7272 + _7279;
    assign _7262 = _7220[244:244];
    assign _7263 = { _8232,
                     _7262 };
    assign _7259 = _7220[245:245];
    assign _7260 = { _8232,
                     _7259 };
    assign _7264 = _7260 + _7263;
    assign _7255 = _7220[246:246];
    assign _7256 = { _8232,
                     _7255 };
    assign _7252 = _7220[247:247];
    assign _7253 = { _8232,
                     _7252 };
    assign _7257 = _7253 + _7256;
    assign _7265 = _7257 + _7264;
    assign _7281 = _7265 + _7280;
    assign _7246 = _7220[248:248];
    assign _7247 = { _8232,
                     _7246 };
    assign _7243 = _7220[249:249];
    assign _7244 = { _8232,
                     _7243 };
    assign _7248 = _7244 + _7247;
    assign _7239 = _7220[250:250];
    assign _7240 = { _8232,
                     _7239 };
    assign _7236 = _7220[251:251];
    assign _7237 = { _8232,
                     _7236 };
    assign _7241 = _7237 + _7240;
    assign _7249 = _7241 + _7248;
    assign _7231 = _7220[252:252];
    assign _7232 = { _8232,
                     _7231 };
    assign _7228 = _7220[253:253];
    assign _7229 = { _8232,
                     _7228 };
    assign _7233 = _7229 + _7232;
    assign _7224 = _7220[254:254];
    assign _7225 = { _8232,
                     _7224 };
    assign _5396 = vdd ^ _303;
    assign _5397 = ~ _5396;
    assign _7212 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    assign _7209 = 8'b11111111;
    assign _7210 = _7 == _7209;
    assign _7213 = _7210 ? _7212 : _290;
    assign _5376 = gnd ^ _303;
    assign _5377 = ~ _5376;
    assign _7202 = 8'b11111110;
    assign _7203 = _7 == _7202;
    assign _7206 = _7203 ? _7212 : _290;
    assign _5400 = _5398 ? _5391 : _290;
    assign _5356 = vdd ^ _303;
    assign _5357 = ~ _5356;
    assign _7195 = 8'b11111101;
    assign _7196 = _7 == _7195;
    assign _7199 = _7196 ? _7212 : _290;
    assign _5380 = _5378 ? _5371 : _290;
    assign _5336 = gnd ^ _303;
    assign _5337 = ~ _5336;
    assign _7188 = 8'b11111100;
    assign _7189 = _7 == _7188;
    assign _7192 = _7189 ? _7212 : _290;
    assign _5360 = _5358 ? _5351 : _290;
    assign _5316 = vdd ^ _303;
    assign _5317 = ~ _5316;
    assign _7181 = 8'b11111011;
    assign _7182 = _7 == _7181;
    assign _7185 = _7182 ? _7212 : _290;
    assign _5340 = _5338 ? _5331 : _290;
    assign _5296 = gnd ^ _303;
    assign _5297 = ~ _5296;
    assign _7174 = 8'b11111010;
    assign _7175 = _7 == _7174;
    assign _7178 = _7175 ? _7212 : _290;
    assign _5320 = _5318 ? _5311 : _290;
    assign _5276 = vdd ^ _303;
    assign _5277 = ~ _5276;
    assign _7167 = 8'b11111001;
    assign _7168 = _7 == _7167;
    assign _7171 = _7168 ? _7212 : _290;
    assign _5300 = _5298 ? _5291 : _290;
    assign _5256 = gnd ^ _303;
    assign _5257 = ~ _5256;
    assign _7160 = 8'b11111000;
    assign _7161 = _7 == _7160;
    assign _7164 = _7161 ? _7212 : _290;
    assign _5280 = _5278 ? _5271 : _290;
    assign _5236 = vdd ^ _303;
    assign _5237 = ~ _5236;
    assign _7153 = 8'b11110111;
    assign _7154 = _7 == _7153;
    assign _7157 = _7154 ? _7212 : _290;
    assign _5260 = _5258 ? _5251 : _290;
    assign _5216 = gnd ^ _303;
    assign _5217 = ~ _5216;
    assign _7146 = 8'b11110110;
    assign _7147 = _7 == _7146;
    assign _7150 = _7147 ? _7212 : _290;
    assign _5240 = _5238 ? _5231 : _290;
    assign _5196 = vdd ^ _303;
    assign _5197 = ~ _5196;
    assign _7139 = 8'b11110101;
    assign _7140 = _7 == _7139;
    assign _7143 = _7140 ? _7212 : _290;
    assign _5220 = _5218 ? _5211 : _290;
    assign _5176 = gnd ^ _303;
    assign _5177 = ~ _5176;
    assign _7132 = 8'b11110100;
    assign _7133 = _7 == _7132;
    assign _7136 = _7133 ? _7212 : _290;
    assign _5200 = _5198 ? _5191 : _290;
    assign _5156 = vdd ^ _303;
    assign _5157 = ~ _5156;
    assign _7125 = 8'b11110011;
    assign _7126 = _7 == _7125;
    assign _7129 = _7126 ? _7212 : _290;
    assign _5180 = _5178 ? _5171 : _290;
    assign _5136 = gnd ^ _303;
    assign _5137 = ~ _5136;
    assign _7118 = 8'b11110010;
    assign _7119 = _7 == _7118;
    assign _7122 = _7119 ? _7212 : _290;
    assign _5160 = _5158 ? _5151 : _290;
    assign _5116 = vdd ^ _303;
    assign _5117 = ~ _5116;
    assign _7111 = 8'b11110001;
    assign _7112 = _7 == _7111;
    assign _7115 = _7112 ? _7212 : _290;
    assign _5140 = _5138 ? _5131 : _290;
    assign _5096 = gnd ^ _303;
    assign _5097 = ~ _5096;
    assign _7104 = 8'b11110000;
    assign _7105 = _7 == _7104;
    assign _7108 = _7105 ? _7212 : _290;
    assign _5120 = _5118 ? _5111 : _290;
    assign _5076 = vdd ^ _303;
    assign _5077 = ~ _5076;
    assign _7097 = 8'b11101111;
    assign _7098 = _7 == _7097;
    assign _7101 = _7098 ? _7212 : _290;
    assign _5100 = _5098 ? _5091 : _290;
    assign _5056 = gnd ^ _303;
    assign _5057 = ~ _5056;
    assign _7090 = 8'b11101110;
    assign _7091 = _7 == _7090;
    assign _7094 = _7091 ? _7212 : _290;
    assign _5080 = _5078 ? _5071 : _290;
    assign _5036 = vdd ^ _303;
    assign _5037 = ~ _5036;
    assign _7083 = 8'b11101101;
    assign _7084 = _7 == _7083;
    assign _7087 = _7084 ? _7212 : _290;
    assign _5060 = _5058 ? _5051 : _290;
    assign _5016 = gnd ^ _303;
    assign _5017 = ~ _5016;
    assign _7076 = 8'b11101100;
    assign _7077 = _7 == _7076;
    assign _7080 = _7077 ? _7212 : _290;
    assign _5040 = _5038 ? _5031 : _290;
    assign _4996 = vdd ^ _303;
    assign _4997 = ~ _4996;
    assign _7069 = 8'b11101011;
    assign _7070 = _7 == _7069;
    assign _7073 = _7070 ? _7212 : _290;
    assign _5020 = _5018 ? _5011 : _290;
    assign _4976 = gnd ^ _303;
    assign _4977 = ~ _4976;
    assign _7062 = 8'b11101010;
    assign _7063 = _7 == _7062;
    assign _7066 = _7063 ? _7212 : _290;
    assign _5000 = _4998 ? _4991 : _290;
    assign _4956 = vdd ^ _303;
    assign _4957 = ~ _4956;
    assign _7055 = 8'b11101001;
    assign _7056 = _7 == _7055;
    assign _7059 = _7056 ? _7212 : _290;
    assign _4980 = _4978 ? _4971 : _290;
    assign _4936 = gnd ^ _303;
    assign _4937 = ~ _4936;
    assign _7048 = 8'b11101000;
    assign _7049 = _7 == _7048;
    assign _7052 = _7049 ? _7212 : _290;
    assign _4960 = _4958 ? _4951 : _290;
    assign _4916 = vdd ^ _303;
    assign _4917 = ~ _4916;
    assign _7041 = 8'b11100111;
    assign _7042 = _7 == _7041;
    assign _7045 = _7042 ? _7212 : _290;
    assign _4940 = _4938 ? _4931 : _290;
    assign _4896 = gnd ^ _303;
    assign _4897 = ~ _4896;
    assign _7034 = 8'b11100110;
    assign _7035 = _7 == _7034;
    assign _7038 = _7035 ? _7212 : _290;
    assign _4920 = _4918 ? _4911 : _290;
    assign _4876 = vdd ^ _303;
    assign _4877 = ~ _4876;
    assign _7027 = 8'b11100101;
    assign _7028 = _7 == _7027;
    assign _7031 = _7028 ? _7212 : _290;
    assign _4900 = _4898 ? _4891 : _290;
    assign _4856 = gnd ^ _303;
    assign _4857 = ~ _4856;
    assign _7020 = 8'b11100100;
    assign _7021 = _7 == _7020;
    assign _7024 = _7021 ? _7212 : _290;
    assign _4880 = _4878 ? _4871 : _290;
    assign _4836 = vdd ^ _303;
    assign _4837 = ~ _4836;
    assign _7013 = 8'b11100011;
    assign _7014 = _7 == _7013;
    assign _7017 = _7014 ? _7212 : _290;
    assign _4860 = _4858 ? _4851 : _290;
    assign _4816 = gnd ^ _303;
    assign _4817 = ~ _4816;
    assign _7006 = 8'b11100010;
    assign _7007 = _7 == _7006;
    assign _7010 = _7007 ? _7212 : _290;
    assign _4840 = _4838 ? _4831 : _290;
    assign _4796 = vdd ^ _303;
    assign _4797 = ~ _4796;
    assign _6999 = 8'b11100001;
    assign _7000 = _7 == _6999;
    assign _7003 = _7000 ? _7212 : _290;
    assign _4820 = _4818 ? _4811 : _290;
    assign _4776 = gnd ^ _303;
    assign _4777 = ~ _4776;
    assign _6992 = 8'b11100000;
    assign _6993 = _7 == _6992;
    assign _6996 = _6993 ? _7212 : _290;
    assign _4800 = _4798 ? _4791 : _290;
    assign _4756 = vdd ^ _303;
    assign _4757 = ~ _4756;
    assign _6985 = 8'b11011111;
    assign _6986 = _7 == _6985;
    assign _6989 = _6986 ? _7212 : _290;
    assign _4780 = _4778 ? _4771 : _290;
    assign _4736 = gnd ^ _303;
    assign _4737 = ~ _4736;
    assign _6978 = 8'b11011110;
    assign _6979 = _7 == _6978;
    assign _6982 = _6979 ? _7212 : _290;
    assign _4760 = _4758 ? _4751 : _290;
    assign _4716 = vdd ^ _303;
    assign _4717 = ~ _4716;
    assign _6971 = 8'b11011101;
    assign _6972 = _7 == _6971;
    assign _6975 = _6972 ? _7212 : _290;
    assign _4740 = _4738 ? _4731 : _290;
    assign _4696 = gnd ^ _303;
    assign _4697 = ~ _4696;
    assign _6964 = 8'b11011100;
    assign _6965 = _7 == _6964;
    assign _6968 = _6965 ? _7212 : _290;
    assign _4720 = _4718 ? _4711 : _290;
    assign _4676 = vdd ^ _303;
    assign _4677 = ~ _4676;
    assign _6957 = 8'b11011011;
    assign _6958 = _7 == _6957;
    assign _6961 = _6958 ? _7212 : _290;
    assign _4700 = _4698 ? _4691 : _290;
    assign _4656 = gnd ^ _303;
    assign _4657 = ~ _4656;
    assign _6950 = 8'b11011010;
    assign _6951 = _7 == _6950;
    assign _6954 = _6951 ? _7212 : _290;
    assign _4680 = _4678 ? _4671 : _290;
    assign _4636 = vdd ^ _303;
    assign _4637 = ~ _4636;
    assign _6943 = 8'b11011001;
    assign _6944 = _7 == _6943;
    assign _6947 = _6944 ? _7212 : _290;
    assign _4660 = _4658 ? _4651 : _290;
    assign _4616 = gnd ^ _303;
    assign _4617 = ~ _4616;
    assign _6936 = 8'b11011000;
    assign _6937 = _7 == _6936;
    assign _6940 = _6937 ? _7212 : _290;
    assign _4640 = _4638 ? _4631 : _290;
    assign _4596 = vdd ^ _303;
    assign _4597 = ~ _4596;
    assign _6929 = 8'b11010111;
    assign _6930 = _7 == _6929;
    assign _6933 = _6930 ? _7212 : _290;
    assign _4620 = _4618 ? _4611 : _290;
    assign _4576 = gnd ^ _303;
    assign _4577 = ~ _4576;
    assign _6922 = 8'b11010110;
    assign _6923 = _7 == _6922;
    assign _6926 = _6923 ? _7212 : _290;
    assign _4600 = _4598 ? _4591 : _290;
    assign _4556 = vdd ^ _303;
    assign _4557 = ~ _4556;
    assign _6915 = 8'b11010101;
    assign _6916 = _7 == _6915;
    assign _6919 = _6916 ? _7212 : _290;
    assign _4580 = _4578 ? _4571 : _290;
    assign _4536 = gnd ^ _303;
    assign _4537 = ~ _4536;
    assign _6908 = 8'b11010100;
    assign _6909 = _7 == _6908;
    assign _6912 = _6909 ? _7212 : _290;
    assign _4560 = _4558 ? _4551 : _290;
    assign _4516 = vdd ^ _303;
    assign _4517 = ~ _4516;
    assign _6901 = 8'b11010011;
    assign _6902 = _7 == _6901;
    assign _6905 = _6902 ? _7212 : _290;
    assign _4540 = _4538 ? _4531 : _290;
    assign _4496 = gnd ^ _303;
    assign _4497 = ~ _4496;
    assign _6894 = 8'b11010010;
    assign _6895 = _7 == _6894;
    assign _6898 = _6895 ? _7212 : _290;
    assign _4520 = _4518 ? _4511 : _290;
    assign _4476 = vdd ^ _303;
    assign _4477 = ~ _4476;
    assign _6887 = 8'b11010001;
    assign _6888 = _7 == _6887;
    assign _6891 = _6888 ? _7212 : _290;
    assign _4500 = _4498 ? _4491 : _290;
    assign _4456 = gnd ^ _303;
    assign _4457 = ~ _4456;
    assign _6880 = 8'b11010000;
    assign _6881 = _7 == _6880;
    assign _6884 = _6881 ? _7212 : _290;
    assign _4480 = _4478 ? _4471 : _290;
    assign _4436 = vdd ^ _303;
    assign _4437 = ~ _4436;
    assign _6873 = 8'b11001111;
    assign _6874 = _7 == _6873;
    assign _6877 = _6874 ? _7212 : _290;
    assign _4460 = _4458 ? _4451 : _290;
    assign _4416 = gnd ^ _303;
    assign _4417 = ~ _4416;
    assign _6866 = 8'b11001110;
    assign _6867 = _7 == _6866;
    assign _6870 = _6867 ? _7212 : _290;
    assign _4440 = _4438 ? _4431 : _290;
    assign _4396 = vdd ^ _303;
    assign _4397 = ~ _4396;
    assign _6859 = 8'b11001101;
    assign _6860 = _7 == _6859;
    assign _6863 = _6860 ? _7212 : _290;
    assign _4420 = _4418 ? _4411 : _290;
    assign _4376 = gnd ^ _303;
    assign _4377 = ~ _4376;
    assign _6852 = 8'b11001100;
    assign _6853 = _7 == _6852;
    assign _6856 = _6853 ? _7212 : _290;
    assign _4400 = _4398 ? _4391 : _290;
    assign _4356 = vdd ^ _303;
    assign _4357 = ~ _4356;
    assign _6845 = 8'b11001011;
    assign _6846 = _7 == _6845;
    assign _6849 = _6846 ? _7212 : _290;
    assign _4380 = _4378 ? _4371 : _290;
    assign _4336 = gnd ^ _303;
    assign _4337 = ~ _4336;
    assign _6838 = 8'b11001010;
    assign _6839 = _7 == _6838;
    assign _6842 = _6839 ? _7212 : _290;
    assign _4360 = _4358 ? _4351 : _290;
    assign _4316 = vdd ^ _303;
    assign _4317 = ~ _4316;
    assign _6831 = 8'b11001001;
    assign _6832 = _7 == _6831;
    assign _6835 = _6832 ? _7212 : _290;
    assign _4340 = _4338 ? _4331 : _290;
    assign _4296 = gnd ^ _303;
    assign _4297 = ~ _4296;
    assign _6824 = 8'b11001000;
    assign _6825 = _7 == _6824;
    assign _6828 = _6825 ? _7212 : _290;
    assign _4320 = _4318 ? _4311 : _290;
    assign _4276 = vdd ^ _303;
    assign _4277 = ~ _4276;
    assign _6817 = 8'b11000111;
    assign _6818 = _7 == _6817;
    assign _6821 = _6818 ? _7212 : _290;
    assign _4300 = _4298 ? _4291 : _290;
    assign _4256 = gnd ^ _303;
    assign _4257 = ~ _4256;
    assign _6810 = 8'b11000110;
    assign _6811 = _7 == _6810;
    assign _6814 = _6811 ? _7212 : _290;
    assign _4280 = _4278 ? _4271 : _290;
    assign _4236 = vdd ^ _303;
    assign _4237 = ~ _4236;
    assign _6803 = 8'b11000101;
    assign _6804 = _7 == _6803;
    assign _6807 = _6804 ? _7212 : _290;
    assign _4260 = _4258 ? _4251 : _290;
    assign _4216 = gnd ^ _303;
    assign _4217 = ~ _4216;
    assign _6796 = 8'b11000100;
    assign _6797 = _7 == _6796;
    assign _6800 = _6797 ? _7212 : _290;
    assign _4240 = _4238 ? _4231 : _290;
    assign _4196 = vdd ^ _303;
    assign _4197 = ~ _4196;
    assign _6789 = 8'b11000011;
    assign _6790 = _7 == _6789;
    assign _6793 = _6790 ? _7212 : _290;
    assign _4220 = _4218 ? _4211 : _290;
    assign _4176 = gnd ^ _303;
    assign _4177 = ~ _4176;
    assign _6782 = 8'b11000010;
    assign _6783 = _7 == _6782;
    assign _6786 = _6783 ? _7212 : _290;
    assign _4200 = _4198 ? _4191 : _290;
    assign _4156 = vdd ^ _303;
    assign _4157 = ~ _4156;
    assign _6775 = 8'b11000001;
    assign _6776 = _7 == _6775;
    assign _6779 = _6776 ? _7212 : _290;
    assign _4180 = _4178 ? _4171 : _290;
    assign _4136 = gnd ^ _303;
    assign _4137 = ~ _4136;
    assign _6768 = 8'b11000000;
    assign _6769 = _7 == _6768;
    assign _6772 = _6769 ? _7212 : _290;
    assign _4160 = _4158 ? _4151 : _290;
    assign _4116 = vdd ^ _303;
    assign _4117 = ~ _4116;
    assign _6761 = 8'b10111111;
    assign _6762 = _7 == _6761;
    assign _6765 = _6762 ? _7212 : _290;
    assign _4140 = _4138 ? _4131 : _290;
    assign _4096 = gnd ^ _303;
    assign _4097 = ~ _4096;
    assign _6754 = 8'b10111110;
    assign _6755 = _7 == _6754;
    assign _6758 = _6755 ? _7212 : _290;
    assign _4120 = _4118 ? _4111 : _290;
    assign _4076 = vdd ^ _303;
    assign _4077 = ~ _4076;
    assign _6747 = 8'b10111101;
    assign _6748 = _7 == _6747;
    assign _6751 = _6748 ? _7212 : _290;
    assign _4100 = _4098 ? _4091 : _290;
    assign _4056 = gnd ^ _303;
    assign _4057 = ~ _4056;
    assign _6740 = 8'b10111100;
    assign _6741 = _7 == _6740;
    assign _6744 = _6741 ? _7212 : _290;
    assign _4080 = _4078 ? _4071 : _290;
    assign _4036 = vdd ^ _303;
    assign _4037 = ~ _4036;
    assign _6733 = 8'b10111011;
    assign _6734 = _7 == _6733;
    assign _6737 = _6734 ? _7212 : _290;
    assign _4060 = _4058 ? _4051 : _290;
    assign _4016 = gnd ^ _303;
    assign _4017 = ~ _4016;
    assign _6726 = 8'b10111010;
    assign _6727 = _7 == _6726;
    assign _6730 = _6727 ? _7212 : _290;
    assign _4040 = _4038 ? _4031 : _290;
    assign _3996 = vdd ^ _303;
    assign _3997 = ~ _3996;
    assign _6719 = 8'b10111001;
    assign _6720 = _7 == _6719;
    assign _6723 = _6720 ? _7212 : _290;
    assign _4020 = _4018 ? _4011 : _290;
    assign _3976 = gnd ^ _303;
    assign _3977 = ~ _3976;
    assign _6712 = 8'b10111000;
    assign _6713 = _7 == _6712;
    assign _6716 = _6713 ? _7212 : _290;
    assign _4000 = _3998 ? _3991 : _290;
    assign _3956 = vdd ^ _303;
    assign _3957 = ~ _3956;
    assign _6705 = 8'b10110111;
    assign _6706 = _7 == _6705;
    assign _6709 = _6706 ? _7212 : _290;
    assign _3980 = _3978 ? _3971 : _290;
    assign _3936 = gnd ^ _303;
    assign _3937 = ~ _3936;
    assign _6698 = 8'b10110110;
    assign _6699 = _7 == _6698;
    assign _6702 = _6699 ? _7212 : _290;
    assign _3960 = _3958 ? _3951 : _290;
    assign _3916 = vdd ^ _303;
    assign _3917 = ~ _3916;
    assign _6691 = 8'b10110101;
    assign _6692 = _7 == _6691;
    assign _6695 = _6692 ? _7212 : _290;
    assign _3940 = _3938 ? _3931 : _290;
    assign _3896 = gnd ^ _303;
    assign _3897 = ~ _3896;
    assign _6684 = 8'b10110100;
    assign _6685 = _7 == _6684;
    assign _6688 = _6685 ? _7212 : _290;
    assign _3920 = _3918 ? _3911 : _290;
    assign _3876 = vdd ^ _303;
    assign _3877 = ~ _3876;
    assign _6677 = 8'b10110011;
    assign _6678 = _7 == _6677;
    assign _6681 = _6678 ? _7212 : _290;
    assign _3900 = _3898 ? _3891 : _290;
    assign _3856 = gnd ^ _303;
    assign _3857 = ~ _3856;
    assign _6670 = 8'b10110010;
    assign _6671 = _7 == _6670;
    assign _6674 = _6671 ? _7212 : _290;
    assign _3880 = _3878 ? _3871 : _290;
    assign _3836 = vdd ^ _303;
    assign _3837 = ~ _3836;
    assign _6663 = 8'b10110001;
    assign _6664 = _7 == _6663;
    assign _6667 = _6664 ? _7212 : _290;
    assign _3860 = _3858 ? _3851 : _290;
    assign _3816 = gnd ^ _303;
    assign _3817 = ~ _3816;
    assign _6656 = 8'b10110000;
    assign _6657 = _7 == _6656;
    assign _6660 = _6657 ? _7212 : _290;
    assign _3840 = _3838 ? _3831 : _290;
    assign _3796 = vdd ^ _303;
    assign _3797 = ~ _3796;
    assign _6649 = 8'b10101111;
    assign _6650 = _7 == _6649;
    assign _6653 = _6650 ? _7212 : _290;
    assign _3820 = _3818 ? _3811 : _290;
    assign _3776 = gnd ^ _303;
    assign _3777 = ~ _3776;
    assign _6642 = 8'b10101110;
    assign _6643 = _7 == _6642;
    assign _6646 = _6643 ? _7212 : _290;
    assign _3800 = _3798 ? _3791 : _290;
    assign _3756 = vdd ^ _303;
    assign _3757 = ~ _3756;
    assign _6635 = 8'b10101101;
    assign _6636 = _7 == _6635;
    assign _6639 = _6636 ? _7212 : _290;
    assign _3780 = _3778 ? _3771 : _290;
    assign _3736 = gnd ^ _303;
    assign _3737 = ~ _3736;
    assign _6628 = 8'b10101100;
    assign _6629 = _7 == _6628;
    assign _6632 = _6629 ? _7212 : _290;
    assign _3760 = _3758 ? _3751 : _290;
    assign _3716 = vdd ^ _303;
    assign _3717 = ~ _3716;
    assign _6621 = 8'b10101011;
    assign _6622 = _7 == _6621;
    assign _6625 = _6622 ? _7212 : _290;
    assign _3740 = _3738 ? _3731 : _290;
    assign _3696 = gnd ^ _303;
    assign _3697 = ~ _3696;
    assign _6614 = 8'b10101010;
    assign _6615 = _7 == _6614;
    assign _6618 = _6615 ? _7212 : _290;
    assign _3720 = _3718 ? _3711 : _290;
    assign _3676 = vdd ^ _303;
    assign _3677 = ~ _3676;
    assign _6607 = 8'b10101001;
    assign _6608 = _7 == _6607;
    assign _6611 = _6608 ? _7212 : _290;
    assign _3700 = _3698 ? _3691 : _290;
    assign _3656 = gnd ^ _303;
    assign _3657 = ~ _3656;
    assign _6600 = 8'b10101000;
    assign _6601 = _7 == _6600;
    assign _6604 = _6601 ? _7212 : _290;
    assign _3680 = _3678 ? _3671 : _290;
    assign _3636 = vdd ^ _303;
    assign _3637 = ~ _3636;
    assign _6593 = 8'b10100111;
    assign _6594 = _7 == _6593;
    assign _6597 = _6594 ? _7212 : _290;
    assign _3660 = _3658 ? _3651 : _290;
    assign _3616 = gnd ^ _303;
    assign _3617 = ~ _3616;
    assign _6586 = 8'b10100110;
    assign _6587 = _7 == _6586;
    assign _6590 = _6587 ? _7212 : _290;
    assign _3640 = _3638 ? _3631 : _290;
    assign _3596 = vdd ^ _303;
    assign _3597 = ~ _3596;
    assign _6579 = 8'b10100101;
    assign _6580 = _7 == _6579;
    assign _6583 = _6580 ? _7212 : _290;
    assign _3620 = _3618 ? _3611 : _290;
    assign _3576 = gnd ^ _303;
    assign _3577 = ~ _3576;
    assign _6572 = 8'b10100100;
    assign _6573 = _7 == _6572;
    assign _6576 = _6573 ? _7212 : _290;
    assign _3600 = _3598 ? _3591 : _290;
    assign _3556 = vdd ^ _303;
    assign _3557 = ~ _3556;
    assign _6565 = 8'b10100011;
    assign _6566 = _7 == _6565;
    assign _6569 = _6566 ? _7212 : _290;
    assign _3580 = _3578 ? _3571 : _290;
    assign _3536 = gnd ^ _303;
    assign _3537 = ~ _3536;
    assign _6558 = 8'b10100010;
    assign _6559 = _7 == _6558;
    assign _6562 = _6559 ? _7212 : _290;
    assign _3560 = _3558 ? _3551 : _290;
    assign _3516 = vdd ^ _303;
    assign _3517 = ~ _3516;
    assign _6551 = 8'b10100001;
    assign _6552 = _7 == _6551;
    assign _6555 = _6552 ? _7212 : _290;
    assign _3540 = _3538 ? _3531 : _290;
    assign _3496 = gnd ^ _303;
    assign _3497 = ~ _3496;
    assign _6544 = 8'b10100000;
    assign _6545 = _7 == _6544;
    assign _6548 = _6545 ? _7212 : _290;
    assign _3520 = _3518 ? _3511 : _290;
    assign _3476 = vdd ^ _303;
    assign _3477 = ~ _3476;
    assign _6537 = 8'b10011111;
    assign _6538 = _7 == _6537;
    assign _6541 = _6538 ? _7212 : _290;
    assign _3500 = _3498 ? _3491 : _290;
    assign _3456 = gnd ^ _303;
    assign _3457 = ~ _3456;
    assign _6530 = 8'b10011110;
    assign _6531 = _7 == _6530;
    assign _6534 = _6531 ? _7212 : _290;
    assign _3480 = _3478 ? _3471 : _290;
    assign _3436 = vdd ^ _303;
    assign _3437 = ~ _3436;
    assign _6523 = 8'b10011101;
    assign _6524 = _7 == _6523;
    assign _6527 = _6524 ? _7212 : _290;
    assign _3460 = _3458 ? _3451 : _290;
    assign _3416 = gnd ^ _303;
    assign _3417 = ~ _3416;
    assign _6516 = 8'b10011100;
    assign _6517 = _7 == _6516;
    assign _6520 = _6517 ? _7212 : _290;
    assign _3440 = _3438 ? _3431 : _290;
    assign _3396 = vdd ^ _303;
    assign _3397 = ~ _3396;
    assign _6509 = 8'b10011011;
    assign _6510 = _7 == _6509;
    assign _6513 = _6510 ? _7212 : _290;
    assign _3420 = _3418 ? _3411 : _290;
    assign _3376 = gnd ^ _303;
    assign _3377 = ~ _3376;
    assign _6502 = 8'b10011010;
    assign _6503 = _7 == _6502;
    assign _6506 = _6503 ? _7212 : _290;
    assign _3400 = _3398 ? _3391 : _290;
    assign _3356 = vdd ^ _303;
    assign _3357 = ~ _3356;
    assign _6495 = 8'b10011001;
    assign _6496 = _7 == _6495;
    assign _6499 = _6496 ? _7212 : _290;
    assign _3380 = _3378 ? _3371 : _290;
    assign _3336 = gnd ^ _303;
    assign _3337 = ~ _3336;
    assign _6488 = 8'b10011000;
    assign _6489 = _7 == _6488;
    assign _6492 = _6489 ? _7212 : _290;
    assign _3360 = _3358 ? _3351 : _290;
    assign _3316 = vdd ^ _303;
    assign _3317 = ~ _3316;
    assign _6481 = 8'b10010111;
    assign _6482 = _7 == _6481;
    assign _6485 = _6482 ? _7212 : _290;
    assign _3340 = _3338 ? _3331 : _290;
    assign _3296 = gnd ^ _303;
    assign _3297 = ~ _3296;
    assign _6474 = 8'b10010110;
    assign _6475 = _7 == _6474;
    assign _6478 = _6475 ? _7212 : _290;
    assign _3320 = _3318 ? _3311 : _290;
    assign _3276 = vdd ^ _303;
    assign _3277 = ~ _3276;
    assign _6467 = 8'b10010101;
    assign _6468 = _7 == _6467;
    assign _6471 = _6468 ? _7212 : _290;
    assign _3300 = _3298 ? _3291 : _290;
    assign _3256 = gnd ^ _303;
    assign _3257 = ~ _3256;
    assign _6460 = 8'b10010100;
    assign _6461 = _7 == _6460;
    assign _6464 = _6461 ? _7212 : _290;
    assign _3280 = _3278 ? _3271 : _290;
    assign _3236 = vdd ^ _303;
    assign _3237 = ~ _3236;
    assign _6453 = 8'b10010011;
    assign _6454 = _7 == _6453;
    assign _6457 = _6454 ? _7212 : _290;
    assign _3260 = _3258 ? _3251 : _290;
    assign _3216 = gnd ^ _303;
    assign _3217 = ~ _3216;
    assign _6446 = 8'b10010010;
    assign _6447 = _7 == _6446;
    assign _6450 = _6447 ? _7212 : _290;
    assign _3240 = _3238 ? _3231 : _290;
    assign _3196 = vdd ^ _303;
    assign _3197 = ~ _3196;
    assign _6439 = 8'b10010001;
    assign _6440 = _7 == _6439;
    assign _6443 = _6440 ? _7212 : _290;
    assign _3220 = _3218 ? _3211 : _290;
    assign _3176 = gnd ^ _303;
    assign _3177 = ~ _3176;
    assign _6432 = 8'b10010000;
    assign _6433 = _7 == _6432;
    assign _6436 = _6433 ? _7212 : _290;
    assign _3200 = _3198 ? _3191 : _290;
    assign _3156 = vdd ^ _303;
    assign _3157 = ~ _3156;
    assign _6425 = 8'b10001111;
    assign _6426 = _7 == _6425;
    assign _6429 = _6426 ? _7212 : _290;
    assign _3180 = _3178 ? _3171 : _290;
    assign _3136 = gnd ^ _303;
    assign _3137 = ~ _3136;
    assign _6418 = 8'b10001110;
    assign _6419 = _7 == _6418;
    assign _6422 = _6419 ? _7212 : _290;
    assign _3160 = _3158 ? _3151 : _290;
    assign _3116 = vdd ^ _303;
    assign _3117 = ~ _3116;
    assign _6411 = 8'b10001101;
    assign _6412 = _7 == _6411;
    assign _6415 = _6412 ? _7212 : _290;
    assign _3140 = _3138 ? _3131 : _290;
    assign _3096 = gnd ^ _303;
    assign _3097 = ~ _3096;
    assign _6404 = 8'b10001100;
    assign _6405 = _7 == _6404;
    assign _6408 = _6405 ? _7212 : _290;
    assign _3120 = _3118 ? _3111 : _290;
    assign _3076 = vdd ^ _303;
    assign _3077 = ~ _3076;
    assign _6397 = 8'b10001011;
    assign _6398 = _7 == _6397;
    assign _6401 = _6398 ? _7212 : _290;
    assign _3100 = _3098 ? _3091 : _290;
    assign _3056 = gnd ^ _303;
    assign _3057 = ~ _3056;
    assign _6390 = 8'b10001010;
    assign _6391 = _7 == _6390;
    assign _6394 = _6391 ? _7212 : _290;
    assign _3080 = _3078 ? _3071 : _290;
    assign _3036 = vdd ^ _303;
    assign _3037 = ~ _3036;
    assign _6383 = 8'b10001001;
    assign _6384 = _7 == _6383;
    assign _6387 = _6384 ? _7212 : _290;
    assign _3060 = _3058 ? _3051 : _290;
    assign _3016 = gnd ^ _303;
    assign _3017 = ~ _3016;
    assign _6376 = 8'b10001000;
    assign _6377 = _7 == _6376;
    assign _6380 = _6377 ? _7212 : _290;
    assign _3040 = _3038 ? _3031 : _290;
    assign _2996 = vdd ^ _303;
    assign _2997 = ~ _2996;
    assign _6369 = 8'b10000111;
    assign _6370 = _7 == _6369;
    assign _6373 = _6370 ? _7212 : _290;
    assign _3020 = _3018 ? _3011 : _290;
    assign _2976 = gnd ^ _303;
    assign _2977 = ~ _2976;
    assign _6362 = 8'b10000110;
    assign _6363 = _7 == _6362;
    assign _6366 = _6363 ? _7212 : _290;
    assign _3000 = _2998 ? _2991 : _290;
    assign _2956 = vdd ^ _303;
    assign _2957 = ~ _2956;
    assign _6355 = 8'b10000101;
    assign _6356 = _7 == _6355;
    assign _6359 = _6356 ? _7212 : _290;
    assign _2980 = _2978 ? _2971 : _290;
    assign _2936 = gnd ^ _303;
    assign _2937 = ~ _2936;
    assign _6348 = 8'b10000100;
    assign _6349 = _7 == _6348;
    assign _6352 = _6349 ? _7212 : _290;
    assign _2960 = _2958 ? _2951 : _290;
    assign _2916 = vdd ^ _303;
    assign _2917 = ~ _2916;
    assign _6341 = 8'b10000011;
    assign _6342 = _7 == _6341;
    assign _6345 = _6342 ? _7212 : _290;
    assign _2940 = _2938 ? _2931 : _290;
    assign _2896 = gnd ^ _303;
    assign _2897 = ~ _2896;
    assign _6334 = 8'b10000010;
    assign _6335 = _7 == _6334;
    assign _6338 = _6335 ? _7212 : _290;
    assign _2920 = _2918 ? _2911 : _290;
    assign _2876 = vdd ^ _303;
    assign _2877 = ~ _2876;
    assign _6327 = 8'b10000001;
    assign _6328 = _7 == _6327;
    assign _6331 = _6328 ? _7212 : _290;
    assign _2900 = _2898 ? _2891 : _290;
    assign _2856 = gnd ^ _303;
    assign _2857 = ~ _2856;
    assign _6320 = 8'b10000000;
    assign _6321 = _7 == _6320;
    assign _6324 = _6321 ? _7212 : _290;
    assign _2880 = _2878 ? _2871 : _290;
    assign _2836 = vdd ^ _303;
    assign _2837 = ~ _2836;
    assign _6313 = 8'b01111111;
    assign _6314 = _7 == _6313;
    assign _6317 = _6314 ? _7212 : _290;
    assign _2860 = _2858 ? _2851 : _290;
    assign _2816 = gnd ^ _303;
    assign _2817 = ~ _2816;
    assign _6306 = 8'b01111110;
    assign _6307 = _7 == _6306;
    assign _6310 = _6307 ? _7212 : _290;
    assign _2840 = _2838 ? _2831 : _290;
    assign _2796 = vdd ^ _303;
    assign _2797 = ~ _2796;
    assign _6299 = 8'b01111101;
    assign _6300 = _7 == _6299;
    assign _6303 = _6300 ? _7212 : _290;
    assign _2820 = _2818 ? _2811 : _290;
    assign _2776 = gnd ^ _303;
    assign _2777 = ~ _2776;
    assign _6292 = 8'b01111100;
    assign _6293 = _7 == _6292;
    assign _6296 = _6293 ? _7212 : _290;
    assign _2800 = _2798 ? _2791 : _290;
    assign _2756 = vdd ^ _303;
    assign _2757 = ~ _2756;
    assign _6285 = 8'b01111011;
    assign _6286 = _7 == _6285;
    assign _6289 = _6286 ? _7212 : _290;
    assign _2780 = _2778 ? _2771 : _290;
    assign _2736 = gnd ^ _303;
    assign _2737 = ~ _2736;
    assign _6278 = 8'b01111010;
    assign _6279 = _7 == _6278;
    assign _6282 = _6279 ? _7212 : _290;
    assign _2760 = _2758 ? _2751 : _290;
    assign _2716 = vdd ^ _303;
    assign _2717 = ~ _2716;
    assign _6271 = 8'b01111001;
    assign _6272 = _7 == _6271;
    assign _6275 = _6272 ? _7212 : _290;
    assign _2740 = _2738 ? _2731 : _290;
    assign _2696 = gnd ^ _303;
    assign _2697 = ~ _2696;
    assign _6264 = 8'b01111000;
    assign _6265 = _7 == _6264;
    assign _6268 = _6265 ? _7212 : _290;
    assign _2720 = _2718 ? _2711 : _290;
    assign _2676 = vdd ^ _303;
    assign _2677 = ~ _2676;
    assign _6257 = 8'b01110111;
    assign _6258 = _7 == _6257;
    assign _6261 = _6258 ? _7212 : _290;
    assign _2700 = _2698 ? _2691 : _290;
    assign _2656 = gnd ^ _303;
    assign _2657 = ~ _2656;
    assign _6250 = 8'b01110110;
    assign _6251 = _7 == _6250;
    assign _6254 = _6251 ? _7212 : _290;
    assign _2680 = _2678 ? _2671 : _290;
    assign _2636 = vdd ^ _303;
    assign _2637 = ~ _2636;
    assign _6243 = 8'b01110101;
    assign _6244 = _7 == _6243;
    assign _6247 = _6244 ? _7212 : _290;
    assign _2660 = _2658 ? _2651 : _290;
    assign _2616 = gnd ^ _303;
    assign _2617 = ~ _2616;
    assign _6236 = 8'b01110100;
    assign _6237 = _7 == _6236;
    assign _6240 = _6237 ? _7212 : _290;
    assign _2640 = _2638 ? _2631 : _290;
    assign _2596 = vdd ^ _303;
    assign _2597 = ~ _2596;
    assign _6229 = 8'b01110011;
    assign _6230 = _7 == _6229;
    assign _6233 = _6230 ? _7212 : _290;
    assign _2620 = _2618 ? _2611 : _290;
    assign _2576 = gnd ^ _303;
    assign _2577 = ~ _2576;
    assign _6222 = 8'b01110010;
    assign _6223 = _7 == _6222;
    assign _6226 = _6223 ? _7212 : _290;
    assign _2600 = _2598 ? _2591 : _290;
    assign _2556 = vdd ^ _303;
    assign _2557 = ~ _2556;
    assign _6215 = 8'b01110001;
    assign _6216 = _7 == _6215;
    assign _6219 = _6216 ? _7212 : _290;
    assign _2580 = _2578 ? _2571 : _290;
    assign _2536 = gnd ^ _303;
    assign _2537 = ~ _2536;
    assign _6208 = 8'b01110000;
    assign _6209 = _7 == _6208;
    assign _6212 = _6209 ? _7212 : _290;
    assign _2560 = _2558 ? _2551 : _290;
    assign _2516 = vdd ^ _303;
    assign _2517 = ~ _2516;
    assign _6201 = 8'b01101111;
    assign _6202 = _7 == _6201;
    assign _6205 = _6202 ? _7212 : _290;
    assign _2540 = _2538 ? _2531 : _290;
    assign _2496 = gnd ^ _303;
    assign _2497 = ~ _2496;
    assign _6194 = 8'b01101110;
    assign _6195 = _7 == _6194;
    assign _6198 = _6195 ? _7212 : _290;
    assign _2520 = _2518 ? _2511 : _290;
    assign _2476 = vdd ^ _303;
    assign _2477 = ~ _2476;
    assign _6187 = 8'b01101101;
    assign _6188 = _7 == _6187;
    assign _6191 = _6188 ? _7212 : _290;
    assign _2500 = _2498 ? _2491 : _290;
    assign _2456 = gnd ^ _303;
    assign _2457 = ~ _2456;
    assign _6180 = 8'b01101100;
    assign _6181 = _7 == _6180;
    assign _6184 = _6181 ? _7212 : _290;
    assign _2480 = _2478 ? _2471 : _290;
    assign _2436 = vdd ^ _303;
    assign _2437 = ~ _2436;
    assign _6173 = 8'b01101011;
    assign _6174 = _7 == _6173;
    assign _6177 = _6174 ? _7212 : _290;
    assign _2460 = _2458 ? _2451 : _290;
    assign _2416 = gnd ^ _303;
    assign _2417 = ~ _2416;
    assign _6166 = 8'b01101010;
    assign _6167 = _7 == _6166;
    assign _6170 = _6167 ? _7212 : _290;
    assign _2440 = _2438 ? _2431 : _290;
    assign _2396 = vdd ^ _303;
    assign _2397 = ~ _2396;
    assign _6159 = 8'b01101001;
    assign _6160 = _7 == _6159;
    assign _6163 = _6160 ? _7212 : _290;
    assign _2420 = _2418 ? _2411 : _290;
    assign _2376 = gnd ^ _303;
    assign _2377 = ~ _2376;
    assign _6152 = 8'b01101000;
    assign _6153 = _7 == _6152;
    assign _6156 = _6153 ? _7212 : _290;
    assign _2400 = _2398 ? _2391 : _290;
    assign _2356 = vdd ^ _303;
    assign _2357 = ~ _2356;
    assign _6145 = 8'b01100111;
    assign _6146 = _7 == _6145;
    assign _6149 = _6146 ? _7212 : _290;
    assign _2380 = _2378 ? _2371 : _290;
    assign _2336 = gnd ^ _303;
    assign _2337 = ~ _2336;
    assign _6138 = 8'b01100110;
    assign _6139 = _7 == _6138;
    assign _6142 = _6139 ? _7212 : _290;
    assign _2360 = _2358 ? _2351 : _290;
    assign _2316 = vdd ^ _303;
    assign _2317 = ~ _2316;
    assign _6131 = 8'b01100101;
    assign _6132 = _7 == _6131;
    assign _6135 = _6132 ? _7212 : _290;
    assign _2340 = _2338 ? _2331 : _290;
    assign _2296 = gnd ^ _303;
    assign _2297 = ~ _2296;
    assign _6124 = 8'b01100100;
    assign _6125 = _7 == _6124;
    assign _6128 = _6125 ? _7212 : _290;
    assign _2320 = _2318 ? _2311 : _290;
    assign _2276 = vdd ^ _303;
    assign _2277 = ~ _2276;
    assign _6117 = 8'b01100011;
    assign _6118 = _7 == _6117;
    assign _6121 = _6118 ? _7212 : _290;
    assign _2300 = _2298 ? _2291 : _290;
    assign _2256 = gnd ^ _303;
    assign _2257 = ~ _2256;
    assign _6110 = 8'b01100010;
    assign _6111 = _7 == _6110;
    assign _6114 = _6111 ? _7212 : _290;
    assign _2280 = _2278 ? _2271 : _290;
    assign _2236 = vdd ^ _303;
    assign _2237 = ~ _2236;
    assign _6103 = 8'b01100001;
    assign _6104 = _7 == _6103;
    assign _6107 = _6104 ? _7212 : _290;
    assign _2260 = _2258 ? _2251 : _290;
    assign _2216 = gnd ^ _303;
    assign _2217 = ~ _2216;
    assign _6096 = 8'b01100000;
    assign _6097 = _7 == _6096;
    assign _6100 = _6097 ? _7212 : _290;
    assign _2240 = _2238 ? _2231 : _290;
    assign _2196 = vdd ^ _303;
    assign _2197 = ~ _2196;
    assign _6089 = 8'b01011111;
    assign _6090 = _7 == _6089;
    assign _6093 = _6090 ? _7212 : _290;
    assign _2220 = _2218 ? _2211 : _290;
    assign _2176 = gnd ^ _303;
    assign _2177 = ~ _2176;
    assign _6082 = 8'b01011110;
    assign _6083 = _7 == _6082;
    assign _6086 = _6083 ? _7212 : _290;
    assign _2200 = _2198 ? _2191 : _290;
    assign _2156 = vdd ^ _303;
    assign _2157 = ~ _2156;
    assign _6075 = 8'b01011101;
    assign _6076 = _7 == _6075;
    assign _6079 = _6076 ? _7212 : _290;
    assign _2180 = _2178 ? _2171 : _290;
    assign _2136 = gnd ^ _303;
    assign _2137 = ~ _2136;
    assign _6068 = 8'b01011100;
    assign _6069 = _7 == _6068;
    assign _6072 = _6069 ? _7212 : _290;
    assign _2160 = _2158 ? _2151 : _290;
    assign _2116 = vdd ^ _303;
    assign _2117 = ~ _2116;
    assign _6061 = 8'b01011011;
    assign _6062 = _7 == _6061;
    assign _6065 = _6062 ? _7212 : _290;
    assign _2140 = _2138 ? _2131 : _290;
    assign _2096 = gnd ^ _303;
    assign _2097 = ~ _2096;
    assign _6054 = 8'b01011010;
    assign _6055 = _7 == _6054;
    assign _6058 = _6055 ? _7212 : _290;
    assign _2120 = _2118 ? _2111 : _290;
    assign _2076 = vdd ^ _303;
    assign _2077 = ~ _2076;
    assign _6047 = 8'b01011001;
    assign _6048 = _7 == _6047;
    assign _6051 = _6048 ? _7212 : _290;
    assign _2100 = _2098 ? _2091 : _290;
    assign _2056 = gnd ^ _303;
    assign _2057 = ~ _2056;
    assign _6040 = 8'b01011000;
    assign _6041 = _7 == _6040;
    assign _6044 = _6041 ? _7212 : _290;
    assign _2080 = _2078 ? _2071 : _290;
    assign _2036 = vdd ^ _303;
    assign _2037 = ~ _2036;
    assign _6033 = 8'b01010111;
    assign _6034 = _7 == _6033;
    assign _6037 = _6034 ? _7212 : _290;
    assign _2060 = _2058 ? _2051 : _290;
    assign _2016 = gnd ^ _303;
    assign _2017 = ~ _2016;
    assign _6026 = 8'b01010110;
    assign _6027 = _7 == _6026;
    assign _6030 = _6027 ? _7212 : _290;
    assign _2040 = _2038 ? _2031 : _290;
    assign _1996 = vdd ^ _303;
    assign _1997 = ~ _1996;
    assign _6019 = 8'b01010101;
    assign _6020 = _7 == _6019;
    assign _6023 = _6020 ? _7212 : _290;
    assign _2020 = _2018 ? _2011 : _290;
    assign _1976 = gnd ^ _303;
    assign _1977 = ~ _1976;
    assign _6012 = 8'b01010100;
    assign _6013 = _7 == _6012;
    assign _6016 = _6013 ? _7212 : _290;
    assign _2000 = _1998 ? _1991 : _290;
    assign _1956 = vdd ^ _303;
    assign _1957 = ~ _1956;
    assign _6005 = 8'b01010011;
    assign _6006 = _7 == _6005;
    assign _6009 = _6006 ? _7212 : _290;
    assign _1980 = _1978 ? _1971 : _290;
    assign _1936 = gnd ^ _303;
    assign _1937 = ~ _1936;
    assign _5998 = 8'b01010010;
    assign _5999 = _7 == _5998;
    assign _6002 = _5999 ? _7212 : _290;
    assign _1960 = _1958 ? _1951 : _290;
    assign _1916 = vdd ^ _303;
    assign _1917 = ~ _1916;
    assign _5991 = 8'b01010001;
    assign _5992 = _7 == _5991;
    assign _5995 = _5992 ? _7212 : _290;
    assign _1940 = _1938 ? _1931 : _290;
    assign _1896 = gnd ^ _303;
    assign _1897 = ~ _1896;
    assign _5984 = 8'b01010000;
    assign _5985 = _7 == _5984;
    assign _5988 = _5985 ? _7212 : _290;
    assign _1920 = _1918 ? _1911 : _290;
    assign _1876 = vdd ^ _303;
    assign _1877 = ~ _1876;
    assign _5977 = 8'b01001111;
    assign _5978 = _7 == _5977;
    assign _5981 = _5978 ? _7212 : _290;
    assign _1900 = _1898 ? _1891 : _290;
    assign _1856 = gnd ^ _303;
    assign _1857 = ~ _1856;
    assign _5970 = 8'b01001110;
    assign _5971 = _7 == _5970;
    assign _5974 = _5971 ? _7212 : _290;
    assign _1880 = _1878 ? _1871 : _290;
    assign _1836 = vdd ^ _303;
    assign _1837 = ~ _1836;
    assign _5963 = 8'b01001101;
    assign _5964 = _7 == _5963;
    assign _5967 = _5964 ? _7212 : _290;
    assign _1860 = _1858 ? _1851 : _290;
    assign _1816 = gnd ^ _303;
    assign _1817 = ~ _1816;
    assign _5956 = 8'b01001100;
    assign _5957 = _7 == _5956;
    assign _5960 = _5957 ? _7212 : _290;
    assign _1840 = _1838 ? _1831 : _290;
    assign _1796 = vdd ^ _303;
    assign _1797 = ~ _1796;
    assign _5949 = 8'b01001011;
    assign _5950 = _7 == _5949;
    assign _5953 = _5950 ? _7212 : _290;
    assign _1820 = _1818 ? _1811 : _290;
    assign _1776 = gnd ^ _303;
    assign _1777 = ~ _1776;
    assign _5942 = 8'b01001010;
    assign _5943 = _7 == _5942;
    assign _5946 = _5943 ? _7212 : _290;
    assign _1800 = _1798 ? _1791 : _290;
    assign _1756 = vdd ^ _303;
    assign _1757 = ~ _1756;
    assign _5935 = 8'b01001001;
    assign _5936 = _7 == _5935;
    assign _5939 = _5936 ? _7212 : _290;
    assign _1780 = _1778 ? _1771 : _290;
    assign _1736 = gnd ^ _303;
    assign _1737 = ~ _1736;
    assign _5928 = 8'b01001000;
    assign _5929 = _7 == _5928;
    assign _5932 = _5929 ? _7212 : _290;
    assign _1760 = _1758 ? _1751 : _290;
    assign _1716 = vdd ^ _303;
    assign _1717 = ~ _1716;
    assign _5921 = 8'b01000111;
    assign _5922 = _7 == _5921;
    assign _5925 = _5922 ? _7212 : _290;
    assign _1740 = _1738 ? _1731 : _290;
    assign _1696 = gnd ^ _303;
    assign _1697 = ~ _1696;
    assign _5914 = 8'b01000110;
    assign _5915 = _7 == _5914;
    assign _5918 = _5915 ? _7212 : _290;
    assign _1720 = _1718 ? _1711 : _290;
    assign _1676 = vdd ^ _303;
    assign _1677 = ~ _1676;
    assign _5907 = 8'b01000101;
    assign _5908 = _7 == _5907;
    assign _5911 = _5908 ? _7212 : _290;
    assign _1700 = _1698 ? _1691 : _290;
    assign _1656 = gnd ^ _303;
    assign _1657 = ~ _1656;
    assign _5900 = 8'b01000100;
    assign _5901 = _7 == _5900;
    assign _5904 = _5901 ? _7212 : _290;
    assign _1680 = _1678 ? _1671 : _290;
    assign _1636 = vdd ^ _303;
    assign _1637 = ~ _1636;
    assign _5893 = 8'b01000011;
    assign _5894 = _7 == _5893;
    assign _5897 = _5894 ? _7212 : _290;
    assign _1660 = _1658 ? _1651 : _290;
    assign _1616 = gnd ^ _303;
    assign _1617 = ~ _1616;
    assign _5886 = 8'b01000010;
    assign _5887 = _7 == _5886;
    assign _5890 = _5887 ? _7212 : _290;
    assign _1640 = _1638 ? _1631 : _290;
    assign _1596 = vdd ^ _303;
    assign _1597 = ~ _1596;
    assign _5879 = 8'b01000001;
    assign _5880 = _7 == _5879;
    assign _5883 = _5880 ? _7212 : _290;
    assign _1620 = _1618 ? _1611 : _290;
    assign _1576 = gnd ^ _303;
    assign _1577 = ~ _1576;
    assign _5872 = 8'b01000000;
    assign _5873 = _7 == _5872;
    assign _5876 = _5873 ? _7212 : _290;
    assign _1600 = _1598 ? _1591 : _290;
    assign _1556 = vdd ^ _303;
    assign _1557 = ~ _1556;
    assign _5865 = 8'b00111111;
    assign _5866 = _7 == _5865;
    assign _5869 = _5866 ? _7212 : _290;
    assign _1580 = _1578 ? _1571 : _290;
    assign _1536 = gnd ^ _303;
    assign _1537 = ~ _1536;
    assign _5858 = 8'b00111110;
    assign _5859 = _7 == _5858;
    assign _5862 = _5859 ? _7212 : _290;
    assign _1560 = _1558 ? _1551 : _290;
    assign _1516 = vdd ^ _303;
    assign _1517 = ~ _1516;
    assign _5851 = 8'b00111101;
    assign _5852 = _7 == _5851;
    assign _5855 = _5852 ? _7212 : _290;
    assign _1540 = _1538 ? _1531 : _290;
    assign _1496 = gnd ^ _303;
    assign _1497 = ~ _1496;
    assign _5844 = 8'b00111100;
    assign _5845 = _7 == _5844;
    assign _5848 = _5845 ? _7212 : _290;
    assign _1520 = _1518 ? _1511 : _290;
    assign _1476 = vdd ^ _303;
    assign _1477 = ~ _1476;
    assign _5837 = 8'b00111011;
    assign _5838 = _7 == _5837;
    assign _5841 = _5838 ? _7212 : _290;
    assign _1500 = _1498 ? _1491 : _290;
    assign _1456 = gnd ^ _303;
    assign _1457 = ~ _1456;
    assign _5830 = 8'b00111010;
    assign _5831 = _7 == _5830;
    assign _5834 = _5831 ? _7212 : _290;
    assign _1480 = _1478 ? _1471 : _290;
    assign _1436 = vdd ^ _303;
    assign _1437 = ~ _1436;
    assign _5823 = 8'b00111001;
    assign _5824 = _7 == _5823;
    assign _5827 = _5824 ? _7212 : _290;
    assign _1460 = _1458 ? _1451 : _290;
    assign _1416 = gnd ^ _303;
    assign _1417 = ~ _1416;
    assign _5816 = 8'b00111000;
    assign _5817 = _7 == _5816;
    assign _5820 = _5817 ? _7212 : _290;
    assign _1440 = _1438 ? _1431 : _290;
    assign _1396 = vdd ^ _303;
    assign _1397 = ~ _1396;
    assign _5809 = 8'b00110111;
    assign _5810 = _7 == _5809;
    assign _5813 = _5810 ? _7212 : _290;
    assign _1420 = _1418 ? _1411 : _290;
    assign _1376 = gnd ^ _303;
    assign _1377 = ~ _1376;
    assign _5802 = 8'b00110110;
    assign _5803 = _7 == _5802;
    assign _5806 = _5803 ? _7212 : _290;
    assign _1400 = _1398 ? _1391 : _290;
    assign _1356 = vdd ^ _303;
    assign _1357 = ~ _1356;
    assign _5795 = 8'b00110101;
    assign _5796 = _7 == _5795;
    assign _5799 = _5796 ? _7212 : _290;
    assign _1380 = _1378 ? _1371 : _290;
    assign _1336 = gnd ^ _303;
    assign _1337 = ~ _1336;
    assign _5788 = 8'b00110100;
    assign _5789 = _7 == _5788;
    assign _5792 = _5789 ? _7212 : _290;
    assign _1360 = _1358 ? _1351 : _290;
    assign _1316 = vdd ^ _303;
    assign _1317 = ~ _1316;
    assign _5781 = 8'b00110011;
    assign _5782 = _7 == _5781;
    assign _5785 = _5782 ? _7212 : _290;
    assign _1340 = _1338 ? _1331 : _290;
    assign _1296 = gnd ^ _303;
    assign _1297 = ~ _1296;
    assign _5774 = 8'b00110010;
    assign _5775 = _7 == _5774;
    assign _5778 = _5775 ? _7212 : _290;
    assign _1320 = _1318 ? _1311 : _290;
    assign _1276 = vdd ^ _303;
    assign _1277 = ~ _1276;
    assign _5767 = 8'b00110001;
    assign _5768 = _7 == _5767;
    assign _5771 = _5768 ? _7212 : _290;
    assign _1300 = _1298 ? _1291 : _290;
    assign _1256 = gnd ^ _303;
    assign _1257 = ~ _1256;
    assign _5760 = 8'b00110000;
    assign _5761 = _7 == _5760;
    assign _5764 = _5761 ? _7212 : _290;
    assign _1280 = _1278 ? _1271 : _290;
    assign _1236 = vdd ^ _303;
    assign _1237 = ~ _1236;
    assign _5753 = 8'b00101111;
    assign _5754 = _7 == _5753;
    assign _5757 = _5754 ? _7212 : _290;
    assign _1260 = _1258 ? _1251 : _290;
    assign _1216 = gnd ^ _303;
    assign _1217 = ~ _1216;
    assign _5746 = 8'b00101110;
    assign _5747 = _7 == _5746;
    assign _5750 = _5747 ? _7212 : _290;
    assign _1240 = _1238 ? _1231 : _290;
    assign _1196 = vdd ^ _303;
    assign _1197 = ~ _1196;
    assign _5739 = 8'b00101101;
    assign _5740 = _7 == _5739;
    assign _5743 = _5740 ? _7212 : _290;
    assign _1220 = _1218 ? _1211 : _290;
    assign _1176 = gnd ^ _303;
    assign _1177 = ~ _1176;
    assign _5732 = 8'b00101100;
    assign _5733 = _7 == _5732;
    assign _5736 = _5733 ? _7212 : _290;
    assign _1200 = _1198 ? _1191 : _290;
    assign _1156 = vdd ^ _303;
    assign _1157 = ~ _1156;
    assign _5725 = 8'b00101011;
    assign _5726 = _7 == _5725;
    assign _5729 = _5726 ? _7212 : _290;
    assign _1180 = _1178 ? _1171 : _290;
    assign _1136 = gnd ^ _303;
    assign _1137 = ~ _1136;
    assign _5718 = 8'b00101010;
    assign _5719 = _7 == _5718;
    assign _5722 = _5719 ? _7212 : _290;
    assign _1160 = _1158 ? _1151 : _290;
    assign _1116 = vdd ^ _303;
    assign _1117 = ~ _1116;
    assign _5711 = 8'b00101001;
    assign _5712 = _7 == _5711;
    assign _5715 = _5712 ? _7212 : _290;
    assign _1140 = _1138 ? _1131 : _290;
    assign _1096 = gnd ^ _303;
    assign _1097 = ~ _1096;
    assign _5704 = 8'b00101000;
    assign _5705 = _7 == _5704;
    assign _5708 = _5705 ? _7212 : _290;
    assign _1120 = _1118 ? _1111 : _290;
    assign _1076 = vdd ^ _303;
    assign _1077 = ~ _1076;
    assign _5697 = 8'b00100111;
    assign _5698 = _7 == _5697;
    assign _5701 = _5698 ? _7212 : _290;
    assign _1100 = _1098 ? _1091 : _290;
    assign _1056 = gnd ^ _303;
    assign _1057 = ~ _1056;
    assign _5690 = 8'b00100110;
    assign _5691 = _7 == _5690;
    assign _5694 = _5691 ? _7212 : _290;
    assign _1080 = _1078 ? _1071 : _290;
    assign _1036 = vdd ^ _303;
    assign _1037 = ~ _1036;
    assign _5683 = 8'b00100101;
    assign _5684 = _7 == _5683;
    assign _5687 = _5684 ? _7212 : _290;
    assign _1060 = _1058 ? _1051 : _290;
    assign _1016 = gnd ^ _303;
    assign _1017 = ~ _1016;
    assign _5676 = 8'b00100100;
    assign _5677 = _7 == _5676;
    assign _5680 = _5677 ? _7212 : _290;
    assign _1040 = _1038 ? _1031 : _290;
    assign _996 = vdd ^ _303;
    assign _997 = ~ _996;
    assign _5669 = 8'b00100011;
    assign _5670 = _7 == _5669;
    assign _5673 = _5670 ? _7212 : _290;
    assign _1020 = _1018 ? _1011 : _290;
    assign _976 = gnd ^ _303;
    assign _977 = ~ _976;
    assign _5662 = 8'b00100010;
    assign _5663 = _7 == _5662;
    assign _5666 = _5663 ? _7212 : _290;
    assign _1000 = _998 ? _991 : _290;
    assign _956 = vdd ^ _303;
    assign _957 = ~ _956;
    assign _5655 = 8'b00100001;
    assign _5656 = _7 == _5655;
    assign _5659 = _5656 ? _7212 : _290;
    assign _980 = _978 ? _971 : _290;
    assign _936 = gnd ^ _303;
    assign _937 = ~ _936;
    assign _5648 = 8'b00100000;
    assign _5649 = _7 == _5648;
    assign _5652 = _5649 ? _7212 : _290;
    assign _960 = _958 ? _951 : _290;
    assign _916 = vdd ^ _303;
    assign _917 = ~ _916;
    assign _5641 = 8'b00011111;
    assign _5642 = _7 == _5641;
    assign _5645 = _5642 ? _7212 : _290;
    assign _940 = _938 ? _931 : _290;
    assign _896 = gnd ^ _303;
    assign _897 = ~ _896;
    assign _5634 = 8'b00011110;
    assign _5635 = _7 == _5634;
    assign _5638 = _5635 ? _7212 : _290;
    assign _920 = _918 ? _911 : _290;
    assign _876 = vdd ^ _303;
    assign _877 = ~ _876;
    assign _5627 = 8'b00011101;
    assign _5628 = _7 == _5627;
    assign _5631 = _5628 ? _7212 : _290;
    assign _900 = _898 ? _891 : _290;
    assign _856 = gnd ^ _303;
    assign _857 = ~ _856;
    assign _5620 = 8'b00011100;
    assign _5621 = _7 == _5620;
    assign _5624 = _5621 ? _7212 : _290;
    assign _880 = _878 ? _871 : _290;
    assign _836 = vdd ^ _303;
    assign _837 = ~ _836;
    assign _5613 = 8'b00011011;
    assign _5614 = _7 == _5613;
    assign _5617 = _5614 ? _7212 : _290;
    assign _860 = _858 ? _851 : _290;
    assign _816 = gnd ^ _303;
    assign _817 = ~ _816;
    assign _5606 = 8'b00011010;
    assign _5607 = _7 == _5606;
    assign _5610 = _5607 ? _7212 : _290;
    assign _840 = _838 ? _831 : _290;
    assign _796 = vdd ^ _303;
    assign _797 = ~ _796;
    assign _5599 = 8'b00011001;
    assign _5600 = _7 == _5599;
    assign _5603 = _5600 ? _7212 : _290;
    assign _820 = _818 ? _811 : _290;
    assign _776 = gnd ^ _303;
    assign _777 = ~ _776;
    assign _5592 = 8'b00011000;
    assign _5593 = _7 == _5592;
    assign _5596 = _5593 ? _7212 : _290;
    assign _800 = _798 ? _791 : _290;
    assign _756 = vdd ^ _303;
    assign _757 = ~ _756;
    assign _5585 = 8'b00010111;
    assign _5586 = _7 == _5585;
    assign _5589 = _5586 ? _7212 : _290;
    assign _780 = _778 ? _771 : _290;
    assign _736 = gnd ^ _303;
    assign _737 = ~ _736;
    assign _5578 = 8'b00010110;
    assign _5579 = _7 == _5578;
    assign _5582 = _5579 ? _7212 : _290;
    assign _760 = _758 ? _751 : _290;
    assign _716 = vdd ^ _303;
    assign _717 = ~ _716;
    assign _5571 = 8'b00010101;
    assign _5572 = _7 == _5571;
    assign _5575 = _5572 ? _7212 : _290;
    assign _740 = _738 ? _731 : _290;
    assign _696 = gnd ^ _303;
    assign _697 = ~ _696;
    assign _5564 = 8'b00010100;
    assign _5565 = _7 == _5564;
    assign _5568 = _5565 ? _7212 : _290;
    assign _720 = _718 ? _711 : _290;
    assign _676 = vdd ^ _303;
    assign _677 = ~ _676;
    assign _5557 = 8'b00010011;
    assign _5558 = _7 == _5557;
    assign _5561 = _5558 ? _7212 : _290;
    assign _700 = _698 ? _691 : _290;
    assign _656 = gnd ^ _303;
    assign _657 = ~ _656;
    assign _5550 = 8'b00010010;
    assign _5551 = _7 == _5550;
    assign _5554 = _5551 ? _7212 : _290;
    assign _680 = _678 ? _671 : _290;
    assign _636 = vdd ^ _303;
    assign _637 = ~ _636;
    assign _5543 = 8'b00010001;
    assign _5544 = _7 == _5543;
    assign _5547 = _5544 ? _7212 : _290;
    assign _660 = _658 ? _651 : _290;
    assign _616 = gnd ^ _303;
    assign _617 = ~ _616;
    assign _5536 = 8'b00010000;
    assign _5537 = _7 == _5536;
    assign _5540 = _5537 ? _7212 : _290;
    assign _640 = _638 ? _631 : _290;
    assign _596 = vdd ^ _303;
    assign _597 = ~ _596;
    assign _5529 = 8'b00001111;
    assign _5530 = _7 == _5529;
    assign _5533 = _5530 ? _7212 : _290;
    assign _620 = _618 ? _611 : _290;
    assign _576 = gnd ^ _303;
    assign _577 = ~ _576;
    assign _5522 = 8'b00001110;
    assign _5523 = _7 == _5522;
    assign _5526 = _5523 ? _7212 : _290;
    assign _600 = _598 ? _591 : _290;
    assign _556 = vdd ^ _303;
    assign _557 = ~ _556;
    assign _5515 = 8'b00001101;
    assign _5516 = _7 == _5515;
    assign _5519 = _5516 ? _7212 : _290;
    assign _580 = _578 ? _571 : _290;
    assign _536 = gnd ^ _303;
    assign _537 = ~ _536;
    assign _5508 = 8'b00001100;
    assign _5509 = _7 == _5508;
    assign _5512 = _5509 ? _7212 : _290;
    assign _560 = _558 ? _551 : _290;
    assign _516 = vdd ^ _303;
    assign _517 = ~ _516;
    assign _5501 = 8'b00001011;
    assign _5502 = _7 == _5501;
    assign _5505 = _5502 ? _7212 : _290;
    assign _540 = _538 ? _531 : _290;
    assign _496 = gnd ^ _303;
    assign _497 = ~ _496;
    assign _5494 = 8'b00001010;
    assign _5495 = _7 == _5494;
    assign _5498 = _5495 ? _7212 : _290;
    assign _520 = _518 ? _511 : _290;
    assign _476 = vdd ^ _303;
    assign _477 = ~ _476;
    assign _5487 = 8'b00001001;
    assign _5488 = _7 == _5487;
    assign _5491 = _5488 ? _7212 : _290;
    assign _500 = _498 ? _491 : _290;
    assign _456 = gnd ^ _303;
    assign _457 = ~ _456;
    assign _5480 = 8'b00001000;
    assign _5481 = _7 == _5480;
    assign _5484 = _5481 ? _7212 : _290;
    assign _480 = _478 ? _471 : _290;
    assign _436 = vdd ^ _303;
    assign _437 = ~ _436;
    assign _5473 = 8'b00000111;
    assign _5474 = _7 == _5473;
    assign _5477 = _5474 ? _7212 : _290;
    assign _460 = _458 ? _451 : _290;
    assign _416 = gnd ^ _303;
    assign _417 = ~ _416;
    assign _5466 = 8'b00000110;
    assign _5467 = _7 == _5466;
    assign _5470 = _5467 ? _7212 : _290;
    assign _440 = _438 ? _431 : _290;
    assign _396 = vdd ^ _303;
    assign _397 = ~ _396;
    assign _5459 = 8'b00000101;
    assign _5460 = _7 == _5459;
    assign _5463 = _5460 ? _7212 : _290;
    assign _420 = _418 ? _411 : _290;
    assign _376 = gnd ^ _303;
    assign _377 = ~ _376;
    assign _5452 = 8'b00000100;
    assign _5453 = _7 == _5452;
    assign _5456 = _5453 ? _7212 : _290;
    assign _400 = _398 ? _391 : _290;
    assign _356 = vdd ^ _303;
    assign _357 = ~ _356;
    assign _5445 = 8'b00000011;
    assign _5446 = _7 == _5445;
    assign _5449 = _5446 ? _7212 : _290;
    assign _380 = _378 ? _371 : _290;
    assign _336 = gnd ^ _303;
    assign _337 = ~ _336;
    assign _5438 = 8'b00000010;
    assign _5439 = _7 == _5438;
    assign _5442 = _5439 ? _7212 : _290;
    assign _360 = _358 ? _351 : _290;
    assign _317 = vdd ^ _303;
    assign _318 = ~ _317;
    assign _5431 = 8'b00000001;
    assign _5432 = _7 == _5431;
    assign _5435 = _5432 ? _7212 : _290;
    assign _340 = _338 ? _331 : _290;
    assign _302 = 1'b0;
    assign _5414 = _7[0:0];
    assign _5412 = ~ _303;
    assign _5413 = _287 ? _5412 : _303;
    assign _5415 = _278 ? _5414 : _5413;
    assign _4 = _5415;
    always @(posedge _272) begin
        if (_270)
            _303 <= _302;
        else
            _303 <= _4;
    end
    assign gnd = 1'b0;
    assign _304 = gnd ^ _303;
    assign _305 = ~ _304;
    assign _6 = width;
    assign _5420 = _6[7:1];
    assign _5421 = { _302,
                     _5420 };
    always @(posedge _272) begin
        if (_270)
            _5418 <= _8232;
        else
            _5418 <= _7;
    end
    assign _5422 = _278 ? _5421 : _5418;
    assign _7 = _5422;
    assign _5425 = _7 == _8232;
    assign _5428 = _5425 ? _7212 : _290;
    assign _321 = _319 ? _312 : _290;
    assign _308 = _306 ? _290 : _295;
    assign _322 = _308 + _321;
    assign _5423 = _287 ? _322 : _295;
    assign _5429 = _278 ? _5428 : _5423;
    assign _8 = _5429;
    always @(posedge _272) begin
        if (_270)
            _295 <= _290;
        else
            _295 <= _8;
    end
    assign _297 = _295 == _290;
    assign _298 = ~ _297;
    assign _292 = _265[0:0];
    assign _299 = _292 & _298;
    assign _306 = _299 & _305;
    assign _326 = _306 ? _295 : _290;
    assign _324 = _319 ? _290 : _312;
    assign _327 = _324 + _326;
    assign _341 = _327 + _340;
    assign _5430 = _287 ? _341 : _312;
    assign _5436 = _278 ? _5435 : _5430;
    assign _9 = _5436;
    always @(posedge _272) begin
        if (_270)
            _312 <= _290;
        else
            _312 <= _9;
    end
    assign _314 = _312 == _290;
    assign _315 = ~ _314;
    assign _309 = _265[1:1];
    assign _316 = _309 & _315;
    assign _319 = _316 & _318;
    assign _346 = _319 ? _312 : _290;
    assign _344 = _338 ? _290 : _331;
    assign _347 = _344 + _346;
    assign _361 = _347 + _360;
    assign _5437 = _287 ? _361 : _331;
    assign _5443 = _278 ? _5442 : _5437;
    assign _10 = _5443;
    always @(posedge _272) begin
        if (_270)
            _331 <= _290;
        else
            _331 <= _10;
    end
    assign _333 = _331 == _290;
    assign _334 = ~ _333;
    assign _328 = _265[2:2];
    assign _335 = _328 & _334;
    assign _338 = _335 & _337;
    assign _366 = _338 ? _331 : _290;
    assign _364 = _358 ? _290 : _351;
    assign _367 = _364 + _366;
    assign _381 = _367 + _380;
    assign _5444 = _287 ? _381 : _351;
    assign _5450 = _278 ? _5449 : _5444;
    assign _11 = _5450;
    always @(posedge _272) begin
        if (_270)
            _351 <= _290;
        else
            _351 <= _11;
    end
    assign _353 = _351 == _290;
    assign _354 = ~ _353;
    assign _348 = _265[3:3];
    assign _355 = _348 & _354;
    assign _358 = _355 & _357;
    assign _386 = _358 ? _351 : _290;
    assign _384 = _378 ? _290 : _371;
    assign _387 = _384 + _386;
    assign _401 = _387 + _400;
    assign _5451 = _287 ? _401 : _371;
    assign _5457 = _278 ? _5456 : _5451;
    assign _12 = _5457;
    always @(posedge _272) begin
        if (_270)
            _371 <= _290;
        else
            _371 <= _12;
    end
    assign _373 = _371 == _290;
    assign _374 = ~ _373;
    assign _368 = _265[4:4];
    assign _375 = _368 & _374;
    assign _378 = _375 & _377;
    assign _406 = _378 ? _371 : _290;
    assign _404 = _398 ? _290 : _391;
    assign _407 = _404 + _406;
    assign _421 = _407 + _420;
    assign _5458 = _287 ? _421 : _391;
    assign _5464 = _278 ? _5463 : _5458;
    assign _13 = _5464;
    always @(posedge _272) begin
        if (_270)
            _391 <= _290;
        else
            _391 <= _13;
    end
    assign _393 = _391 == _290;
    assign _394 = ~ _393;
    assign _388 = _265[5:5];
    assign _395 = _388 & _394;
    assign _398 = _395 & _397;
    assign _426 = _398 ? _391 : _290;
    assign _424 = _418 ? _290 : _411;
    assign _427 = _424 + _426;
    assign _441 = _427 + _440;
    assign _5465 = _287 ? _441 : _411;
    assign _5471 = _278 ? _5470 : _5465;
    assign _14 = _5471;
    always @(posedge _272) begin
        if (_270)
            _411 <= _290;
        else
            _411 <= _14;
    end
    assign _413 = _411 == _290;
    assign _414 = ~ _413;
    assign _408 = _265[6:6];
    assign _415 = _408 & _414;
    assign _418 = _415 & _417;
    assign _446 = _418 ? _411 : _290;
    assign _444 = _438 ? _290 : _431;
    assign _447 = _444 + _446;
    assign _461 = _447 + _460;
    assign _5472 = _287 ? _461 : _431;
    assign _5478 = _278 ? _5477 : _5472;
    assign _15 = _5478;
    always @(posedge _272) begin
        if (_270)
            _431 <= _290;
        else
            _431 <= _15;
    end
    assign _433 = _431 == _290;
    assign _434 = ~ _433;
    assign _428 = _265[7:7];
    assign _435 = _428 & _434;
    assign _438 = _435 & _437;
    assign _466 = _438 ? _431 : _290;
    assign _464 = _458 ? _290 : _451;
    assign _467 = _464 + _466;
    assign _481 = _467 + _480;
    assign _5479 = _287 ? _481 : _451;
    assign _5485 = _278 ? _5484 : _5479;
    assign _16 = _5485;
    always @(posedge _272) begin
        if (_270)
            _451 <= _290;
        else
            _451 <= _16;
    end
    assign _453 = _451 == _290;
    assign _454 = ~ _453;
    assign _448 = _265[8:8];
    assign _455 = _448 & _454;
    assign _458 = _455 & _457;
    assign _486 = _458 ? _451 : _290;
    assign _484 = _478 ? _290 : _471;
    assign _487 = _484 + _486;
    assign _501 = _487 + _500;
    assign _5486 = _287 ? _501 : _471;
    assign _5492 = _278 ? _5491 : _5486;
    assign _17 = _5492;
    always @(posedge _272) begin
        if (_270)
            _471 <= _290;
        else
            _471 <= _17;
    end
    assign _473 = _471 == _290;
    assign _474 = ~ _473;
    assign _468 = _265[9:9];
    assign _475 = _468 & _474;
    assign _478 = _475 & _477;
    assign _506 = _478 ? _471 : _290;
    assign _504 = _498 ? _290 : _491;
    assign _507 = _504 + _506;
    assign _521 = _507 + _520;
    assign _5493 = _287 ? _521 : _491;
    assign _5499 = _278 ? _5498 : _5493;
    assign _18 = _5499;
    always @(posedge _272) begin
        if (_270)
            _491 <= _290;
        else
            _491 <= _18;
    end
    assign _493 = _491 == _290;
    assign _494 = ~ _493;
    assign _488 = _265[10:10];
    assign _495 = _488 & _494;
    assign _498 = _495 & _497;
    assign _526 = _498 ? _491 : _290;
    assign _524 = _518 ? _290 : _511;
    assign _527 = _524 + _526;
    assign _541 = _527 + _540;
    assign _5500 = _287 ? _541 : _511;
    assign _5506 = _278 ? _5505 : _5500;
    assign _19 = _5506;
    always @(posedge _272) begin
        if (_270)
            _511 <= _290;
        else
            _511 <= _19;
    end
    assign _513 = _511 == _290;
    assign _514 = ~ _513;
    assign _508 = _265[11:11];
    assign _515 = _508 & _514;
    assign _518 = _515 & _517;
    assign _546 = _518 ? _511 : _290;
    assign _544 = _538 ? _290 : _531;
    assign _547 = _544 + _546;
    assign _561 = _547 + _560;
    assign _5507 = _287 ? _561 : _531;
    assign _5513 = _278 ? _5512 : _5507;
    assign _20 = _5513;
    always @(posedge _272) begin
        if (_270)
            _531 <= _290;
        else
            _531 <= _20;
    end
    assign _533 = _531 == _290;
    assign _534 = ~ _533;
    assign _528 = _265[12:12];
    assign _535 = _528 & _534;
    assign _538 = _535 & _537;
    assign _566 = _538 ? _531 : _290;
    assign _564 = _558 ? _290 : _551;
    assign _567 = _564 + _566;
    assign _581 = _567 + _580;
    assign _5514 = _287 ? _581 : _551;
    assign _5520 = _278 ? _5519 : _5514;
    assign _21 = _5520;
    always @(posedge _272) begin
        if (_270)
            _551 <= _290;
        else
            _551 <= _21;
    end
    assign _553 = _551 == _290;
    assign _554 = ~ _553;
    assign _548 = _265[13:13];
    assign _555 = _548 & _554;
    assign _558 = _555 & _557;
    assign _586 = _558 ? _551 : _290;
    assign _584 = _578 ? _290 : _571;
    assign _587 = _584 + _586;
    assign _601 = _587 + _600;
    assign _5521 = _287 ? _601 : _571;
    assign _5527 = _278 ? _5526 : _5521;
    assign _22 = _5527;
    always @(posedge _272) begin
        if (_270)
            _571 <= _290;
        else
            _571 <= _22;
    end
    assign _573 = _571 == _290;
    assign _574 = ~ _573;
    assign _568 = _265[14:14];
    assign _575 = _568 & _574;
    assign _578 = _575 & _577;
    assign _606 = _578 ? _571 : _290;
    assign _604 = _598 ? _290 : _591;
    assign _607 = _604 + _606;
    assign _621 = _607 + _620;
    assign _5528 = _287 ? _621 : _591;
    assign _5534 = _278 ? _5533 : _5528;
    assign _23 = _5534;
    always @(posedge _272) begin
        if (_270)
            _591 <= _290;
        else
            _591 <= _23;
    end
    assign _593 = _591 == _290;
    assign _594 = ~ _593;
    assign _588 = _265[15:15];
    assign _595 = _588 & _594;
    assign _598 = _595 & _597;
    assign _626 = _598 ? _591 : _290;
    assign _624 = _618 ? _290 : _611;
    assign _627 = _624 + _626;
    assign _641 = _627 + _640;
    assign _5535 = _287 ? _641 : _611;
    assign _5541 = _278 ? _5540 : _5535;
    assign _24 = _5541;
    always @(posedge _272) begin
        if (_270)
            _611 <= _290;
        else
            _611 <= _24;
    end
    assign _613 = _611 == _290;
    assign _614 = ~ _613;
    assign _608 = _265[16:16];
    assign _615 = _608 & _614;
    assign _618 = _615 & _617;
    assign _646 = _618 ? _611 : _290;
    assign _644 = _638 ? _290 : _631;
    assign _647 = _644 + _646;
    assign _661 = _647 + _660;
    assign _5542 = _287 ? _661 : _631;
    assign _5548 = _278 ? _5547 : _5542;
    assign _25 = _5548;
    always @(posedge _272) begin
        if (_270)
            _631 <= _290;
        else
            _631 <= _25;
    end
    assign _633 = _631 == _290;
    assign _634 = ~ _633;
    assign _628 = _265[17:17];
    assign _635 = _628 & _634;
    assign _638 = _635 & _637;
    assign _666 = _638 ? _631 : _290;
    assign _664 = _658 ? _290 : _651;
    assign _667 = _664 + _666;
    assign _681 = _667 + _680;
    assign _5549 = _287 ? _681 : _651;
    assign _5555 = _278 ? _5554 : _5549;
    assign _26 = _5555;
    always @(posedge _272) begin
        if (_270)
            _651 <= _290;
        else
            _651 <= _26;
    end
    assign _653 = _651 == _290;
    assign _654 = ~ _653;
    assign _648 = _265[18:18];
    assign _655 = _648 & _654;
    assign _658 = _655 & _657;
    assign _686 = _658 ? _651 : _290;
    assign _684 = _678 ? _290 : _671;
    assign _687 = _684 + _686;
    assign _701 = _687 + _700;
    assign _5556 = _287 ? _701 : _671;
    assign _5562 = _278 ? _5561 : _5556;
    assign _27 = _5562;
    always @(posedge _272) begin
        if (_270)
            _671 <= _290;
        else
            _671 <= _27;
    end
    assign _673 = _671 == _290;
    assign _674 = ~ _673;
    assign _668 = _265[19:19];
    assign _675 = _668 & _674;
    assign _678 = _675 & _677;
    assign _706 = _678 ? _671 : _290;
    assign _704 = _698 ? _290 : _691;
    assign _707 = _704 + _706;
    assign _721 = _707 + _720;
    assign _5563 = _287 ? _721 : _691;
    assign _5569 = _278 ? _5568 : _5563;
    assign _28 = _5569;
    always @(posedge _272) begin
        if (_270)
            _691 <= _290;
        else
            _691 <= _28;
    end
    assign _693 = _691 == _290;
    assign _694 = ~ _693;
    assign _688 = _265[20:20];
    assign _695 = _688 & _694;
    assign _698 = _695 & _697;
    assign _726 = _698 ? _691 : _290;
    assign _724 = _718 ? _290 : _711;
    assign _727 = _724 + _726;
    assign _741 = _727 + _740;
    assign _5570 = _287 ? _741 : _711;
    assign _5576 = _278 ? _5575 : _5570;
    assign _29 = _5576;
    always @(posedge _272) begin
        if (_270)
            _711 <= _290;
        else
            _711 <= _29;
    end
    assign _713 = _711 == _290;
    assign _714 = ~ _713;
    assign _708 = _265[21:21];
    assign _715 = _708 & _714;
    assign _718 = _715 & _717;
    assign _746 = _718 ? _711 : _290;
    assign _744 = _738 ? _290 : _731;
    assign _747 = _744 + _746;
    assign _761 = _747 + _760;
    assign _5577 = _287 ? _761 : _731;
    assign _5583 = _278 ? _5582 : _5577;
    assign _30 = _5583;
    always @(posedge _272) begin
        if (_270)
            _731 <= _290;
        else
            _731 <= _30;
    end
    assign _733 = _731 == _290;
    assign _734 = ~ _733;
    assign _728 = _265[22:22];
    assign _735 = _728 & _734;
    assign _738 = _735 & _737;
    assign _766 = _738 ? _731 : _290;
    assign _764 = _758 ? _290 : _751;
    assign _767 = _764 + _766;
    assign _781 = _767 + _780;
    assign _5584 = _287 ? _781 : _751;
    assign _5590 = _278 ? _5589 : _5584;
    assign _31 = _5590;
    always @(posedge _272) begin
        if (_270)
            _751 <= _290;
        else
            _751 <= _31;
    end
    assign _753 = _751 == _290;
    assign _754 = ~ _753;
    assign _748 = _265[23:23];
    assign _755 = _748 & _754;
    assign _758 = _755 & _757;
    assign _786 = _758 ? _751 : _290;
    assign _784 = _778 ? _290 : _771;
    assign _787 = _784 + _786;
    assign _801 = _787 + _800;
    assign _5591 = _287 ? _801 : _771;
    assign _5597 = _278 ? _5596 : _5591;
    assign _32 = _5597;
    always @(posedge _272) begin
        if (_270)
            _771 <= _290;
        else
            _771 <= _32;
    end
    assign _773 = _771 == _290;
    assign _774 = ~ _773;
    assign _768 = _265[24:24];
    assign _775 = _768 & _774;
    assign _778 = _775 & _777;
    assign _806 = _778 ? _771 : _290;
    assign _804 = _798 ? _290 : _791;
    assign _807 = _804 + _806;
    assign _821 = _807 + _820;
    assign _5598 = _287 ? _821 : _791;
    assign _5604 = _278 ? _5603 : _5598;
    assign _33 = _5604;
    always @(posedge _272) begin
        if (_270)
            _791 <= _290;
        else
            _791 <= _33;
    end
    assign _793 = _791 == _290;
    assign _794 = ~ _793;
    assign _788 = _265[25:25];
    assign _795 = _788 & _794;
    assign _798 = _795 & _797;
    assign _826 = _798 ? _791 : _290;
    assign _824 = _818 ? _290 : _811;
    assign _827 = _824 + _826;
    assign _841 = _827 + _840;
    assign _5605 = _287 ? _841 : _811;
    assign _5611 = _278 ? _5610 : _5605;
    assign _34 = _5611;
    always @(posedge _272) begin
        if (_270)
            _811 <= _290;
        else
            _811 <= _34;
    end
    assign _813 = _811 == _290;
    assign _814 = ~ _813;
    assign _808 = _265[26:26];
    assign _815 = _808 & _814;
    assign _818 = _815 & _817;
    assign _846 = _818 ? _811 : _290;
    assign _844 = _838 ? _290 : _831;
    assign _847 = _844 + _846;
    assign _861 = _847 + _860;
    assign _5612 = _287 ? _861 : _831;
    assign _5618 = _278 ? _5617 : _5612;
    assign _35 = _5618;
    always @(posedge _272) begin
        if (_270)
            _831 <= _290;
        else
            _831 <= _35;
    end
    assign _833 = _831 == _290;
    assign _834 = ~ _833;
    assign _828 = _265[27:27];
    assign _835 = _828 & _834;
    assign _838 = _835 & _837;
    assign _866 = _838 ? _831 : _290;
    assign _864 = _858 ? _290 : _851;
    assign _867 = _864 + _866;
    assign _881 = _867 + _880;
    assign _5619 = _287 ? _881 : _851;
    assign _5625 = _278 ? _5624 : _5619;
    assign _36 = _5625;
    always @(posedge _272) begin
        if (_270)
            _851 <= _290;
        else
            _851 <= _36;
    end
    assign _853 = _851 == _290;
    assign _854 = ~ _853;
    assign _848 = _265[28:28];
    assign _855 = _848 & _854;
    assign _858 = _855 & _857;
    assign _886 = _858 ? _851 : _290;
    assign _884 = _878 ? _290 : _871;
    assign _887 = _884 + _886;
    assign _901 = _887 + _900;
    assign _5626 = _287 ? _901 : _871;
    assign _5632 = _278 ? _5631 : _5626;
    assign _37 = _5632;
    always @(posedge _272) begin
        if (_270)
            _871 <= _290;
        else
            _871 <= _37;
    end
    assign _873 = _871 == _290;
    assign _874 = ~ _873;
    assign _868 = _265[29:29];
    assign _875 = _868 & _874;
    assign _878 = _875 & _877;
    assign _906 = _878 ? _871 : _290;
    assign _904 = _898 ? _290 : _891;
    assign _907 = _904 + _906;
    assign _921 = _907 + _920;
    assign _5633 = _287 ? _921 : _891;
    assign _5639 = _278 ? _5638 : _5633;
    assign _38 = _5639;
    always @(posedge _272) begin
        if (_270)
            _891 <= _290;
        else
            _891 <= _38;
    end
    assign _893 = _891 == _290;
    assign _894 = ~ _893;
    assign _888 = _265[30:30];
    assign _895 = _888 & _894;
    assign _898 = _895 & _897;
    assign _926 = _898 ? _891 : _290;
    assign _924 = _918 ? _290 : _911;
    assign _927 = _924 + _926;
    assign _941 = _927 + _940;
    assign _5640 = _287 ? _941 : _911;
    assign _5646 = _278 ? _5645 : _5640;
    assign _39 = _5646;
    always @(posedge _272) begin
        if (_270)
            _911 <= _290;
        else
            _911 <= _39;
    end
    assign _913 = _911 == _290;
    assign _914 = ~ _913;
    assign _908 = _265[31:31];
    assign _915 = _908 & _914;
    assign _918 = _915 & _917;
    assign _946 = _918 ? _911 : _290;
    assign _944 = _938 ? _290 : _931;
    assign _947 = _944 + _946;
    assign _961 = _947 + _960;
    assign _5647 = _287 ? _961 : _931;
    assign _5653 = _278 ? _5652 : _5647;
    assign _40 = _5653;
    always @(posedge _272) begin
        if (_270)
            _931 <= _290;
        else
            _931 <= _40;
    end
    assign _933 = _931 == _290;
    assign _934 = ~ _933;
    assign _928 = _265[32:32];
    assign _935 = _928 & _934;
    assign _938 = _935 & _937;
    assign _966 = _938 ? _931 : _290;
    assign _964 = _958 ? _290 : _951;
    assign _967 = _964 + _966;
    assign _981 = _967 + _980;
    assign _5654 = _287 ? _981 : _951;
    assign _5660 = _278 ? _5659 : _5654;
    assign _41 = _5660;
    always @(posedge _272) begin
        if (_270)
            _951 <= _290;
        else
            _951 <= _41;
    end
    assign _953 = _951 == _290;
    assign _954 = ~ _953;
    assign _948 = _265[33:33];
    assign _955 = _948 & _954;
    assign _958 = _955 & _957;
    assign _986 = _958 ? _951 : _290;
    assign _984 = _978 ? _290 : _971;
    assign _987 = _984 + _986;
    assign _1001 = _987 + _1000;
    assign _5661 = _287 ? _1001 : _971;
    assign _5667 = _278 ? _5666 : _5661;
    assign _42 = _5667;
    always @(posedge _272) begin
        if (_270)
            _971 <= _290;
        else
            _971 <= _42;
    end
    assign _973 = _971 == _290;
    assign _974 = ~ _973;
    assign _968 = _265[34:34];
    assign _975 = _968 & _974;
    assign _978 = _975 & _977;
    assign _1006 = _978 ? _971 : _290;
    assign _1004 = _998 ? _290 : _991;
    assign _1007 = _1004 + _1006;
    assign _1021 = _1007 + _1020;
    assign _5668 = _287 ? _1021 : _991;
    assign _5674 = _278 ? _5673 : _5668;
    assign _43 = _5674;
    always @(posedge _272) begin
        if (_270)
            _991 <= _290;
        else
            _991 <= _43;
    end
    assign _993 = _991 == _290;
    assign _994 = ~ _993;
    assign _988 = _265[35:35];
    assign _995 = _988 & _994;
    assign _998 = _995 & _997;
    assign _1026 = _998 ? _991 : _290;
    assign _1024 = _1018 ? _290 : _1011;
    assign _1027 = _1024 + _1026;
    assign _1041 = _1027 + _1040;
    assign _5675 = _287 ? _1041 : _1011;
    assign _5681 = _278 ? _5680 : _5675;
    assign _44 = _5681;
    always @(posedge _272) begin
        if (_270)
            _1011 <= _290;
        else
            _1011 <= _44;
    end
    assign _1013 = _1011 == _290;
    assign _1014 = ~ _1013;
    assign _1008 = _265[36:36];
    assign _1015 = _1008 & _1014;
    assign _1018 = _1015 & _1017;
    assign _1046 = _1018 ? _1011 : _290;
    assign _1044 = _1038 ? _290 : _1031;
    assign _1047 = _1044 + _1046;
    assign _1061 = _1047 + _1060;
    assign _5682 = _287 ? _1061 : _1031;
    assign _5688 = _278 ? _5687 : _5682;
    assign _45 = _5688;
    always @(posedge _272) begin
        if (_270)
            _1031 <= _290;
        else
            _1031 <= _45;
    end
    assign _1033 = _1031 == _290;
    assign _1034 = ~ _1033;
    assign _1028 = _265[37:37];
    assign _1035 = _1028 & _1034;
    assign _1038 = _1035 & _1037;
    assign _1066 = _1038 ? _1031 : _290;
    assign _1064 = _1058 ? _290 : _1051;
    assign _1067 = _1064 + _1066;
    assign _1081 = _1067 + _1080;
    assign _5689 = _287 ? _1081 : _1051;
    assign _5695 = _278 ? _5694 : _5689;
    assign _46 = _5695;
    always @(posedge _272) begin
        if (_270)
            _1051 <= _290;
        else
            _1051 <= _46;
    end
    assign _1053 = _1051 == _290;
    assign _1054 = ~ _1053;
    assign _1048 = _265[38:38];
    assign _1055 = _1048 & _1054;
    assign _1058 = _1055 & _1057;
    assign _1086 = _1058 ? _1051 : _290;
    assign _1084 = _1078 ? _290 : _1071;
    assign _1087 = _1084 + _1086;
    assign _1101 = _1087 + _1100;
    assign _5696 = _287 ? _1101 : _1071;
    assign _5702 = _278 ? _5701 : _5696;
    assign _47 = _5702;
    always @(posedge _272) begin
        if (_270)
            _1071 <= _290;
        else
            _1071 <= _47;
    end
    assign _1073 = _1071 == _290;
    assign _1074 = ~ _1073;
    assign _1068 = _265[39:39];
    assign _1075 = _1068 & _1074;
    assign _1078 = _1075 & _1077;
    assign _1106 = _1078 ? _1071 : _290;
    assign _1104 = _1098 ? _290 : _1091;
    assign _1107 = _1104 + _1106;
    assign _1121 = _1107 + _1120;
    assign _5703 = _287 ? _1121 : _1091;
    assign _5709 = _278 ? _5708 : _5703;
    assign _48 = _5709;
    always @(posedge _272) begin
        if (_270)
            _1091 <= _290;
        else
            _1091 <= _48;
    end
    assign _1093 = _1091 == _290;
    assign _1094 = ~ _1093;
    assign _1088 = _265[40:40];
    assign _1095 = _1088 & _1094;
    assign _1098 = _1095 & _1097;
    assign _1126 = _1098 ? _1091 : _290;
    assign _1124 = _1118 ? _290 : _1111;
    assign _1127 = _1124 + _1126;
    assign _1141 = _1127 + _1140;
    assign _5710 = _287 ? _1141 : _1111;
    assign _5716 = _278 ? _5715 : _5710;
    assign _49 = _5716;
    always @(posedge _272) begin
        if (_270)
            _1111 <= _290;
        else
            _1111 <= _49;
    end
    assign _1113 = _1111 == _290;
    assign _1114 = ~ _1113;
    assign _1108 = _265[41:41];
    assign _1115 = _1108 & _1114;
    assign _1118 = _1115 & _1117;
    assign _1146 = _1118 ? _1111 : _290;
    assign _1144 = _1138 ? _290 : _1131;
    assign _1147 = _1144 + _1146;
    assign _1161 = _1147 + _1160;
    assign _5717 = _287 ? _1161 : _1131;
    assign _5723 = _278 ? _5722 : _5717;
    assign _50 = _5723;
    always @(posedge _272) begin
        if (_270)
            _1131 <= _290;
        else
            _1131 <= _50;
    end
    assign _1133 = _1131 == _290;
    assign _1134 = ~ _1133;
    assign _1128 = _265[42:42];
    assign _1135 = _1128 & _1134;
    assign _1138 = _1135 & _1137;
    assign _1166 = _1138 ? _1131 : _290;
    assign _1164 = _1158 ? _290 : _1151;
    assign _1167 = _1164 + _1166;
    assign _1181 = _1167 + _1180;
    assign _5724 = _287 ? _1181 : _1151;
    assign _5730 = _278 ? _5729 : _5724;
    assign _51 = _5730;
    always @(posedge _272) begin
        if (_270)
            _1151 <= _290;
        else
            _1151 <= _51;
    end
    assign _1153 = _1151 == _290;
    assign _1154 = ~ _1153;
    assign _1148 = _265[43:43];
    assign _1155 = _1148 & _1154;
    assign _1158 = _1155 & _1157;
    assign _1186 = _1158 ? _1151 : _290;
    assign _1184 = _1178 ? _290 : _1171;
    assign _1187 = _1184 + _1186;
    assign _1201 = _1187 + _1200;
    assign _5731 = _287 ? _1201 : _1171;
    assign _5737 = _278 ? _5736 : _5731;
    assign _52 = _5737;
    always @(posedge _272) begin
        if (_270)
            _1171 <= _290;
        else
            _1171 <= _52;
    end
    assign _1173 = _1171 == _290;
    assign _1174 = ~ _1173;
    assign _1168 = _265[44:44];
    assign _1175 = _1168 & _1174;
    assign _1178 = _1175 & _1177;
    assign _1206 = _1178 ? _1171 : _290;
    assign _1204 = _1198 ? _290 : _1191;
    assign _1207 = _1204 + _1206;
    assign _1221 = _1207 + _1220;
    assign _5738 = _287 ? _1221 : _1191;
    assign _5744 = _278 ? _5743 : _5738;
    assign _53 = _5744;
    always @(posedge _272) begin
        if (_270)
            _1191 <= _290;
        else
            _1191 <= _53;
    end
    assign _1193 = _1191 == _290;
    assign _1194 = ~ _1193;
    assign _1188 = _265[45:45];
    assign _1195 = _1188 & _1194;
    assign _1198 = _1195 & _1197;
    assign _1226 = _1198 ? _1191 : _290;
    assign _1224 = _1218 ? _290 : _1211;
    assign _1227 = _1224 + _1226;
    assign _1241 = _1227 + _1240;
    assign _5745 = _287 ? _1241 : _1211;
    assign _5751 = _278 ? _5750 : _5745;
    assign _54 = _5751;
    always @(posedge _272) begin
        if (_270)
            _1211 <= _290;
        else
            _1211 <= _54;
    end
    assign _1213 = _1211 == _290;
    assign _1214 = ~ _1213;
    assign _1208 = _265[46:46];
    assign _1215 = _1208 & _1214;
    assign _1218 = _1215 & _1217;
    assign _1246 = _1218 ? _1211 : _290;
    assign _1244 = _1238 ? _290 : _1231;
    assign _1247 = _1244 + _1246;
    assign _1261 = _1247 + _1260;
    assign _5752 = _287 ? _1261 : _1231;
    assign _5758 = _278 ? _5757 : _5752;
    assign _55 = _5758;
    always @(posedge _272) begin
        if (_270)
            _1231 <= _290;
        else
            _1231 <= _55;
    end
    assign _1233 = _1231 == _290;
    assign _1234 = ~ _1233;
    assign _1228 = _265[47:47];
    assign _1235 = _1228 & _1234;
    assign _1238 = _1235 & _1237;
    assign _1266 = _1238 ? _1231 : _290;
    assign _1264 = _1258 ? _290 : _1251;
    assign _1267 = _1264 + _1266;
    assign _1281 = _1267 + _1280;
    assign _5759 = _287 ? _1281 : _1251;
    assign _5765 = _278 ? _5764 : _5759;
    assign _56 = _5765;
    always @(posedge _272) begin
        if (_270)
            _1251 <= _290;
        else
            _1251 <= _56;
    end
    assign _1253 = _1251 == _290;
    assign _1254 = ~ _1253;
    assign _1248 = _265[48:48];
    assign _1255 = _1248 & _1254;
    assign _1258 = _1255 & _1257;
    assign _1286 = _1258 ? _1251 : _290;
    assign _1284 = _1278 ? _290 : _1271;
    assign _1287 = _1284 + _1286;
    assign _1301 = _1287 + _1300;
    assign _5766 = _287 ? _1301 : _1271;
    assign _5772 = _278 ? _5771 : _5766;
    assign _57 = _5772;
    always @(posedge _272) begin
        if (_270)
            _1271 <= _290;
        else
            _1271 <= _57;
    end
    assign _1273 = _1271 == _290;
    assign _1274 = ~ _1273;
    assign _1268 = _265[49:49];
    assign _1275 = _1268 & _1274;
    assign _1278 = _1275 & _1277;
    assign _1306 = _1278 ? _1271 : _290;
    assign _1304 = _1298 ? _290 : _1291;
    assign _1307 = _1304 + _1306;
    assign _1321 = _1307 + _1320;
    assign _5773 = _287 ? _1321 : _1291;
    assign _5779 = _278 ? _5778 : _5773;
    assign _58 = _5779;
    always @(posedge _272) begin
        if (_270)
            _1291 <= _290;
        else
            _1291 <= _58;
    end
    assign _1293 = _1291 == _290;
    assign _1294 = ~ _1293;
    assign _1288 = _265[50:50];
    assign _1295 = _1288 & _1294;
    assign _1298 = _1295 & _1297;
    assign _1326 = _1298 ? _1291 : _290;
    assign _1324 = _1318 ? _290 : _1311;
    assign _1327 = _1324 + _1326;
    assign _1341 = _1327 + _1340;
    assign _5780 = _287 ? _1341 : _1311;
    assign _5786 = _278 ? _5785 : _5780;
    assign _59 = _5786;
    always @(posedge _272) begin
        if (_270)
            _1311 <= _290;
        else
            _1311 <= _59;
    end
    assign _1313 = _1311 == _290;
    assign _1314 = ~ _1313;
    assign _1308 = _265[51:51];
    assign _1315 = _1308 & _1314;
    assign _1318 = _1315 & _1317;
    assign _1346 = _1318 ? _1311 : _290;
    assign _1344 = _1338 ? _290 : _1331;
    assign _1347 = _1344 + _1346;
    assign _1361 = _1347 + _1360;
    assign _5787 = _287 ? _1361 : _1331;
    assign _5793 = _278 ? _5792 : _5787;
    assign _60 = _5793;
    always @(posedge _272) begin
        if (_270)
            _1331 <= _290;
        else
            _1331 <= _60;
    end
    assign _1333 = _1331 == _290;
    assign _1334 = ~ _1333;
    assign _1328 = _265[52:52];
    assign _1335 = _1328 & _1334;
    assign _1338 = _1335 & _1337;
    assign _1366 = _1338 ? _1331 : _290;
    assign _1364 = _1358 ? _290 : _1351;
    assign _1367 = _1364 + _1366;
    assign _1381 = _1367 + _1380;
    assign _5794 = _287 ? _1381 : _1351;
    assign _5800 = _278 ? _5799 : _5794;
    assign _61 = _5800;
    always @(posedge _272) begin
        if (_270)
            _1351 <= _290;
        else
            _1351 <= _61;
    end
    assign _1353 = _1351 == _290;
    assign _1354 = ~ _1353;
    assign _1348 = _265[53:53];
    assign _1355 = _1348 & _1354;
    assign _1358 = _1355 & _1357;
    assign _1386 = _1358 ? _1351 : _290;
    assign _1384 = _1378 ? _290 : _1371;
    assign _1387 = _1384 + _1386;
    assign _1401 = _1387 + _1400;
    assign _5801 = _287 ? _1401 : _1371;
    assign _5807 = _278 ? _5806 : _5801;
    assign _62 = _5807;
    always @(posedge _272) begin
        if (_270)
            _1371 <= _290;
        else
            _1371 <= _62;
    end
    assign _1373 = _1371 == _290;
    assign _1374 = ~ _1373;
    assign _1368 = _265[54:54];
    assign _1375 = _1368 & _1374;
    assign _1378 = _1375 & _1377;
    assign _1406 = _1378 ? _1371 : _290;
    assign _1404 = _1398 ? _290 : _1391;
    assign _1407 = _1404 + _1406;
    assign _1421 = _1407 + _1420;
    assign _5808 = _287 ? _1421 : _1391;
    assign _5814 = _278 ? _5813 : _5808;
    assign _63 = _5814;
    always @(posedge _272) begin
        if (_270)
            _1391 <= _290;
        else
            _1391 <= _63;
    end
    assign _1393 = _1391 == _290;
    assign _1394 = ~ _1393;
    assign _1388 = _265[55:55];
    assign _1395 = _1388 & _1394;
    assign _1398 = _1395 & _1397;
    assign _1426 = _1398 ? _1391 : _290;
    assign _1424 = _1418 ? _290 : _1411;
    assign _1427 = _1424 + _1426;
    assign _1441 = _1427 + _1440;
    assign _5815 = _287 ? _1441 : _1411;
    assign _5821 = _278 ? _5820 : _5815;
    assign _64 = _5821;
    always @(posedge _272) begin
        if (_270)
            _1411 <= _290;
        else
            _1411 <= _64;
    end
    assign _1413 = _1411 == _290;
    assign _1414 = ~ _1413;
    assign _1408 = _265[56:56];
    assign _1415 = _1408 & _1414;
    assign _1418 = _1415 & _1417;
    assign _1446 = _1418 ? _1411 : _290;
    assign _1444 = _1438 ? _290 : _1431;
    assign _1447 = _1444 + _1446;
    assign _1461 = _1447 + _1460;
    assign _5822 = _287 ? _1461 : _1431;
    assign _5828 = _278 ? _5827 : _5822;
    assign _65 = _5828;
    always @(posedge _272) begin
        if (_270)
            _1431 <= _290;
        else
            _1431 <= _65;
    end
    assign _1433 = _1431 == _290;
    assign _1434 = ~ _1433;
    assign _1428 = _265[57:57];
    assign _1435 = _1428 & _1434;
    assign _1438 = _1435 & _1437;
    assign _1466 = _1438 ? _1431 : _290;
    assign _1464 = _1458 ? _290 : _1451;
    assign _1467 = _1464 + _1466;
    assign _1481 = _1467 + _1480;
    assign _5829 = _287 ? _1481 : _1451;
    assign _5835 = _278 ? _5834 : _5829;
    assign _66 = _5835;
    always @(posedge _272) begin
        if (_270)
            _1451 <= _290;
        else
            _1451 <= _66;
    end
    assign _1453 = _1451 == _290;
    assign _1454 = ~ _1453;
    assign _1448 = _265[58:58];
    assign _1455 = _1448 & _1454;
    assign _1458 = _1455 & _1457;
    assign _1486 = _1458 ? _1451 : _290;
    assign _1484 = _1478 ? _290 : _1471;
    assign _1487 = _1484 + _1486;
    assign _1501 = _1487 + _1500;
    assign _5836 = _287 ? _1501 : _1471;
    assign _5842 = _278 ? _5841 : _5836;
    assign _67 = _5842;
    always @(posedge _272) begin
        if (_270)
            _1471 <= _290;
        else
            _1471 <= _67;
    end
    assign _1473 = _1471 == _290;
    assign _1474 = ~ _1473;
    assign _1468 = _265[59:59];
    assign _1475 = _1468 & _1474;
    assign _1478 = _1475 & _1477;
    assign _1506 = _1478 ? _1471 : _290;
    assign _1504 = _1498 ? _290 : _1491;
    assign _1507 = _1504 + _1506;
    assign _1521 = _1507 + _1520;
    assign _5843 = _287 ? _1521 : _1491;
    assign _5849 = _278 ? _5848 : _5843;
    assign _68 = _5849;
    always @(posedge _272) begin
        if (_270)
            _1491 <= _290;
        else
            _1491 <= _68;
    end
    assign _1493 = _1491 == _290;
    assign _1494 = ~ _1493;
    assign _1488 = _265[60:60];
    assign _1495 = _1488 & _1494;
    assign _1498 = _1495 & _1497;
    assign _1526 = _1498 ? _1491 : _290;
    assign _1524 = _1518 ? _290 : _1511;
    assign _1527 = _1524 + _1526;
    assign _1541 = _1527 + _1540;
    assign _5850 = _287 ? _1541 : _1511;
    assign _5856 = _278 ? _5855 : _5850;
    assign _69 = _5856;
    always @(posedge _272) begin
        if (_270)
            _1511 <= _290;
        else
            _1511 <= _69;
    end
    assign _1513 = _1511 == _290;
    assign _1514 = ~ _1513;
    assign _1508 = _265[61:61];
    assign _1515 = _1508 & _1514;
    assign _1518 = _1515 & _1517;
    assign _1546 = _1518 ? _1511 : _290;
    assign _1544 = _1538 ? _290 : _1531;
    assign _1547 = _1544 + _1546;
    assign _1561 = _1547 + _1560;
    assign _5857 = _287 ? _1561 : _1531;
    assign _5863 = _278 ? _5862 : _5857;
    assign _70 = _5863;
    always @(posedge _272) begin
        if (_270)
            _1531 <= _290;
        else
            _1531 <= _70;
    end
    assign _1533 = _1531 == _290;
    assign _1534 = ~ _1533;
    assign _1528 = _265[62:62];
    assign _1535 = _1528 & _1534;
    assign _1538 = _1535 & _1537;
    assign _1566 = _1538 ? _1531 : _290;
    assign _1564 = _1558 ? _290 : _1551;
    assign _1567 = _1564 + _1566;
    assign _1581 = _1567 + _1580;
    assign _5864 = _287 ? _1581 : _1551;
    assign _5870 = _278 ? _5869 : _5864;
    assign _71 = _5870;
    always @(posedge _272) begin
        if (_270)
            _1551 <= _290;
        else
            _1551 <= _71;
    end
    assign _1553 = _1551 == _290;
    assign _1554 = ~ _1553;
    assign _1548 = _265[63:63];
    assign _1555 = _1548 & _1554;
    assign _1558 = _1555 & _1557;
    assign _1586 = _1558 ? _1551 : _290;
    assign _1584 = _1578 ? _290 : _1571;
    assign _1587 = _1584 + _1586;
    assign _1601 = _1587 + _1600;
    assign _5871 = _287 ? _1601 : _1571;
    assign _5877 = _278 ? _5876 : _5871;
    assign _72 = _5877;
    always @(posedge _272) begin
        if (_270)
            _1571 <= _290;
        else
            _1571 <= _72;
    end
    assign _1573 = _1571 == _290;
    assign _1574 = ~ _1573;
    assign _1568 = _265[64:64];
    assign _1575 = _1568 & _1574;
    assign _1578 = _1575 & _1577;
    assign _1606 = _1578 ? _1571 : _290;
    assign _1604 = _1598 ? _290 : _1591;
    assign _1607 = _1604 + _1606;
    assign _1621 = _1607 + _1620;
    assign _5878 = _287 ? _1621 : _1591;
    assign _5884 = _278 ? _5883 : _5878;
    assign _73 = _5884;
    always @(posedge _272) begin
        if (_270)
            _1591 <= _290;
        else
            _1591 <= _73;
    end
    assign _1593 = _1591 == _290;
    assign _1594 = ~ _1593;
    assign _1588 = _265[65:65];
    assign _1595 = _1588 & _1594;
    assign _1598 = _1595 & _1597;
    assign _1626 = _1598 ? _1591 : _290;
    assign _1624 = _1618 ? _290 : _1611;
    assign _1627 = _1624 + _1626;
    assign _1641 = _1627 + _1640;
    assign _5885 = _287 ? _1641 : _1611;
    assign _5891 = _278 ? _5890 : _5885;
    assign _74 = _5891;
    always @(posedge _272) begin
        if (_270)
            _1611 <= _290;
        else
            _1611 <= _74;
    end
    assign _1613 = _1611 == _290;
    assign _1614 = ~ _1613;
    assign _1608 = _265[66:66];
    assign _1615 = _1608 & _1614;
    assign _1618 = _1615 & _1617;
    assign _1646 = _1618 ? _1611 : _290;
    assign _1644 = _1638 ? _290 : _1631;
    assign _1647 = _1644 + _1646;
    assign _1661 = _1647 + _1660;
    assign _5892 = _287 ? _1661 : _1631;
    assign _5898 = _278 ? _5897 : _5892;
    assign _75 = _5898;
    always @(posedge _272) begin
        if (_270)
            _1631 <= _290;
        else
            _1631 <= _75;
    end
    assign _1633 = _1631 == _290;
    assign _1634 = ~ _1633;
    assign _1628 = _265[67:67];
    assign _1635 = _1628 & _1634;
    assign _1638 = _1635 & _1637;
    assign _1666 = _1638 ? _1631 : _290;
    assign _1664 = _1658 ? _290 : _1651;
    assign _1667 = _1664 + _1666;
    assign _1681 = _1667 + _1680;
    assign _5899 = _287 ? _1681 : _1651;
    assign _5905 = _278 ? _5904 : _5899;
    assign _76 = _5905;
    always @(posedge _272) begin
        if (_270)
            _1651 <= _290;
        else
            _1651 <= _76;
    end
    assign _1653 = _1651 == _290;
    assign _1654 = ~ _1653;
    assign _1648 = _265[68:68];
    assign _1655 = _1648 & _1654;
    assign _1658 = _1655 & _1657;
    assign _1686 = _1658 ? _1651 : _290;
    assign _1684 = _1678 ? _290 : _1671;
    assign _1687 = _1684 + _1686;
    assign _1701 = _1687 + _1700;
    assign _5906 = _287 ? _1701 : _1671;
    assign _5912 = _278 ? _5911 : _5906;
    assign _77 = _5912;
    always @(posedge _272) begin
        if (_270)
            _1671 <= _290;
        else
            _1671 <= _77;
    end
    assign _1673 = _1671 == _290;
    assign _1674 = ~ _1673;
    assign _1668 = _265[69:69];
    assign _1675 = _1668 & _1674;
    assign _1678 = _1675 & _1677;
    assign _1706 = _1678 ? _1671 : _290;
    assign _1704 = _1698 ? _290 : _1691;
    assign _1707 = _1704 + _1706;
    assign _1721 = _1707 + _1720;
    assign _5913 = _287 ? _1721 : _1691;
    assign _5919 = _278 ? _5918 : _5913;
    assign _78 = _5919;
    always @(posedge _272) begin
        if (_270)
            _1691 <= _290;
        else
            _1691 <= _78;
    end
    assign _1693 = _1691 == _290;
    assign _1694 = ~ _1693;
    assign _1688 = _265[70:70];
    assign _1695 = _1688 & _1694;
    assign _1698 = _1695 & _1697;
    assign _1726 = _1698 ? _1691 : _290;
    assign _1724 = _1718 ? _290 : _1711;
    assign _1727 = _1724 + _1726;
    assign _1741 = _1727 + _1740;
    assign _5920 = _287 ? _1741 : _1711;
    assign _5926 = _278 ? _5925 : _5920;
    assign _79 = _5926;
    always @(posedge _272) begin
        if (_270)
            _1711 <= _290;
        else
            _1711 <= _79;
    end
    assign _1713 = _1711 == _290;
    assign _1714 = ~ _1713;
    assign _1708 = _265[71:71];
    assign _1715 = _1708 & _1714;
    assign _1718 = _1715 & _1717;
    assign _1746 = _1718 ? _1711 : _290;
    assign _1744 = _1738 ? _290 : _1731;
    assign _1747 = _1744 + _1746;
    assign _1761 = _1747 + _1760;
    assign _5927 = _287 ? _1761 : _1731;
    assign _5933 = _278 ? _5932 : _5927;
    assign _80 = _5933;
    always @(posedge _272) begin
        if (_270)
            _1731 <= _290;
        else
            _1731 <= _80;
    end
    assign _1733 = _1731 == _290;
    assign _1734 = ~ _1733;
    assign _1728 = _265[72:72];
    assign _1735 = _1728 & _1734;
    assign _1738 = _1735 & _1737;
    assign _1766 = _1738 ? _1731 : _290;
    assign _1764 = _1758 ? _290 : _1751;
    assign _1767 = _1764 + _1766;
    assign _1781 = _1767 + _1780;
    assign _5934 = _287 ? _1781 : _1751;
    assign _5940 = _278 ? _5939 : _5934;
    assign _81 = _5940;
    always @(posedge _272) begin
        if (_270)
            _1751 <= _290;
        else
            _1751 <= _81;
    end
    assign _1753 = _1751 == _290;
    assign _1754 = ~ _1753;
    assign _1748 = _265[73:73];
    assign _1755 = _1748 & _1754;
    assign _1758 = _1755 & _1757;
    assign _1786 = _1758 ? _1751 : _290;
    assign _1784 = _1778 ? _290 : _1771;
    assign _1787 = _1784 + _1786;
    assign _1801 = _1787 + _1800;
    assign _5941 = _287 ? _1801 : _1771;
    assign _5947 = _278 ? _5946 : _5941;
    assign _82 = _5947;
    always @(posedge _272) begin
        if (_270)
            _1771 <= _290;
        else
            _1771 <= _82;
    end
    assign _1773 = _1771 == _290;
    assign _1774 = ~ _1773;
    assign _1768 = _265[74:74];
    assign _1775 = _1768 & _1774;
    assign _1778 = _1775 & _1777;
    assign _1806 = _1778 ? _1771 : _290;
    assign _1804 = _1798 ? _290 : _1791;
    assign _1807 = _1804 + _1806;
    assign _1821 = _1807 + _1820;
    assign _5948 = _287 ? _1821 : _1791;
    assign _5954 = _278 ? _5953 : _5948;
    assign _83 = _5954;
    always @(posedge _272) begin
        if (_270)
            _1791 <= _290;
        else
            _1791 <= _83;
    end
    assign _1793 = _1791 == _290;
    assign _1794 = ~ _1793;
    assign _1788 = _265[75:75];
    assign _1795 = _1788 & _1794;
    assign _1798 = _1795 & _1797;
    assign _1826 = _1798 ? _1791 : _290;
    assign _1824 = _1818 ? _290 : _1811;
    assign _1827 = _1824 + _1826;
    assign _1841 = _1827 + _1840;
    assign _5955 = _287 ? _1841 : _1811;
    assign _5961 = _278 ? _5960 : _5955;
    assign _84 = _5961;
    always @(posedge _272) begin
        if (_270)
            _1811 <= _290;
        else
            _1811 <= _84;
    end
    assign _1813 = _1811 == _290;
    assign _1814 = ~ _1813;
    assign _1808 = _265[76:76];
    assign _1815 = _1808 & _1814;
    assign _1818 = _1815 & _1817;
    assign _1846 = _1818 ? _1811 : _290;
    assign _1844 = _1838 ? _290 : _1831;
    assign _1847 = _1844 + _1846;
    assign _1861 = _1847 + _1860;
    assign _5962 = _287 ? _1861 : _1831;
    assign _5968 = _278 ? _5967 : _5962;
    assign _85 = _5968;
    always @(posedge _272) begin
        if (_270)
            _1831 <= _290;
        else
            _1831 <= _85;
    end
    assign _1833 = _1831 == _290;
    assign _1834 = ~ _1833;
    assign _1828 = _265[77:77];
    assign _1835 = _1828 & _1834;
    assign _1838 = _1835 & _1837;
    assign _1866 = _1838 ? _1831 : _290;
    assign _1864 = _1858 ? _290 : _1851;
    assign _1867 = _1864 + _1866;
    assign _1881 = _1867 + _1880;
    assign _5969 = _287 ? _1881 : _1851;
    assign _5975 = _278 ? _5974 : _5969;
    assign _86 = _5975;
    always @(posedge _272) begin
        if (_270)
            _1851 <= _290;
        else
            _1851 <= _86;
    end
    assign _1853 = _1851 == _290;
    assign _1854 = ~ _1853;
    assign _1848 = _265[78:78];
    assign _1855 = _1848 & _1854;
    assign _1858 = _1855 & _1857;
    assign _1886 = _1858 ? _1851 : _290;
    assign _1884 = _1878 ? _290 : _1871;
    assign _1887 = _1884 + _1886;
    assign _1901 = _1887 + _1900;
    assign _5976 = _287 ? _1901 : _1871;
    assign _5982 = _278 ? _5981 : _5976;
    assign _87 = _5982;
    always @(posedge _272) begin
        if (_270)
            _1871 <= _290;
        else
            _1871 <= _87;
    end
    assign _1873 = _1871 == _290;
    assign _1874 = ~ _1873;
    assign _1868 = _265[79:79];
    assign _1875 = _1868 & _1874;
    assign _1878 = _1875 & _1877;
    assign _1906 = _1878 ? _1871 : _290;
    assign _1904 = _1898 ? _290 : _1891;
    assign _1907 = _1904 + _1906;
    assign _1921 = _1907 + _1920;
    assign _5983 = _287 ? _1921 : _1891;
    assign _5989 = _278 ? _5988 : _5983;
    assign _88 = _5989;
    always @(posedge _272) begin
        if (_270)
            _1891 <= _290;
        else
            _1891 <= _88;
    end
    assign _1893 = _1891 == _290;
    assign _1894 = ~ _1893;
    assign _1888 = _265[80:80];
    assign _1895 = _1888 & _1894;
    assign _1898 = _1895 & _1897;
    assign _1926 = _1898 ? _1891 : _290;
    assign _1924 = _1918 ? _290 : _1911;
    assign _1927 = _1924 + _1926;
    assign _1941 = _1927 + _1940;
    assign _5990 = _287 ? _1941 : _1911;
    assign _5996 = _278 ? _5995 : _5990;
    assign _89 = _5996;
    always @(posedge _272) begin
        if (_270)
            _1911 <= _290;
        else
            _1911 <= _89;
    end
    assign _1913 = _1911 == _290;
    assign _1914 = ~ _1913;
    assign _1908 = _265[81:81];
    assign _1915 = _1908 & _1914;
    assign _1918 = _1915 & _1917;
    assign _1946 = _1918 ? _1911 : _290;
    assign _1944 = _1938 ? _290 : _1931;
    assign _1947 = _1944 + _1946;
    assign _1961 = _1947 + _1960;
    assign _5997 = _287 ? _1961 : _1931;
    assign _6003 = _278 ? _6002 : _5997;
    assign _90 = _6003;
    always @(posedge _272) begin
        if (_270)
            _1931 <= _290;
        else
            _1931 <= _90;
    end
    assign _1933 = _1931 == _290;
    assign _1934 = ~ _1933;
    assign _1928 = _265[82:82];
    assign _1935 = _1928 & _1934;
    assign _1938 = _1935 & _1937;
    assign _1966 = _1938 ? _1931 : _290;
    assign _1964 = _1958 ? _290 : _1951;
    assign _1967 = _1964 + _1966;
    assign _1981 = _1967 + _1980;
    assign _6004 = _287 ? _1981 : _1951;
    assign _6010 = _278 ? _6009 : _6004;
    assign _91 = _6010;
    always @(posedge _272) begin
        if (_270)
            _1951 <= _290;
        else
            _1951 <= _91;
    end
    assign _1953 = _1951 == _290;
    assign _1954 = ~ _1953;
    assign _1948 = _265[83:83];
    assign _1955 = _1948 & _1954;
    assign _1958 = _1955 & _1957;
    assign _1986 = _1958 ? _1951 : _290;
    assign _1984 = _1978 ? _290 : _1971;
    assign _1987 = _1984 + _1986;
    assign _2001 = _1987 + _2000;
    assign _6011 = _287 ? _2001 : _1971;
    assign _6017 = _278 ? _6016 : _6011;
    assign _92 = _6017;
    always @(posedge _272) begin
        if (_270)
            _1971 <= _290;
        else
            _1971 <= _92;
    end
    assign _1973 = _1971 == _290;
    assign _1974 = ~ _1973;
    assign _1968 = _265[84:84];
    assign _1975 = _1968 & _1974;
    assign _1978 = _1975 & _1977;
    assign _2006 = _1978 ? _1971 : _290;
    assign _2004 = _1998 ? _290 : _1991;
    assign _2007 = _2004 + _2006;
    assign _2021 = _2007 + _2020;
    assign _6018 = _287 ? _2021 : _1991;
    assign _6024 = _278 ? _6023 : _6018;
    assign _93 = _6024;
    always @(posedge _272) begin
        if (_270)
            _1991 <= _290;
        else
            _1991 <= _93;
    end
    assign _1993 = _1991 == _290;
    assign _1994 = ~ _1993;
    assign _1988 = _265[85:85];
    assign _1995 = _1988 & _1994;
    assign _1998 = _1995 & _1997;
    assign _2026 = _1998 ? _1991 : _290;
    assign _2024 = _2018 ? _290 : _2011;
    assign _2027 = _2024 + _2026;
    assign _2041 = _2027 + _2040;
    assign _6025 = _287 ? _2041 : _2011;
    assign _6031 = _278 ? _6030 : _6025;
    assign _94 = _6031;
    always @(posedge _272) begin
        if (_270)
            _2011 <= _290;
        else
            _2011 <= _94;
    end
    assign _2013 = _2011 == _290;
    assign _2014 = ~ _2013;
    assign _2008 = _265[86:86];
    assign _2015 = _2008 & _2014;
    assign _2018 = _2015 & _2017;
    assign _2046 = _2018 ? _2011 : _290;
    assign _2044 = _2038 ? _290 : _2031;
    assign _2047 = _2044 + _2046;
    assign _2061 = _2047 + _2060;
    assign _6032 = _287 ? _2061 : _2031;
    assign _6038 = _278 ? _6037 : _6032;
    assign _95 = _6038;
    always @(posedge _272) begin
        if (_270)
            _2031 <= _290;
        else
            _2031 <= _95;
    end
    assign _2033 = _2031 == _290;
    assign _2034 = ~ _2033;
    assign _2028 = _265[87:87];
    assign _2035 = _2028 & _2034;
    assign _2038 = _2035 & _2037;
    assign _2066 = _2038 ? _2031 : _290;
    assign _2064 = _2058 ? _290 : _2051;
    assign _2067 = _2064 + _2066;
    assign _2081 = _2067 + _2080;
    assign _6039 = _287 ? _2081 : _2051;
    assign _6045 = _278 ? _6044 : _6039;
    assign _96 = _6045;
    always @(posedge _272) begin
        if (_270)
            _2051 <= _290;
        else
            _2051 <= _96;
    end
    assign _2053 = _2051 == _290;
    assign _2054 = ~ _2053;
    assign _2048 = _265[88:88];
    assign _2055 = _2048 & _2054;
    assign _2058 = _2055 & _2057;
    assign _2086 = _2058 ? _2051 : _290;
    assign _2084 = _2078 ? _290 : _2071;
    assign _2087 = _2084 + _2086;
    assign _2101 = _2087 + _2100;
    assign _6046 = _287 ? _2101 : _2071;
    assign _6052 = _278 ? _6051 : _6046;
    assign _97 = _6052;
    always @(posedge _272) begin
        if (_270)
            _2071 <= _290;
        else
            _2071 <= _97;
    end
    assign _2073 = _2071 == _290;
    assign _2074 = ~ _2073;
    assign _2068 = _265[89:89];
    assign _2075 = _2068 & _2074;
    assign _2078 = _2075 & _2077;
    assign _2106 = _2078 ? _2071 : _290;
    assign _2104 = _2098 ? _290 : _2091;
    assign _2107 = _2104 + _2106;
    assign _2121 = _2107 + _2120;
    assign _6053 = _287 ? _2121 : _2091;
    assign _6059 = _278 ? _6058 : _6053;
    assign _98 = _6059;
    always @(posedge _272) begin
        if (_270)
            _2091 <= _290;
        else
            _2091 <= _98;
    end
    assign _2093 = _2091 == _290;
    assign _2094 = ~ _2093;
    assign _2088 = _265[90:90];
    assign _2095 = _2088 & _2094;
    assign _2098 = _2095 & _2097;
    assign _2126 = _2098 ? _2091 : _290;
    assign _2124 = _2118 ? _290 : _2111;
    assign _2127 = _2124 + _2126;
    assign _2141 = _2127 + _2140;
    assign _6060 = _287 ? _2141 : _2111;
    assign _6066 = _278 ? _6065 : _6060;
    assign _99 = _6066;
    always @(posedge _272) begin
        if (_270)
            _2111 <= _290;
        else
            _2111 <= _99;
    end
    assign _2113 = _2111 == _290;
    assign _2114 = ~ _2113;
    assign _2108 = _265[91:91];
    assign _2115 = _2108 & _2114;
    assign _2118 = _2115 & _2117;
    assign _2146 = _2118 ? _2111 : _290;
    assign _2144 = _2138 ? _290 : _2131;
    assign _2147 = _2144 + _2146;
    assign _2161 = _2147 + _2160;
    assign _6067 = _287 ? _2161 : _2131;
    assign _6073 = _278 ? _6072 : _6067;
    assign _100 = _6073;
    always @(posedge _272) begin
        if (_270)
            _2131 <= _290;
        else
            _2131 <= _100;
    end
    assign _2133 = _2131 == _290;
    assign _2134 = ~ _2133;
    assign _2128 = _265[92:92];
    assign _2135 = _2128 & _2134;
    assign _2138 = _2135 & _2137;
    assign _2166 = _2138 ? _2131 : _290;
    assign _2164 = _2158 ? _290 : _2151;
    assign _2167 = _2164 + _2166;
    assign _2181 = _2167 + _2180;
    assign _6074 = _287 ? _2181 : _2151;
    assign _6080 = _278 ? _6079 : _6074;
    assign _101 = _6080;
    always @(posedge _272) begin
        if (_270)
            _2151 <= _290;
        else
            _2151 <= _101;
    end
    assign _2153 = _2151 == _290;
    assign _2154 = ~ _2153;
    assign _2148 = _265[93:93];
    assign _2155 = _2148 & _2154;
    assign _2158 = _2155 & _2157;
    assign _2186 = _2158 ? _2151 : _290;
    assign _2184 = _2178 ? _290 : _2171;
    assign _2187 = _2184 + _2186;
    assign _2201 = _2187 + _2200;
    assign _6081 = _287 ? _2201 : _2171;
    assign _6087 = _278 ? _6086 : _6081;
    assign _102 = _6087;
    always @(posedge _272) begin
        if (_270)
            _2171 <= _290;
        else
            _2171 <= _102;
    end
    assign _2173 = _2171 == _290;
    assign _2174 = ~ _2173;
    assign _2168 = _265[94:94];
    assign _2175 = _2168 & _2174;
    assign _2178 = _2175 & _2177;
    assign _2206 = _2178 ? _2171 : _290;
    assign _2204 = _2198 ? _290 : _2191;
    assign _2207 = _2204 + _2206;
    assign _2221 = _2207 + _2220;
    assign _6088 = _287 ? _2221 : _2191;
    assign _6094 = _278 ? _6093 : _6088;
    assign _103 = _6094;
    always @(posedge _272) begin
        if (_270)
            _2191 <= _290;
        else
            _2191 <= _103;
    end
    assign _2193 = _2191 == _290;
    assign _2194 = ~ _2193;
    assign _2188 = _265[95:95];
    assign _2195 = _2188 & _2194;
    assign _2198 = _2195 & _2197;
    assign _2226 = _2198 ? _2191 : _290;
    assign _2224 = _2218 ? _290 : _2211;
    assign _2227 = _2224 + _2226;
    assign _2241 = _2227 + _2240;
    assign _6095 = _287 ? _2241 : _2211;
    assign _6101 = _278 ? _6100 : _6095;
    assign _104 = _6101;
    always @(posedge _272) begin
        if (_270)
            _2211 <= _290;
        else
            _2211 <= _104;
    end
    assign _2213 = _2211 == _290;
    assign _2214 = ~ _2213;
    assign _2208 = _265[96:96];
    assign _2215 = _2208 & _2214;
    assign _2218 = _2215 & _2217;
    assign _2246 = _2218 ? _2211 : _290;
    assign _2244 = _2238 ? _290 : _2231;
    assign _2247 = _2244 + _2246;
    assign _2261 = _2247 + _2260;
    assign _6102 = _287 ? _2261 : _2231;
    assign _6108 = _278 ? _6107 : _6102;
    assign _105 = _6108;
    always @(posedge _272) begin
        if (_270)
            _2231 <= _290;
        else
            _2231 <= _105;
    end
    assign _2233 = _2231 == _290;
    assign _2234 = ~ _2233;
    assign _2228 = _265[97:97];
    assign _2235 = _2228 & _2234;
    assign _2238 = _2235 & _2237;
    assign _2266 = _2238 ? _2231 : _290;
    assign _2264 = _2258 ? _290 : _2251;
    assign _2267 = _2264 + _2266;
    assign _2281 = _2267 + _2280;
    assign _6109 = _287 ? _2281 : _2251;
    assign _6115 = _278 ? _6114 : _6109;
    assign _106 = _6115;
    always @(posedge _272) begin
        if (_270)
            _2251 <= _290;
        else
            _2251 <= _106;
    end
    assign _2253 = _2251 == _290;
    assign _2254 = ~ _2253;
    assign _2248 = _265[98:98];
    assign _2255 = _2248 & _2254;
    assign _2258 = _2255 & _2257;
    assign _2286 = _2258 ? _2251 : _290;
    assign _2284 = _2278 ? _290 : _2271;
    assign _2287 = _2284 + _2286;
    assign _2301 = _2287 + _2300;
    assign _6116 = _287 ? _2301 : _2271;
    assign _6122 = _278 ? _6121 : _6116;
    assign _107 = _6122;
    always @(posedge _272) begin
        if (_270)
            _2271 <= _290;
        else
            _2271 <= _107;
    end
    assign _2273 = _2271 == _290;
    assign _2274 = ~ _2273;
    assign _2268 = _265[99:99];
    assign _2275 = _2268 & _2274;
    assign _2278 = _2275 & _2277;
    assign _2306 = _2278 ? _2271 : _290;
    assign _2304 = _2298 ? _290 : _2291;
    assign _2307 = _2304 + _2306;
    assign _2321 = _2307 + _2320;
    assign _6123 = _287 ? _2321 : _2291;
    assign _6129 = _278 ? _6128 : _6123;
    assign _108 = _6129;
    always @(posedge _272) begin
        if (_270)
            _2291 <= _290;
        else
            _2291 <= _108;
    end
    assign _2293 = _2291 == _290;
    assign _2294 = ~ _2293;
    assign _2288 = _265[100:100];
    assign _2295 = _2288 & _2294;
    assign _2298 = _2295 & _2297;
    assign _2326 = _2298 ? _2291 : _290;
    assign _2324 = _2318 ? _290 : _2311;
    assign _2327 = _2324 + _2326;
    assign _2341 = _2327 + _2340;
    assign _6130 = _287 ? _2341 : _2311;
    assign _6136 = _278 ? _6135 : _6130;
    assign _109 = _6136;
    always @(posedge _272) begin
        if (_270)
            _2311 <= _290;
        else
            _2311 <= _109;
    end
    assign _2313 = _2311 == _290;
    assign _2314 = ~ _2313;
    assign _2308 = _265[101:101];
    assign _2315 = _2308 & _2314;
    assign _2318 = _2315 & _2317;
    assign _2346 = _2318 ? _2311 : _290;
    assign _2344 = _2338 ? _290 : _2331;
    assign _2347 = _2344 + _2346;
    assign _2361 = _2347 + _2360;
    assign _6137 = _287 ? _2361 : _2331;
    assign _6143 = _278 ? _6142 : _6137;
    assign _110 = _6143;
    always @(posedge _272) begin
        if (_270)
            _2331 <= _290;
        else
            _2331 <= _110;
    end
    assign _2333 = _2331 == _290;
    assign _2334 = ~ _2333;
    assign _2328 = _265[102:102];
    assign _2335 = _2328 & _2334;
    assign _2338 = _2335 & _2337;
    assign _2366 = _2338 ? _2331 : _290;
    assign _2364 = _2358 ? _290 : _2351;
    assign _2367 = _2364 + _2366;
    assign _2381 = _2367 + _2380;
    assign _6144 = _287 ? _2381 : _2351;
    assign _6150 = _278 ? _6149 : _6144;
    assign _111 = _6150;
    always @(posedge _272) begin
        if (_270)
            _2351 <= _290;
        else
            _2351 <= _111;
    end
    assign _2353 = _2351 == _290;
    assign _2354 = ~ _2353;
    assign _2348 = _265[103:103];
    assign _2355 = _2348 & _2354;
    assign _2358 = _2355 & _2357;
    assign _2386 = _2358 ? _2351 : _290;
    assign _2384 = _2378 ? _290 : _2371;
    assign _2387 = _2384 + _2386;
    assign _2401 = _2387 + _2400;
    assign _6151 = _287 ? _2401 : _2371;
    assign _6157 = _278 ? _6156 : _6151;
    assign _112 = _6157;
    always @(posedge _272) begin
        if (_270)
            _2371 <= _290;
        else
            _2371 <= _112;
    end
    assign _2373 = _2371 == _290;
    assign _2374 = ~ _2373;
    assign _2368 = _265[104:104];
    assign _2375 = _2368 & _2374;
    assign _2378 = _2375 & _2377;
    assign _2406 = _2378 ? _2371 : _290;
    assign _2404 = _2398 ? _290 : _2391;
    assign _2407 = _2404 + _2406;
    assign _2421 = _2407 + _2420;
    assign _6158 = _287 ? _2421 : _2391;
    assign _6164 = _278 ? _6163 : _6158;
    assign _113 = _6164;
    always @(posedge _272) begin
        if (_270)
            _2391 <= _290;
        else
            _2391 <= _113;
    end
    assign _2393 = _2391 == _290;
    assign _2394 = ~ _2393;
    assign _2388 = _265[105:105];
    assign _2395 = _2388 & _2394;
    assign _2398 = _2395 & _2397;
    assign _2426 = _2398 ? _2391 : _290;
    assign _2424 = _2418 ? _290 : _2411;
    assign _2427 = _2424 + _2426;
    assign _2441 = _2427 + _2440;
    assign _6165 = _287 ? _2441 : _2411;
    assign _6171 = _278 ? _6170 : _6165;
    assign _114 = _6171;
    always @(posedge _272) begin
        if (_270)
            _2411 <= _290;
        else
            _2411 <= _114;
    end
    assign _2413 = _2411 == _290;
    assign _2414 = ~ _2413;
    assign _2408 = _265[106:106];
    assign _2415 = _2408 & _2414;
    assign _2418 = _2415 & _2417;
    assign _2446 = _2418 ? _2411 : _290;
    assign _2444 = _2438 ? _290 : _2431;
    assign _2447 = _2444 + _2446;
    assign _2461 = _2447 + _2460;
    assign _6172 = _287 ? _2461 : _2431;
    assign _6178 = _278 ? _6177 : _6172;
    assign _115 = _6178;
    always @(posedge _272) begin
        if (_270)
            _2431 <= _290;
        else
            _2431 <= _115;
    end
    assign _2433 = _2431 == _290;
    assign _2434 = ~ _2433;
    assign _2428 = _265[107:107];
    assign _2435 = _2428 & _2434;
    assign _2438 = _2435 & _2437;
    assign _2466 = _2438 ? _2431 : _290;
    assign _2464 = _2458 ? _290 : _2451;
    assign _2467 = _2464 + _2466;
    assign _2481 = _2467 + _2480;
    assign _6179 = _287 ? _2481 : _2451;
    assign _6185 = _278 ? _6184 : _6179;
    assign _116 = _6185;
    always @(posedge _272) begin
        if (_270)
            _2451 <= _290;
        else
            _2451 <= _116;
    end
    assign _2453 = _2451 == _290;
    assign _2454 = ~ _2453;
    assign _2448 = _265[108:108];
    assign _2455 = _2448 & _2454;
    assign _2458 = _2455 & _2457;
    assign _2486 = _2458 ? _2451 : _290;
    assign _2484 = _2478 ? _290 : _2471;
    assign _2487 = _2484 + _2486;
    assign _2501 = _2487 + _2500;
    assign _6186 = _287 ? _2501 : _2471;
    assign _6192 = _278 ? _6191 : _6186;
    assign _117 = _6192;
    always @(posedge _272) begin
        if (_270)
            _2471 <= _290;
        else
            _2471 <= _117;
    end
    assign _2473 = _2471 == _290;
    assign _2474 = ~ _2473;
    assign _2468 = _265[109:109];
    assign _2475 = _2468 & _2474;
    assign _2478 = _2475 & _2477;
    assign _2506 = _2478 ? _2471 : _290;
    assign _2504 = _2498 ? _290 : _2491;
    assign _2507 = _2504 + _2506;
    assign _2521 = _2507 + _2520;
    assign _6193 = _287 ? _2521 : _2491;
    assign _6199 = _278 ? _6198 : _6193;
    assign _118 = _6199;
    always @(posedge _272) begin
        if (_270)
            _2491 <= _290;
        else
            _2491 <= _118;
    end
    assign _2493 = _2491 == _290;
    assign _2494 = ~ _2493;
    assign _2488 = _265[110:110];
    assign _2495 = _2488 & _2494;
    assign _2498 = _2495 & _2497;
    assign _2526 = _2498 ? _2491 : _290;
    assign _2524 = _2518 ? _290 : _2511;
    assign _2527 = _2524 + _2526;
    assign _2541 = _2527 + _2540;
    assign _6200 = _287 ? _2541 : _2511;
    assign _6206 = _278 ? _6205 : _6200;
    assign _119 = _6206;
    always @(posedge _272) begin
        if (_270)
            _2511 <= _290;
        else
            _2511 <= _119;
    end
    assign _2513 = _2511 == _290;
    assign _2514 = ~ _2513;
    assign _2508 = _265[111:111];
    assign _2515 = _2508 & _2514;
    assign _2518 = _2515 & _2517;
    assign _2546 = _2518 ? _2511 : _290;
    assign _2544 = _2538 ? _290 : _2531;
    assign _2547 = _2544 + _2546;
    assign _2561 = _2547 + _2560;
    assign _6207 = _287 ? _2561 : _2531;
    assign _6213 = _278 ? _6212 : _6207;
    assign _120 = _6213;
    always @(posedge _272) begin
        if (_270)
            _2531 <= _290;
        else
            _2531 <= _120;
    end
    assign _2533 = _2531 == _290;
    assign _2534 = ~ _2533;
    assign _2528 = _265[112:112];
    assign _2535 = _2528 & _2534;
    assign _2538 = _2535 & _2537;
    assign _2566 = _2538 ? _2531 : _290;
    assign _2564 = _2558 ? _290 : _2551;
    assign _2567 = _2564 + _2566;
    assign _2581 = _2567 + _2580;
    assign _6214 = _287 ? _2581 : _2551;
    assign _6220 = _278 ? _6219 : _6214;
    assign _121 = _6220;
    always @(posedge _272) begin
        if (_270)
            _2551 <= _290;
        else
            _2551 <= _121;
    end
    assign _2553 = _2551 == _290;
    assign _2554 = ~ _2553;
    assign _2548 = _265[113:113];
    assign _2555 = _2548 & _2554;
    assign _2558 = _2555 & _2557;
    assign _2586 = _2558 ? _2551 : _290;
    assign _2584 = _2578 ? _290 : _2571;
    assign _2587 = _2584 + _2586;
    assign _2601 = _2587 + _2600;
    assign _6221 = _287 ? _2601 : _2571;
    assign _6227 = _278 ? _6226 : _6221;
    assign _122 = _6227;
    always @(posedge _272) begin
        if (_270)
            _2571 <= _290;
        else
            _2571 <= _122;
    end
    assign _2573 = _2571 == _290;
    assign _2574 = ~ _2573;
    assign _2568 = _265[114:114];
    assign _2575 = _2568 & _2574;
    assign _2578 = _2575 & _2577;
    assign _2606 = _2578 ? _2571 : _290;
    assign _2604 = _2598 ? _290 : _2591;
    assign _2607 = _2604 + _2606;
    assign _2621 = _2607 + _2620;
    assign _6228 = _287 ? _2621 : _2591;
    assign _6234 = _278 ? _6233 : _6228;
    assign _123 = _6234;
    always @(posedge _272) begin
        if (_270)
            _2591 <= _290;
        else
            _2591 <= _123;
    end
    assign _2593 = _2591 == _290;
    assign _2594 = ~ _2593;
    assign _2588 = _265[115:115];
    assign _2595 = _2588 & _2594;
    assign _2598 = _2595 & _2597;
    assign _2626 = _2598 ? _2591 : _290;
    assign _2624 = _2618 ? _290 : _2611;
    assign _2627 = _2624 + _2626;
    assign _2641 = _2627 + _2640;
    assign _6235 = _287 ? _2641 : _2611;
    assign _6241 = _278 ? _6240 : _6235;
    assign _124 = _6241;
    always @(posedge _272) begin
        if (_270)
            _2611 <= _290;
        else
            _2611 <= _124;
    end
    assign _2613 = _2611 == _290;
    assign _2614 = ~ _2613;
    assign _2608 = _265[116:116];
    assign _2615 = _2608 & _2614;
    assign _2618 = _2615 & _2617;
    assign _2646 = _2618 ? _2611 : _290;
    assign _2644 = _2638 ? _290 : _2631;
    assign _2647 = _2644 + _2646;
    assign _2661 = _2647 + _2660;
    assign _6242 = _287 ? _2661 : _2631;
    assign _6248 = _278 ? _6247 : _6242;
    assign _125 = _6248;
    always @(posedge _272) begin
        if (_270)
            _2631 <= _290;
        else
            _2631 <= _125;
    end
    assign _2633 = _2631 == _290;
    assign _2634 = ~ _2633;
    assign _2628 = _265[117:117];
    assign _2635 = _2628 & _2634;
    assign _2638 = _2635 & _2637;
    assign _2666 = _2638 ? _2631 : _290;
    assign _2664 = _2658 ? _290 : _2651;
    assign _2667 = _2664 + _2666;
    assign _2681 = _2667 + _2680;
    assign _6249 = _287 ? _2681 : _2651;
    assign _6255 = _278 ? _6254 : _6249;
    assign _126 = _6255;
    always @(posedge _272) begin
        if (_270)
            _2651 <= _290;
        else
            _2651 <= _126;
    end
    assign _2653 = _2651 == _290;
    assign _2654 = ~ _2653;
    assign _2648 = _265[118:118];
    assign _2655 = _2648 & _2654;
    assign _2658 = _2655 & _2657;
    assign _2686 = _2658 ? _2651 : _290;
    assign _2684 = _2678 ? _290 : _2671;
    assign _2687 = _2684 + _2686;
    assign _2701 = _2687 + _2700;
    assign _6256 = _287 ? _2701 : _2671;
    assign _6262 = _278 ? _6261 : _6256;
    assign _127 = _6262;
    always @(posedge _272) begin
        if (_270)
            _2671 <= _290;
        else
            _2671 <= _127;
    end
    assign _2673 = _2671 == _290;
    assign _2674 = ~ _2673;
    assign _2668 = _265[119:119];
    assign _2675 = _2668 & _2674;
    assign _2678 = _2675 & _2677;
    assign _2706 = _2678 ? _2671 : _290;
    assign _2704 = _2698 ? _290 : _2691;
    assign _2707 = _2704 + _2706;
    assign _2721 = _2707 + _2720;
    assign _6263 = _287 ? _2721 : _2691;
    assign _6269 = _278 ? _6268 : _6263;
    assign _128 = _6269;
    always @(posedge _272) begin
        if (_270)
            _2691 <= _290;
        else
            _2691 <= _128;
    end
    assign _2693 = _2691 == _290;
    assign _2694 = ~ _2693;
    assign _2688 = _265[120:120];
    assign _2695 = _2688 & _2694;
    assign _2698 = _2695 & _2697;
    assign _2726 = _2698 ? _2691 : _290;
    assign _2724 = _2718 ? _290 : _2711;
    assign _2727 = _2724 + _2726;
    assign _2741 = _2727 + _2740;
    assign _6270 = _287 ? _2741 : _2711;
    assign _6276 = _278 ? _6275 : _6270;
    assign _129 = _6276;
    always @(posedge _272) begin
        if (_270)
            _2711 <= _290;
        else
            _2711 <= _129;
    end
    assign _2713 = _2711 == _290;
    assign _2714 = ~ _2713;
    assign _2708 = _265[121:121];
    assign _2715 = _2708 & _2714;
    assign _2718 = _2715 & _2717;
    assign _2746 = _2718 ? _2711 : _290;
    assign _2744 = _2738 ? _290 : _2731;
    assign _2747 = _2744 + _2746;
    assign _2761 = _2747 + _2760;
    assign _6277 = _287 ? _2761 : _2731;
    assign _6283 = _278 ? _6282 : _6277;
    assign _130 = _6283;
    always @(posedge _272) begin
        if (_270)
            _2731 <= _290;
        else
            _2731 <= _130;
    end
    assign _2733 = _2731 == _290;
    assign _2734 = ~ _2733;
    assign _2728 = _265[122:122];
    assign _2735 = _2728 & _2734;
    assign _2738 = _2735 & _2737;
    assign _2766 = _2738 ? _2731 : _290;
    assign _2764 = _2758 ? _290 : _2751;
    assign _2767 = _2764 + _2766;
    assign _2781 = _2767 + _2780;
    assign _6284 = _287 ? _2781 : _2751;
    assign _6290 = _278 ? _6289 : _6284;
    assign _131 = _6290;
    always @(posedge _272) begin
        if (_270)
            _2751 <= _290;
        else
            _2751 <= _131;
    end
    assign _2753 = _2751 == _290;
    assign _2754 = ~ _2753;
    assign _2748 = _265[123:123];
    assign _2755 = _2748 & _2754;
    assign _2758 = _2755 & _2757;
    assign _2786 = _2758 ? _2751 : _290;
    assign _2784 = _2778 ? _290 : _2771;
    assign _2787 = _2784 + _2786;
    assign _2801 = _2787 + _2800;
    assign _6291 = _287 ? _2801 : _2771;
    assign _6297 = _278 ? _6296 : _6291;
    assign _132 = _6297;
    always @(posedge _272) begin
        if (_270)
            _2771 <= _290;
        else
            _2771 <= _132;
    end
    assign _2773 = _2771 == _290;
    assign _2774 = ~ _2773;
    assign _2768 = _265[124:124];
    assign _2775 = _2768 & _2774;
    assign _2778 = _2775 & _2777;
    assign _2806 = _2778 ? _2771 : _290;
    assign _2804 = _2798 ? _290 : _2791;
    assign _2807 = _2804 + _2806;
    assign _2821 = _2807 + _2820;
    assign _6298 = _287 ? _2821 : _2791;
    assign _6304 = _278 ? _6303 : _6298;
    assign _133 = _6304;
    always @(posedge _272) begin
        if (_270)
            _2791 <= _290;
        else
            _2791 <= _133;
    end
    assign _2793 = _2791 == _290;
    assign _2794 = ~ _2793;
    assign _2788 = _265[125:125];
    assign _2795 = _2788 & _2794;
    assign _2798 = _2795 & _2797;
    assign _2826 = _2798 ? _2791 : _290;
    assign _2824 = _2818 ? _290 : _2811;
    assign _2827 = _2824 + _2826;
    assign _2841 = _2827 + _2840;
    assign _6305 = _287 ? _2841 : _2811;
    assign _6311 = _278 ? _6310 : _6305;
    assign _134 = _6311;
    always @(posedge _272) begin
        if (_270)
            _2811 <= _290;
        else
            _2811 <= _134;
    end
    assign _2813 = _2811 == _290;
    assign _2814 = ~ _2813;
    assign _2808 = _265[126:126];
    assign _2815 = _2808 & _2814;
    assign _2818 = _2815 & _2817;
    assign _2846 = _2818 ? _2811 : _290;
    assign _2844 = _2838 ? _290 : _2831;
    assign _2847 = _2844 + _2846;
    assign _2861 = _2847 + _2860;
    assign _6312 = _287 ? _2861 : _2831;
    assign _6318 = _278 ? _6317 : _6312;
    assign _135 = _6318;
    always @(posedge _272) begin
        if (_270)
            _2831 <= _290;
        else
            _2831 <= _135;
    end
    assign _2833 = _2831 == _290;
    assign _2834 = ~ _2833;
    assign _2828 = _265[127:127];
    assign _2835 = _2828 & _2834;
    assign _2838 = _2835 & _2837;
    assign _2866 = _2838 ? _2831 : _290;
    assign _2864 = _2858 ? _290 : _2851;
    assign _2867 = _2864 + _2866;
    assign _2881 = _2867 + _2880;
    assign _6319 = _287 ? _2881 : _2851;
    assign _6325 = _278 ? _6324 : _6319;
    assign _136 = _6325;
    always @(posedge _272) begin
        if (_270)
            _2851 <= _290;
        else
            _2851 <= _136;
    end
    assign _2853 = _2851 == _290;
    assign _2854 = ~ _2853;
    assign _2848 = _265[128:128];
    assign _2855 = _2848 & _2854;
    assign _2858 = _2855 & _2857;
    assign _2886 = _2858 ? _2851 : _290;
    assign _2884 = _2878 ? _290 : _2871;
    assign _2887 = _2884 + _2886;
    assign _2901 = _2887 + _2900;
    assign _6326 = _287 ? _2901 : _2871;
    assign _6332 = _278 ? _6331 : _6326;
    assign _137 = _6332;
    always @(posedge _272) begin
        if (_270)
            _2871 <= _290;
        else
            _2871 <= _137;
    end
    assign _2873 = _2871 == _290;
    assign _2874 = ~ _2873;
    assign _2868 = _265[129:129];
    assign _2875 = _2868 & _2874;
    assign _2878 = _2875 & _2877;
    assign _2906 = _2878 ? _2871 : _290;
    assign _2904 = _2898 ? _290 : _2891;
    assign _2907 = _2904 + _2906;
    assign _2921 = _2907 + _2920;
    assign _6333 = _287 ? _2921 : _2891;
    assign _6339 = _278 ? _6338 : _6333;
    assign _138 = _6339;
    always @(posedge _272) begin
        if (_270)
            _2891 <= _290;
        else
            _2891 <= _138;
    end
    assign _2893 = _2891 == _290;
    assign _2894 = ~ _2893;
    assign _2888 = _265[130:130];
    assign _2895 = _2888 & _2894;
    assign _2898 = _2895 & _2897;
    assign _2926 = _2898 ? _2891 : _290;
    assign _2924 = _2918 ? _290 : _2911;
    assign _2927 = _2924 + _2926;
    assign _2941 = _2927 + _2940;
    assign _6340 = _287 ? _2941 : _2911;
    assign _6346 = _278 ? _6345 : _6340;
    assign _139 = _6346;
    always @(posedge _272) begin
        if (_270)
            _2911 <= _290;
        else
            _2911 <= _139;
    end
    assign _2913 = _2911 == _290;
    assign _2914 = ~ _2913;
    assign _2908 = _265[131:131];
    assign _2915 = _2908 & _2914;
    assign _2918 = _2915 & _2917;
    assign _2946 = _2918 ? _2911 : _290;
    assign _2944 = _2938 ? _290 : _2931;
    assign _2947 = _2944 + _2946;
    assign _2961 = _2947 + _2960;
    assign _6347 = _287 ? _2961 : _2931;
    assign _6353 = _278 ? _6352 : _6347;
    assign _140 = _6353;
    always @(posedge _272) begin
        if (_270)
            _2931 <= _290;
        else
            _2931 <= _140;
    end
    assign _2933 = _2931 == _290;
    assign _2934 = ~ _2933;
    assign _2928 = _265[132:132];
    assign _2935 = _2928 & _2934;
    assign _2938 = _2935 & _2937;
    assign _2966 = _2938 ? _2931 : _290;
    assign _2964 = _2958 ? _290 : _2951;
    assign _2967 = _2964 + _2966;
    assign _2981 = _2967 + _2980;
    assign _6354 = _287 ? _2981 : _2951;
    assign _6360 = _278 ? _6359 : _6354;
    assign _141 = _6360;
    always @(posedge _272) begin
        if (_270)
            _2951 <= _290;
        else
            _2951 <= _141;
    end
    assign _2953 = _2951 == _290;
    assign _2954 = ~ _2953;
    assign _2948 = _265[133:133];
    assign _2955 = _2948 & _2954;
    assign _2958 = _2955 & _2957;
    assign _2986 = _2958 ? _2951 : _290;
    assign _2984 = _2978 ? _290 : _2971;
    assign _2987 = _2984 + _2986;
    assign _3001 = _2987 + _3000;
    assign _6361 = _287 ? _3001 : _2971;
    assign _6367 = _278 ? _6366 : _6361;
    assign _142 = _6367;
    always @(posedge _272) begin
        if (_270)
            _2971 <= _290;
        else
            _2971 <= _142;
    end
    assign _2973 = _2971 == _290;
    assign _2974 = ~ _2973;
    assign _2968 = _265[134:134];
    assign _2975 = _2968 & _2974;
    assign _2978 = _2975 & _2977;
    assign _3006 = _2978 ? _2971 : _290;
    assign _3004 = _2998 ? _290 : _2991;
    assign _3007 = _3004 + _3006;
    assign _3021 = _3007 + _3020;
    assign _6368 = _287 ? _3021 : _2991;
    assign _6374 = _278 ? _6373 : _6368;
    assign _143 = _6374;
    always @(posedge _272) begin
        if (_270)
            _2991 <= _290;
        else
            _2991 <= _143;
    end
    assign _2993 = _2991 == _290;
    assign _2994 = ~ _2993;
    assign _2988 = _265[135:135];
    assign _2995 = _2988 & _2994;
    assign _2998 = _2995 & _2997;
    assign _3026 = _2998 ? _2991 : _290;
    assign _3024 = _3018 ? _290 : _3011;
    assign _3027 = _3024 + _3026;
    assign _3041 = _3027 + _3040;
    assign _6375 = _287 ? _3041 : _3011;
    assign _6381 = _278 ? _6380 : _6375;
    assign _144 = _6381;
    always @(posedge _272) begin
        if (_270)
            _3011 <= _290;
        else
            _3011 <= _144;
    end
    assign _3013 = _3011 == _290;
    assign _3014 = ~ _3013;
    assign _3008 = _265[136:136];
    assign _3015 = _3008 & _3014;
    assign _3018 = _3015 & _3017;
    assign _3046 = _3018 ? _3011 : _290;
    assign _3044 = _3038 ? _290 : _3031;
    assign _3047 = _3044 + _3046;
    assign _3061 = _3047 + _3060;
    assign _6382 = _287 ? _3061 : _3031;
    assign _6388 = _278 ? _6387 : _6382;
    assign _145 = _6388;
    always @(posedge _272) begin
        if (_270)
            _3031 <= _290;
        else
            _3031 <= _145;
    end
    assign _3033 = _3031 == _290;
    assign _3034 = ~ _3033;
    assign _3028 = _265[137:137];
    assign _3035 = _3028 & _3034;
    assign _3038 = _3035 & _3037;
    assign _3066 = _3038 ? _3031 : _290;
    assign _3064 = _3058 ? _290 : _3051;
    assign _3067 = _3064 + _3066;
    assign _3081 = _3067 + _3080;
    assign _6389 = _287 ? _3081 : _3051;
    assign _6395 = _278 ? _6394 : _6389;
    assign _146 = _6395;
    always @(posedge _272) begin
        if (_270)
            _3051 <= _290;
        else
            _3051 <= _146;
    end
    assign _3053 = _3051 == _290;
    assign _3054 = ~ _3053;
    assign _3048 = _265[138:138];
    assign _3055 = _3048 & _3054;
    assign _3058 = _3055 & _3057;
    assign _3086 = _3058 ? _3051 : _290;
    assign _3084 = _3078 ? _290 : _3071;
    assign _3087 = _3084 + _3086;
    assign _3101 = _3087 + _3100;
    assign _6396 = _287 ? _3101 : _3071;
    assign _6402 = _278 ? _6401 : _6396;
    assign _147 = _6402;
    always @(posedge _272) begin
        if (_270)
            _3071 <= _290;
        else
            _3071 <= _147;
    end
    assign _3073 = _3071 == _290;
    assign _3074 = ~ _3073;
    assign _3068 = _265[139:139];
    assign _3075 = _3068 & _3074;
    assign _3078 = _3075 & _3077;
    assign _3106 = _3078 ? _3071 : _290;
    assign _3104 = _3098 ? _290 : _3091;
    assign _3107 = _3104 + _3106;
    assign _3121 = _3107 + _3120;
    assign _6403 = _287 ? _3121 : _3091;
    assign _6409 = _278 ? _6408 : _6403;
    assign _148 = _6409;
    always @(posedge _272) begin
        if (_270)
            _3091 <= _290;
        else
            _3091 <= _148;
    end
    assign _3093 = _3091 == _290;
    assign _3094 = ~ _3093;
    assign _3088 = _265[140:140];
    assign _3095 = _3088 & _3094;
    assign _3098 = _3095 & _3097;
    assign _3126 = _3098 ? _3091 : _290;
    assign _3124 = _3118 ? _290 : _3111;
    assign _3127 = _3124 + _3126;
    assign _3141 = _3127 + _3140;
    assign _6410 = _287 ? _3141 : _3111;
    assign _6416 = _278 ? _6415 : _6410;
    assign _149 = _6416;
    always @(posedge _272) begin
        if (_270)
            _3111 <= _290;
        else
            _3111 <= _149;
    end
    assign _3113 = _3111 == _290;
    assign _3114 = ~ _3113;
    assign _3108 = _265[141:141];
    assign _3115 = _3108 & _3114;
    assign _3118 = _3115 & _3117;
    assign _3146 = _3118 ? _3111 : _290;
    assign _3144 = _3138 ? _290 : _3131;
    assign _3147 = _3144 + _3146;
    assign _3161 = _3147 + _3160;
    assign _6417 = _287 ? _3161 : _3131;
    assign _6423 = _278 ? _6422 : _6417;
    assign _150 = _6423;
    always @(posedge _272) begin
        if (_270)
            _3131 <= _290;
        else
            _3131 <= _150;
    end
    assign _3133 = _3131 == _290;
    assign _3134 = ~ _3133;
    assign _3128 = _265[142:142];
    assign _3135 = _3128 & _3134;
    assign _3138 = _3135 & _3137;
    assign _3166 = _3138 ? _3131 : _290;
    assign _3164 = _3158 ? _290 : _3151;
    assign _3167 = _3164 + _3166;
    assign _3181 = _3167 + _3180;
    assign _6424 = _287 ? _3181 : _3151;
    assign _6430 = _278 ? _6429 : _6424;
    assign _151 = _6430;
    always @(posedge _272) begin
        if (_270)
            _3151 <= _290;
        else
            _3151 <= _151;
    end
    assign _3153 = _3151 == _290;
    assign _3154 = ~ _3153;
    assign _3148 = _265[143:143];
    assign _3155 = _3148 & _3154;
    assign _3158 = _3155 & _3157;
    assign _3186 = _3158 ? _3151 : _290;
    assign _3184 = _3178 ? _290 : _3171;
    assign _3187 = _3184 + _3186;
    assign _3201 = _3187 + _3200;
    assign _6431 = _287 ? _3201 : _3171;
    assign _6437 = _278 ? _6436 : _6431;
    assign _152 = _6437;
    always @(posedge _272) begin
        if (_270)
            _3171 <= _290;
        else
            _3171 <= _152;
    end
    assign _3173 = _3171 == _290;
    assign _3174 = ~ _3173;
    assign _3168 = _265[144:144];
    assign _3175 = _3168 & _3174;
    assign _3178 = _3175 & _3177;
    assign _3206 = _3178 ? _3171 : _290;
    assign _3204 = _3198 ? _290 : _3191;
    assign _3207 = _3204 + _3206;
    assign _3221 = _3207 + _3220;
    assign _6438 = _287 ? _3221 : _3191;
    assign _6444 = _278 ? _6443 : _6438;
    assign _153 = _6444;
    always @(posedge _272) begin
        if (_270)
            _3191 <= _290;
        else
            _3191 <= _153;
    end
    assign _3193 = _3191 == _290;
    assign _3194 = ~ _3193;
    assign _3188 = _265[145:145];
    assign _3195 = _3188 & _3194;
    assign _3198 = _3195 & _3197;
    assign _3226 = _3198 ? _3191 : _290;
    assign _3224 = _3218 ? _290 : _3211;
    assign _3227 = _3224 + _3226;
    assign _3241 = _3227 + _3240;
    assign _6445 = _287 ? _3241 : _3211;
    assign _6451 = _278 ? _6450 : _6445;
    assign _154 = _6451;
    always @(posedge _272) begin
        if (_270)
            _3211 <= _290;
        else
            _3211 <= _154;
    end
    assign _3213 = _3211 == _290;
    assign _3214 = ~ _3213;
    assign _3208 = _265[146:146];
    assign _3215 = _3208 & _3214;
    assign _3218 = _3215 & _3217;
    assign _3246 = _3218 ? _3211 : _290;
    assign _3244 = _3238 ? _290 : _3231;
    assign _3247 = _3244 + _3246;
    assign _3261 = _3247 + _3260;
    assign _6452 = _287 ? _3261 : _3231;
    assign _6458 = _278 ? _6457 : _6452;
    assign _155 = _6458;
    always @(posedge _272) begin
        if (_270)
            _3231 <= _290;
        else
            _3231 <= _155;
    end
    assign _3233 = _3231 == _290;
    assign _3234 = ~ _3233;
    assign _3228 = _265[147:147];
    assign _3235 = _3228 & _3234;
    assign _3238 = _3235 & _3237;
    assign _3266 = _3238 ? _3231 : _290;
    assign _3264 = _3258 ? _290 : _3251;
    assign _3267 = _3264 + _3266;
    assign _3281 = _3267 + _3280;
    assign _6459 = _287 ? _3281 : _3251;
    assign _6465 = _278 ? _6464 : _6459;
    assign _156 = _6465;
    always @(posedge _272) begin
        if (_270)
            _3251 <= _290;
        else
            _3251 <= _156;
    end
    assign _3253 = _3251 == _290;
    assign _3254 = ~ _3253;
    assign _3248 = _265[148:148];
    assign _3255 = _3248 & _3254;
    assign _3258 = _3255 & _3257;
    assign _3286 = _3258 ? _3251 : _290;
    assign _3284 = _3278 ? _290 : _3271;
    assign _3287 = _3284 + _3286;
    assign _3301 = _3287 + _3300;
    assign _6466 = _287 ? _3301 : _3271;
    assign _6472 = _278 ? _6471 : _6466;
    assign _157 = _6472;
    always @(posedge _272) begin
        if (_270)
            _3271 <= _290;
        else
            _3271 <= _157;
    end
    assign _3273 = _3271 == _290;
    assign _3274 = ~ _3273;
    assign _3268 = _265[149:149];
    assign _3275 = _3268 & _3274;
    assign _3278 = _3275 & _3277;
    assign _3306 = _3278 ? _3271 : _290;
    assign _3304 = _3298 ? _290 : _3291;
    assign _3307 = _3304 + _3306;
    assign _3321 = _3307 + _3320;
    assign _6473 = _287 ? _3321 : _3291;
    assign _6479 = _278 ? _6478 : _6473;
    assign _158 = _6479;
    always @(posedge _272) begin
        if (_270)
            _3291 <= _290;
        else
            _3291 <= _158;
    end
    assign _3293 = _3291 == _290;
    assign _3294 = ~ _3293;
    assign _3288 = _265[150:150];
    assign _3295 = _3288 & _3294;
    assign _3298 = _3295 & _3297;
    assign _3326 = _3298 ? _3291 : _290;
    assign _3324 = _3318 ? _290 : _3311;
    assign _3327 = _3324 + _3326;
    assign _3341 = _3327 + _3340;
    assign _6480 = _287 ? _3341 : _3311;
    assign _6486 = _278 ? _6485 : _6480;
    assign _159 = _6486;
    always @(posedge _272) begin
        if (_270)
            _3311 <= _290;
        else
            _3311 <= _159;
    end
    assign _3313 = _3311 == _290;
    assign _3314 = ~ _3313;
    assign _3308 = _265[151:151];
    assign _3315 = _3308 & _3314;
    assign _3318 = _3315 & _3317;
    assign _3346 = _3318 ? _3311 : _290;
    assign _3344 = _3338 ? _290 : _3331;
    assign _3347 = _3344 + _3346;
    assign _3361 = _3347 + _3360;
    assign _6487 = _287 ? _3361 : _3331;
    assign _6493 = _278 ? _6492 : _6487;
    assign _160 = _6493;
    always @(posedge _272) begin
        if (_270)
            _3331 <= _290;
        else
            _3331 <= _160;
    end
    assign _3333 = _3331 == _290;
    assign _3334 = ~ _3333;
    assign _3328 = _265[152:152];
    assign _3335 = _3328 & _3334;
    assign _3338 = _3335 & _3337;
    assign _3366 = _3338 ? _3331 : _290;
    assign _3364 = _3358 ? _290 : _3351;
    assign _3367 = _3364 + _3366;
    assign _3381 = _3367 + _3380;
    assign _6494 = _287 ? _3381 : _3351;
    assign _6500 = _278 ? _6499 : _6494;
    assign _161 = _6500;
    always @(posedge _272) begin
        if (_270)
            _3351 <= _290;
        else
            _3351 <= _161;
    end
    assign _3353 = _3351 == _290;
    assign _3354 = ~ _3353;
    assign _3348 = _265[153:153];
    assign _3355 = _3348 & _3354;
    assign _3358 = _3355 & _3357;
    assign _3386 = _3358 ? _3351 : _290;
    assign _3384 = _3378 ? _290 : _3371;
    assign _3387 = _3384 + _3386;
    assign _3401 = _3387 + _3400;
    assign _6501 = _287 ? _3401 : _3371;
    assign _6507 = _278 ? _6506 : _6501;
    assign _162 = _6507;
    always @(posedge _272) begin
        if (_270)
            _3371 <= _290;
        else
            _3371 <= _162;
    end
    assign _3373 = _3371 == _290;
    assign _3374 = ~ _3373;
    assign _3368 = _265[154:154];
    assign _3375 = _3368 & _3374;
    assign _3378 = _3375 & _3377;
    assign _3406 = _3378 ? _3371 : _290;
    assign _3404 = _3398 ? _290 : _3391;
    assign _3407 = _3404 + _3406;
    assign _3421 = _3407 + _3420;
    assign _6508 = _287 ? _3421 : _3391;
    assign _6514 = _278 ? _6513 : _6508;
    assign _163 = _6514;
    always @(posedge _272) begin
        if (_270)
            _3391 <= _290;
        else
            _3391 <= _163;
    end
    assign _3393 = _3391 == _290;
    assign _3394 = ~ _3393;
    assign _3388 = _265[155:155];
    assign _3395 = _3388 & _3394;
    assign _3398 = _3395 & _3397;
    assign _3426 = _3398 ? _3391 : _290;
    assign _3424 = _3418 ? _290 : _3411;
    assign _3427 = _3424 + _3426;
    assign _3441 = _3427 + _3440;
    assign _6515 = _287 ? _3441 : _3411;
    assign _6521 = _278 ? _6520 : _6515;
    assign _164 = _6521;
    always @(posedge _272) begin
        if (_270)
            _3411 <= _290;
        else
            _3411 <= _164;
    end
    assign _3413 = _3411 == _290;
    assign _3414 = ~ _3413;
    assign _3408 = _265[156:156];
    assign _3415 = _3408 & _3414;
    assign _3418 = _3415 & _3417;
    assign _3446 = _3418 ? _3411 : _290;
    assign _3444 = _3438 ? _290 : _3431;
    assign _3447 = _3444 + _3446;
    assign _3461 = _3447 + _3460;
    assign _6522 = _287 ? _3461 : _3431;
    assign _6528 = _278 ? _6527 : _6522;
    assign _165 = _6528;
    always @(posedge _272) begin
        if (_270)
            _3431 <= _290;
        else
            _3431 <= _165;
    end
    assign _3433 = _3431 == _290;
    assign _3434 = ~ _3433;
    assign _3428 = _265[157:157];
    assign _3435 = _3428 & _3434;
    assign _3438 = _3435 & _3437;
    assign _3466 = _3438 ? _3431 : _290;
    assign _3464 = _3458 ? _290 : _3451;
    assign _3467 = _3464 + _3466;
    assign _3481 = _3467 + _3480;
    assign _6529 = _287 ? _3481 : _3451;
    assign _6535 = _278 ? _6534 : _6529;
    assign _166 = _6535;
    always @(posedge _272) begin
        if (_270)
            _3451 <= _290;
        else
            _3451 <= _166;
    end
    assign _3453 = _3451 == _290;
    assign _3454 = ~ _3453;
    assign _3448 = _265[158:158];
    assign _3455 = _3448 & _3454;
    assign _3458 = _3455 & _3457;
    assign _3486 = _3458 ? _3451 : _290;
    assign _3484 = _3478 ? _290 : _3471;
    assign _3487 = _3484 + _3486;
    assign _3501 = _3487 + _3500;
    assign _6536 = _287 ? _3501 : _3471;
    assign _6542 = _278 ? _6541 : _6536;
    assign _167 = _6542;
    always @(posedge _272) begin
        if (_270)
            _3471 <= _290;
        else
            _3471 <= _167;
    end
    assign _3473 = _3471 == _290;
    assign _3474 = ~ _3473;
    assign _3468 = _265[159:159];
    assign _3475 = _3468 & _3474;
    assign _3478 = _3475 & _3477;
    assign _3506 = _3478 ? _3471 : _290;
    assign _3504 = _3498 ? _290 : _3491;
    assign _3507 = _3504 + _3506;
    assign _3521 = _3507 + _3520;
    assign _6543 = _287 ? _3521 : _3491;
    assign _6549 = _278 ? _6548 : _6543;
    assign _168 = _6549;
    always @(posedge _272) begin
        if (_270)
            _3491 <= _290;
        else
            _3491 <= _168;
    end
    assign _3493 = _3491 == _290;
    assign _3494 = ~ _3493;
    assign _3488 = _265[160:160];
    assign _3495 = _3488 & _3494;
    assign _3498 = _3495 & _3497;
    assign _3526 = _3498 ? _3491 : _290;
    assign _3524 = _3518 ? _290 : _3511;
    assign _3527 = _3524 + _3526;
    assign _3541 = _3527 + _3540;
    assign _6550 = _287 ? _3541 : _3511;
    assign _6556 = _278 ? _6555 : _6550;
    assign _169 = _6556;
    always @(posedge _272) begin
        if (_270)
            _3511 <= _290;
        else
            _3511 <= _169;
    end
    assign _3513 = _3511 == _290;
    assign _3514 = ~ _3513;
    assign _3508 = _265[161:161];
    assign _3515 = _3508 & _3514;
    assign _3518 = _3515 & _3517;
    assign _3546 = _3518 ? _3511 : _290;
    assign _3544 = _3538 ? _290 : _3531;
    assign _3547 = _3544 + _3546;
    assign _3561 = _3547 + _3560;
    assign _6557 = _287 ? _3561 : _3531;
    assign _6563 = _278 ? _6562 : _6557;
    assign _170 = _6563;
    always @(posedge _272) begin
        if (_270)
            _3531 <= _290;
        else
            _3531 <= _170;
    end
    assign _3533 = _3531 == _290;
    assign _3534 = ~ _3533;
    assign _3528 = _265[162:162];
    assign _3535 = _3528 & _3534;
    assign _3538 = _3535 & _3537;
    assign _3566 = _3538 ? _3531 : _290;
    assign _3564 = _3558 ? _290 : _3551;
    assign _3567 = _3564 + _3566;
    assign _3581 = _3567 + _3580;
    assign _6564 = _287 ? _3581 : _3551;
    assign _6570 = _278 ? _6569 : _6564;
    assign _171 = _6570;
    always @(posedge _272) begin
        if (_270)
            _3551 <= _290;
        else
            _3551 <= _171;
    end
    assign _3553 = _3551 == _290;
    assign _3554 = ~ _3553;
    assign _3548 = _265[163:163];
    assign _3555 = _3548 & _3554;
    assign _3558 = _3555 & _3557;
    assign _3586 = _3558 ? _3551 : _290;
    assign _3584 = _3578 ? _290 : _3571;
    assign _3587 = _3584 + _3586;
    assign _3601 = _3587 + _3600;
    assign _6571 = _287 ? _3601 : _3571;
    assign _6577 = _278 ? _6576 : _6571;
    assign _172 = _6577;
    always @(posedge _272) begin
        if (_270)
            _3571 <= _290;
        else
            _3571 <= _172;
    end
    assign _3573 = _3571 == _290;
    assign _3574 = ~ _3573;
    assign _3568 = _265[164:164];
    assign _3575 = _3568 & _3574;
    assign _3578 = _3575 & _3577;
    assign _3606 = _3578 ? _3571 : _290;
    assign _3604 = _3598 ? _290 : _3591;
    assign _3607 = _3604 + _3606;
    assign _3621 = _3607 + _3620;
    assign _6578 = _287 ? _3621 : _3591;
    assign _6584 = _278 ? _6583 : _6578;
    assign _173 = _6584;
    always @(posedge _272) begin
        if (_270)
            _3591 <= _290;
        else
            _3591 <= _173;
    end
    assign _3593 = _3591 == _290;
    assign _3594 = ~ _3593;
    assign _3588 = _265[165:165];
    assign _3595 = _3588 & _3594;
    assign _3598 = _3595 & _3597;
    assign _3626 = _3598 ? _3591 : _290;
    assign _3624 = _3618 ? _290 : _3611;
    assign _3627 = _3624 + _3626;
    assign _3641 = _3627 + _3640;
    assign _6585 = _287 ? _3641 : _3611;
    assign _6591 = _278 ? _6590 : _6585;
    assign _174 = _6591;
    always @(posedge _272) begin
        if (_270)
            _3611 <= _290;
        else
            _3611 <= _174;
    end
    assign _3613 = _3611 == _290;
    assign _3614 = ~ _3613;
    assign _3608 = _265[166:166];
    assign _3615 = _3608 & _3614;
    assign _3618 = _3615 & _3617;
    assign _3646 = _3618 ? _3611 : _290;
    assign _3644 = _3638 ? _290 : _3631;
    assign _3647 = _3644 + _3646;
    assign _3661 = _3647 + _3660;
    assign _6592 = _287 ? _3661 : _3631;
    assign _6598 = _278 ? _6597 : _6592;
    assign _175 = _6598;
    always @(posedge _272) begin
        if (_270)
            _3631 <= _290;
        else
            _3631 <= _175;
    end
    assign _3633 = _3631 == _290;
    assign _3634 = ~ _3633;
    assign _3628 = _265[167:167];
    assign _3635 = _3628 & _3634;
    assign _3638 = _3635 & _3637;
    assign _3666 = _3638 ? _3631 : _290;
    assign _3664 = _3658 ? _290 : _3651;
    assign _3667 = _3664 + _3666;
    assign _3681 = _3667 + _3680;
    assign _6599 = _287 ? _3681 : _3651;
    assign _6605 = _278 ? _6604 : _6599;
    assign _176 = _6605;
    always @(posedge _272) begin
        if (_270)
            _3651 <= _290;
        else
            _3651 <= _176;
    end
    assign _3653 = _3651 == _290;
    assign _3654 = ~ _3653;
    assign _3648 = _265[168:168];
    assign _3655 = _3648 & _3654;
    assign _3658 = _3655 & _3657;
    assign _3686 = _3658 ? _3651 : _290;
    assign _3684 = _3678 ? _290 : _3671;
    assign _3687 = _3684 + _3686;
    assign _3701 = _3687 + _3700;
    assign _6606 = _287 ? _3701 : _3671;
    assign _6612 = _278 ? _6611 : _6606;
    assign _177 = _6612;
    always @(posedge _272) begin
        if (_270)
            _3671 <= _290;
        else
            _3671 <= _177;
    end
    assign _3673 = _3671 == _290;
    assign _3674 = ~ _3673;
    assign _3668 = _265[169:169];
    assign _3675 = _3668 & _3674;
    assign _3678 = _3675 & _3677;
    assign _3706 = _3678 ? _3671 : _290;
    assign _3704 = _3698 ? _290 : _3691;
    assign _3707 = _3704 + _3706;
    assign _3721 = _3707 + _3720;
    assign _6613 = _287 ? _3721 : _3691;
    assign _6619 = _278 ? _6618 : _6613;
    assign _178 = _6619;
    always @(posedge _272) begin
        if (_270)
            _3691 <= _290;
        else
            _3691 <= _178;
    end
    assign _3693 = _3691 == _290;
    assign _3694 = ~ _3693;
    assign _3688 = _265[170:170];
    assign _3695 = _3688 & _3694;
    assign _3698 = _3695 & _3697;
    assign _3726 = _3698 ? _3691 : _290;
    assign _3724 = _3718 ? _290 : _3711;
    assign _3727 = _3724 + _3726;
    assign _3741 = _3727 + _3740;
    assign _6620 = _287 ? _3741 : _3711;
    assign _6626 = _278 ? _6625 : _6620;
    assign _179 = _6626;
    always @(posedge _272) begin
        if (_270)
            _3711 <= _290;
        else
            _3711 <= _179;
    end
    assign _3713 = _3711 == _290;
    assign _3714 = ~ _3713;
    assign _3708 = _265[171:171];
    assign _3715 = _3708 & _3714;
    assign _3718 = _3715 & _3717;
    assign _3746 = _3718 ? _3711 : _290;
    assign _3744 = _3738 ? _290 : _3731;
    assign _3747 = _3744 + _3746;
    assign _3761 = _3747 + _3760;
    assign _6627 = _287 ? _3761 : _3731;
    assign _6633 = _278 ? _6632 : _6627;
    assign _180 = _6633;
    always @(posedge _272) begin
        if (_270)
            _3731 <= _290;
        else
            _3731 <= _180;
    end
    assign _3733 = _3731 == _290;
    assign _3734 = ~ _3733;
    assign _3728 = _265[172:172];
    assign _3735 = _3728 & _3734;
    assign _3738 = _3735 & _3737;
    assign _3766 = _3738 ? _3731 : _290;
    assign _3764 = _3758 ? _290 : _3751;
    assign _3767 = _3764 + _3766;
    assign _3781 = _3767 + _3780;
    assign _6634 = _287 ? _3781 : _3751;
    assign _6640 = _278 ? _6639 : _6634;
    assign _181 = _6640;
    always @(posedge _272) begin
        if (_270)
            _3751 <= _290;
        else
            _3751 <= _181;
    end
    assign _3753 = _3751 == _290;
    assign _3754 = ~ _3753;
    assign _3748 = _265[173:173];
    assign _3755 = _3748 & _3754;
    assign _3758 = _3755 & _3757;
    assign _3786 = _3758 ? _3751 : _290;
    assign _3784 = _3778 ? _290 : _3771;
    assign _3787 = _3784 + _3786;
    assign _3801 = _3787 + _3800;
    assign _6641 = _287 ? _3801 : _3771;
    assign _6647 = _278 ? _6646 : _6641;
    assign _182 = _6647;
    always @(posedge _272) begin
        if (_270)
            _3771 <= _290;
        else
            _3771 <= _182;
    end
    assign _3773 = _3771 == _290;
    assign _3774 = ~ _3773;
    assign _3768 = _265[174:174];
    assign _3775 = _3768 & _3774;
    assign _3778 = _3775 & _3777;
    assign _3806 = _3778 ? _3771 : _290;
    assign _3804 = _3798 ? _290 : _3791;
    assign _3807 = _3804 + _3806;
    assign _3821 = _3807 + _3820;
    assign _6648 = _287 ? _3821 : _3791;
    assign _6654 = _278 ? _6653 : _6648;
    assign _183 = _6654;
    always @(posedge _272) begin
        if (_270)
            _3791 <= _290;
        else
            _3791 <= _183;
    end
    assign _3793 = _3791 == _290;
    assign _3794 = ~ _3793;
    assign _3788 = _265[175:175];
    assign _3795 = _3788 & _3794;
    assign _3798 = _3795 & _3797;
    assign _3826 = _3798 ? _3791 : _290;
    assign _3824 = _3818 ? _290 : _3811;
    assign _3827 = _3824 + _3826;
    assign _3841 = _3827 + _3840;
    assign _6655 = _287 ? _3841 : _3811;
    assign _6661 = _278 ? _6660 : _6655;
    assign _184 = _6661;
    always @(posedge _272) begin
        if (_270)
            _3811 <= _290;
        else
            _3811 <= _184;
    end
    assign _3813 = _3811 == _290;
    assign _3814 = ~ _3813;
    assign _3808 = _265[176:176];
    assign _3815 = _3808 & _3814;
    assign _3818 = _3815 & _3817;
    assign _3846 = _3818 ? _3811 : _290;
    assign _3844 = _3838 ? _290 : _3831;
    assign _3847 = _3844 + _3846;
    assign _3861 = _3847 + _3860;
    assign _6662 = _287 ? _3861 : _3831;
    assign _6668 = _278 ? _6667 : _6662;
    assign _185 = _6668;
    always @(posedge _272) begin
        if (_270)
            _3831 <= _290;
        else
            _3831 <= _185;
    end
    assign _3833 = _3831 == _290;
    assign _3834 = ~ _3833;
    assign _3828 = _265[177:177];
    assign _3835 = _3828 & _3834;
    assign _3838 = _3835 & _3837;
    assign _3866 = _3838 ? _3831 : _290;
    assign _3864 = _3858 ? _290 : _3851;
    assign _3867 = _3864 + _3866;
    assign _3881 = _3867 + _3880;
    assign _6669 = _287 ? _3881 : _3851;
    assign _6675 = _278 ? _6674 : _6669;
    assign _186 = _6675;
    always @(posedge _272) begin
        if (_270)
            _3851 <= _290;
        else
            _3851 <= _186;
    end
    assign _3853 = _3851 == _290;
    assign _3854 = ~ _3853;
    assign _3848 = _265[178:178];
    assign _3855 = _3848 & _3854;
    assign _3858 = _3855 & _3857;
    assign _3886 = _3858 ? _3851 : _290;
    assign _3884 = _3878 ? _290 : _3871;
    assign _3887 = _3884 + _3886;
    assign _3901 = _3887 + _3900;
    assign _6676 = _287 ? _3901 : _3871;
    assign _6682 = _278 ? _6681 : _6676;
    assign _187 = _6682;
    always @(posedge _272) begin
        if (_270)
            _3871 <= _290;
        else
            _3871 <= _187;
    end
    assign _3873 = _3871 == _290;
    assign _3874 = ~ _3873;
    assign _3868 = _265[179:179];
    assign _3875 = _3868 & _3874;
    assign _3878 = _3875 & _3877;
    assign _3906 = _3878 ? _3871 : _290;
    assign _3904 = _3898 ? _290 : _3891;
    assign _3907 = _3904 + _3906;
    assign _3921 = _3907 + _3920;
    assign _6683 = _287 ? _3921 : _3891;
    assign _6689 = _278 ? _6688 : _6683;
    assign _188 = _6689;
    always @(posedge _272) begin
        if (_270)
            _3891 <= _290;
        else
            _3891 <= _188;
    end
    assign _3893 = _3891 == _290;
    assign _3894 = ~ _3893;
    assign _3888 = _265[180:180];
    assign _3895 = _3888 & _3894;
    assign _3898 = _3895 & _3897;
    assign _3926 = _3898 ? _3891 : _290;
    assign _3924 = _3918 ? _290 : _3911;
    assign _3927 = _3924 + _3926;
    assign _3941 = _3927 + _3940;
    assign _6690 = _287 ? _3941 : _3911;
    assign _6696 = _278 ? _6695 : _6690;
    assign _189 = _6696;
    always @(posedge _272) begin
        if (_270)
            _3911 <= _290;
        else
            _3911 <= _189;
    end
    assign _3913 = _3911 == _290;
    assign _3914 = ~ _3913;
    assign _3908 = _265[181:181];
    assign _3915 = _3908 & _3914;
    assign _3918 = _3915 & _3917;
    assign _3946 = _3918 ? _3911 : _290;
    assign _3944 = _3938 ? _290 : _3931;
    assign _3947 = _3944 + _3946;
    assign _3961 = _3947 + _3960;
    assign _6697 = _287 ? _3961 : _3931;
    assign _6703 = _278 ? _6702 : _6697;
    assign _190 = _6703;
    always @(posedge _272) begin
        if (_270)
            _3931 <= _290;
        else
            _3931 <= _190;
    end
    assign _3933 = _3931 == _290;
    assign _3934 = ~ _3933;
    assign _3928 = _265[182:182];
    assign _3935 = _3928 & _3934;
    assign _3938 = _3935 & _3937;
    assign _3966 = _3938 ? _3931 : _290;
    assign _3964 = _3958 ? _290 : _3951;
    assign _3967 = _3964 + _3966;
    assign _3981 = _3967 + _3980;
    assign _6704 = _287 ? _3981 : _3951;
    assign _6710 = _278 ? _6709 : _6704;
    assign _191 = _6710;
    always @(posedge _272) begin
        if (_270)
            _3951 <= _290;
        else
            _3951 <= _191;
    end
    assign _3953 = _3951 == _290;
    assign _3954 = ~ _3953;
    assign _3948 = _265[183:183];
    assign _3955 = _3948 & _3954;
    assign _3958 = _3955 & _3957;
    assign _3986 = _3958 ? _3951 : _290;
    assign _3984 = _3978 ? _290 : _3971;
    assign _3987 = _3984 + _3986;
    assign _4001 = _3987 + _4000;
    assign _6711 = _287 ? _4001 : _3971;
    assign _6717 = _278 ? _6716 : _6711;
    assign _192 = _6717;
    always @(posedge _272) begin
        if (_270)
            _3971 <= _290;
        else
            _3971 <= _192;
    end
    assign _3973 = _3971 == _290;
    assign _3974 = ~ _3973;
    assign _3968 = _265[184:184];
    assign _3975 = _3968 & _3974;
    assign _3978 = _3975 & _3977;
    assign _4006 = _3978 ? _3971 : _290;
    assign _4004 = _3998 ? _290 : _3991;
    assign _4007 = _4004 + _4006;
    assign _4021 = _4007 + _4020;
    assign _6718 = _287 ? _4021 : _3991;
    assign _6724 = _278 ? _6723 : _6718;
    assign _193 = _6724;
    always @(posedge _272) begin
        if (_270)
            _3991 <= _290;
        else
            _3991 <= _193;
    end
    assign _3993 = _3991 == _290;
    assign _3994 = ~ _3993;
    assign _3988 = _265[185:185];
    assign _3995 = _3988 & _3994;
    assign _3998 = _3995 & _3997;
    assign _4026 = _3998 ? _3991 : _290;
    assign _4024 = _4018 ? _290 : _4011;
    assign _4027 = _4024 + _4026;
    assign _4041 = _4027 + _4040;
    assign _6725 = _287 ? _4041 : _4011;
    assign _6731 = _278 ? _6730 : _6725;
    assign _194 = _6731;
    always @(posedge _272) begin
        if (_270)
            _4011 <= _290;
        else
            _4011 <= _194;
    end
    assign _4013 = _4011 == _290;
    assign _4014 = ~ _4013;
    assign _4008 = _265[186:186];
    assign _4015 = _4008 & _4014;
    assign _4018 = _4015 & _4017;
    assign _4046 = _4018 ? _4011 : _290;
    assign _4044 = _4038 ? _290 : _4031;
    assign _4047 = _4044 + _4046;
    assign _4061 = _4047 + _4060;
    assign _6732 = _287 ? _4061 : _4031;
    assign _6738 = _278 ? _6737 : _6732;
    assign _195 = _6738;
    always @(posedge _272) begin
        if (_270)
            _4031 <= _290;
        else
            _4031 <= _195;
    end
    assign _4033 = _4031 == _290;
    assign _4034 = ~ _4033;
    assign _4028 = _265[187:187];
    assign _4035 = _4028 & _4034;
    assign _4038 = _4035 & _4037;
    assign _4066 = _4038 ? _4031 : _290;
    assign _4064 = _4058 ? _290 : _4051;
    assign _4067 = _4064 + _4066;
    assign _4081 = _4067 + _4080;
    assign _6739 = _287 ? _4081 : _4051;
    assign _6745 = _278 ? _6744 : _6739;
    assign _196 = _6745;
    always @(posedge _272) begin
        if (_270)
            _4051 <= _290;
        else
            _4051 <= _196;
    end
    assign _4053 = _4051 == _290;
    assign _4054 = ~ _4053;
    assign _4048 = _265[188:188];
    assign _4055 = _4048 & _4054;
    assign _4058 = _4055 & _4057;
    assign _4086 = _4058 ? _4051 : _290;
    assign _4084 = _4078 ? _290 : _4071;
    assign _4087 = _4084 + _4086;
    assign _4101 = _4087 + _4100;
    assign _6746 = _287 ? _4101 : _4071;
    assign _6752 = _278 ? _6751 : _6746;
    assign _197 = _6752;
    always @(posedge _272) begin
        if (_270)
            _4071 <= _290;
        else
            _4071 <= _197;
    end
    assign _4073 = _4071 == _290;
    assign _4074 = ~ _4073;
    assign _4068 = _265[189:189];
    assign _4075 = _4068 & _4074;
    assign _4078 = _4075 & _4077;
    assign _4106 = _4078 ? _4071 : _290;
    assign _4104 = _4098 ? _290 : _4091;
    assign _4107 = _4104 + _4106;
    assign _4121 = _4107 + _4120;
    assign _6753 = _287 ? _4121 : _4091;
    assign _6759 = _278 ? _6758 : _6753;
    assign _198 = _6759;
    always @(posedge _272) begin
        if (_270)
            _4091 <= _290;
        else
            _4091 <= _198;
    end
    assign _4093 = _4091 == _290;
    assign _4094 = ~ _4093;
    assign _4088 = _265[190:190];
    assign _4095 = _4088 & _4094;
    assign _4098 = _4095 & _4097;
    assign _4126 = _4098 ? _4091 : _290;
    assign _4124 = _4118 ? _290 : _4111;
    assign _4127 = _4124 + _4126;
    assign _4141 = _4127 + _4140;
    assign _6760 = _287 ? _4141 : _4111;
    assign _6766 = _278 ? _6765 : _6760;
    assign _199 = _6766;
    always @(posedge _272) begin
        if (_270)
            _4111 <= _290;
        else
            _4111 <= _199;
    end
    assign _4113 = _4111 == _290;
    assign _4114 = ~ _4113;
    assign _4108 = _265[191:191];
    assign _4115 = _4108 & _4114;
    assign _4118 = _4115 & _4117;
    assign _4146 = _4118 ? _4111 : _290;
    assign _4144 = _4138 ? _290 : _4131;
    assign _4147 = _4144 + _4146;
    assign _4161 = _4147 + _4160;
    assign _6767 = _287 ? _4161 : _4131;
    assign _6773 = _278 ? _6772 : _6767;
    assign _200 = _6773;
    always @(posedge _272) begin
        if (_270)
            _4131 <= _290;
        else
            _4131 <= _200;
    end
    assign _4133 = _4131 == _290;
    assign _4134 = ~ _4133;
    assign _4128 = _265[192:192];
    assign _4135 = _4128 & _4134;
    assign _4138 = _4135 & _4137;
    assign _4166 = _4138 ? _4131 : _290;
    assign _4164 = _4158 ? _290 : _4151;
    assign _4167 = _4164 + _4166;
    assign _4181 = _4167 + _4180;
    assign _6774 = _287 ? _4181 : _4151;
    assign _6780 = _278 ? _6779 : _6774;
    assign _201 = _6780;
    always @(posedge _272) begin
        if (_270)
            _4151 <= _290;
        else
            _4151 <= _201;
    end
    assign _4153 = _4151 == _290;
    assign _4154 = ~ _4153;
    assign _4148 = _265[193:193];
    assign _4155 = _4148 & _4154;
    assign _4158 = _4155 & _4157;
    assign _4186 = _4158 ? _4151 : _290;
    assign _4184 = _4178 ? _290 : _4171;
    assign _4187 = _4184 + _4186;
    assign _4201 = _4187 + _4200;
    assign _6781 = _287 ? _4201 : _4171;
    assign _6787 = _278 ? _6786 : _6781;
    assign _202 = _6787;
    always @(posedge _272) begin
        if (_270)
            _4171 <= _290;
        else
            _4171 <= _202;
    end
    assign _4173 = _4171 == _290;
    assign _4174 = ~ _4173;
    assign _4168 = _265[194:194];
    assign _4175 = _4168 & _4174;
    assign _4178 = _4175 & _4177;
    assign _4206 = _4178 ? _4171 : _290;
    assign _4204 = _4198 ? _290 : _4191;
    assign _4207 = _4204 + _4206;
    assign _4221 = _4207 + _4220;
    assign _6788 = _287 ? _4221 : _4191;
    assign _6794 = _278 ? _6793 : _6788;
    assign _203 = _6794;
    always @(posedge _272) begin
        if (_270)
            _4191 <= _290;
        else
            _4191 <= _203;
    end
    assign _4193 = _4191 == _290;
    assign _4194 = ~ _4193;
    assign _4188 = _265[195:195];
    assign _4195 = _4188 & _4194;
    assign _4198 = _4195 & _4197;
    assign _4226 = _4198 ? _4191 : _290;
    assign _4224 = _4218 ? _290 : _4211;
    assign _4227 = _4224 + _4226;
    assign _4241 = _4227 + _4240;
    assign _6795 = _287 ? _4241 : _4211;
    assign _6801 = _278 ? _6800 : _6795;
    assign _204 = _6801;
    always @(posedge _272) begin
        if (_270)
            _4211 <= _290;
        else
            _4211 <= _204;
    end
    assign _4213 = _4211 == _290;
    assign _4214 = ~ _4213;
    assign _4208 = _265[196:196];
    assign _4215 = _4208 & _4214;
    assign _4218 = _4215 & _4217;
    assign _4246 = _4218 ? _4211 : _290;
    assign _4244 = _4238 ? _290 : _4231;
    assign _4247 = _4244 + _4246;
    assign _4261 = _4247 + _4260;
    assign _6802 = _287 ? _4261 : _4231;
    assign _6808 = _278 ? _6807 : _6802;
    assign _205 = _6808;
    always @(posedge _272) begin
        if (_270)
            _4231 <= _290;
        else
            _4231 <= _205;
    end
    assign _4233 = _4231 == _290;
    assign _4234 = ~ _4233;
    assign _4228 = _265[197:197];
    assign _4235 = _4228 & _4234;
    assign _4238 = _4235 & _4237;
    assign _4266 = _4238 ? _4231 : _290;
    assign _4264 = _4258 ? _290 : _4251;
    assign _4267 = _4264 + _4266;
    assign _4281 = _4267 + _4280;
    assign _6809 = _287 ? _4281 : _4251;
    assign _6815 = _278 ? _6814 : _6809;
    assign _206 = _6815;
    always @(posedge _272) begin
        if (_270)
            _4251 <= _290;
        else
            _4251 <= _206;
    end
    assign _4253 = _4251 == _290;
    assign _4254 = ~ _4253;
    assign _4248 = _265[198:198];
    assign _4255 = _4248 & _4254;
    assign _4258 = _4255 & _4257;
    assign _4286 = _4258 ? _4251 : _290;
    assign _4284 = _4278 ? _290 : _4271;
    assign _4287 = _4284 + _4286;
    assign _4301 = _4287 + _4300;
    assign _6816 = _287 ? _4301 : _4271;
    assign _6822 = _278 ? _6821 : _6816;
    assign _207 = _6822;
    always @(posedge _272) begin
        if (_270)
            _4271 <= _290;
        else
            _4271 <= _207;
    end
    assign _4273 = _4271 == _290;
    assign _4274 = ~ _4273;
    assign _4268 = _265[199:199];
    assign _4275 = _4268 & _4274;
    assign _4278 = _4275 & _4277;
    assign _4306 = _4278 ? _4271 : _290;
    assign _4304 = _4298 ? _290 : _4291;
    assign _4307 = _4304 + _4306;
    assign _4321 = _4307 + _4320;
    assign _6823 = _287 ? _4321 : _4291;
    assign _6829 = _278 ? _6828 : _6823;
    assign _208 = _6829;
    always @(posedge _272) begin
        if (_270)
            _4291 <= _290;
        else
            _4291 <= _208;
    end
    assign _4293 = _4291 == _290;
    assign _4294 = ~ _4293;
    assign _4288 = _265[200:200];
    assign _4295 = _4288 & _4294;
    assign _4298 = _4295 & _4297;
    assign _4326 = _4298 ? _4291 : _290;
    assign _4324 = _4318 ? _290 : _4311;
    assign _4327 = _4324 + _4326;
    assign _4341 = _4327 + _4340;
    assign _6830 = _287 ? _4341 : _4311;
    assign _6836 = _278 ? _6835 : _6830;
    assign _209 = _6836;
    always @(posedge _272) begin
        if (_270)
            _4311 <= _290;
        else
            _4311 <= _209;
    end
    assign _4313 = _4311 == _290;
    assign _4314 = ~ _4313;
    assign _4308 = _265[201:201];
    assign _4315 = _4308 & _4314;
    assign _4318 = _4315 & _4317;
    assign _4346 = _4318 ? _4311 : _290;
    assign _4344 = _4338 ? _290 : _4331;
    assign _4347 = _4344 + _4346;
    assign _4361 = _4347 + _4360;
    assign _6837 = _287 ? _4361 : _4331;
    assign _6843 = _278 ? _6842 : _6837;
    assign _210 = _6843;
    always @(posedge _272) begin
        if (_270)
            _4331 <= _290;
        else
            _4331 <= _210;
    end
    assign _4333 = _4331 == _290;
    assign _4334 = ~ _4333;
    assign _4328 = _265[202:202];
    assign _4335 = _4328 & _4334;
    assign _4338 = _4335 & _4337;
    assign _4366 = _4338 ? _4331 : _290;
    assign _4364 = _4358 ? _290 : _4351;
    assign _4367 = _4364 + _4366;
    assign _4381 = _4367 + _4380;
    assign _6844 = _287 ? _4381 : _4351;
    assign _6850 = _278 ? _6849 : _6844;
    assign _211 = _6850;
    always @(posedge _272) begin
        if (_270)
            _4351 <= _290;
        else
            _4351 <= _211;
    end
    assign _4353 = _4351 == _290;
    assign _4354 = ~ _4353;
    assign _4348 = _265[203:203];
    assign _4355 = _4348 & _4354;
    assign _4358 = _4355 & _4357;
    assign _4386 = _4358 ? _4351 : _290;
    assign _4384 = _4378 ? _290 : _4371;
    assign _4387 = _4384 + _4386;
    assign _4401 = _4387 + _4400;
    assign _6851 = _287 ? _4401 : _4371;
    assign _6857 = _278 ? _6856 : _6851;
    assign _212 = _6857;
    always @(posedge _272) begin
        if (_270)
            _4371 <= _290;
        else
            _4371 <= _212;
    end
    assign _4373 = _4371 == _290;
    assign _4374 = ~ _4373;
    assign _4368 = _265[204:204];
    assign _4375 = _4368 & _4374;
    assign _4378 = _4375 & _4377;
    assign _4406 = _4378 ? _4371 : _290;
    assign _4404 = _4398 ? _290 : _4391;
    assign _4407 = _4404 + _4406;
    assign _4421 = _4407 + _4420;
    assign _6858 = _287 ? _4421 : _4391;
    assign _6864 = _278 ? _6863 : _6858;
    assign _213 = _6864;
    always @(posedge _272) begin
        if (_270)
            _4391 <= _290;
        else
            _4391 <= _213;
    end
    assign _4393 = _4391 == _290;
    assign _4394 = ~ _4393;
    assign _4388 = _265[205:205];
    assign _4395 = _4388 & _4394;
    assign _4398 = _4395 & _4397;
    assign _4426 = _4398 ? _4391 : _290;
    assign _4424 = _4418 ? _290 : _4411;
    assign _4427 = _4424 + _4426;
    assign _4441 = _4427 + _4440;
    assign _6865 = _287 ? _4441 : _4411;
    assign _6871 = _278 ? _6870 : _6865;
    assign _214 = _6871;
    always @(posedge _272) begin
        if (_270)
            _4411 <= _290;
        else
            _4411 <= _214;
    end
    assign _4413 = _4411 == _290;
    assign _4414 = ~ _4413;
    assign _4408 = _265[206:206];
    assign _4415 = _4408 & _4414;
    assign _4418 = _4415 & _4417;
    assign _4446 = _4418 ? _4411 : _290;
    assign _4444 = _4438 ? _290 : _4431;
    assign _4447 = _4444 + _4446;
    assign _4461 = _4447 + _4460;
    assign _6872 = _287 ? _4461 : _4431;
    assign _6878 = _278 ? _6877 : _6872;
    assign _215 = _6878;
    always @(posedge _272) begin
        if (_270)
            _4431 <= _290;
        else
            _4431 <= _215;
    end
    assign _4433 = _4431 == _290;
    assign _4434 = ~ _4433;
    assign _4428 = _265[207:207];
    assign _4435 = _4428 & _4434;
    assign _4438 = _4435 & _4437;
    assign _4466 = _4438 ? _4431 : _290;
    assign _4464 = _4458 ? _290 : _4451;
    assign _4467 = _4464 + _4466;
    assign _4481 = _4467 + _4480;
    assign _6879 = _287 ? _4481 : _4451;
    assign _6885 = _278 ? _6884 : _6879;
    assign _216 = _6885;
    always @(posedge _272) begin
        if (_270)
            _4451 <= _290;
        else
            _4451 <= _216;
    end
    assign _4453 = _4451 == _290;
    assign _4454 = ~ _4453;
    assign _4448 = _265[208:208];
    assign _4455 = _4448 & _4454;
    assign _4458 = _4455 & _4457;
    assign _4486 = _4458 ? _4451 : _290;
    assign _4484 = _4478 ? _290 : _4471;
    assign _4487 = _4484 + _4486;
    assign _4501 = _4487 + _4500;
    assign _6886 = _287 ? _4501 : _4471;
    assign _6892 = _278 ? _6891 : _6886;
    assign _217 = _6892;
    always @(posedge _272) begin
        if (_270)
            _4471 <= _290;
        else
            _4471 <= _217;
    end
    assign _4473 = _4471 == _290;
    assign _4474 = ~ _4473;
    assign _4468 = _265[209:209];
    assign _4475 = _4468 & _4474;
    assign _4478 = _4475 & _4477;
    assign _4506 = _4478 ? _4471 : _290;
    assign _4504 = _4498 ? _290 : _4491;
    assign _4507 = _4504 + _4506;
    assign _4521 = _4507 + _4520;
    assign _6893 = _287 ? _4521 : _4491;
    assign _6899 = _278 ? _6898 : _6893;
    assign _218 = _6899;
    always @(posedge _272) begin
        if (_270)
            _4491 <= _290;
        else
            _4491 <= _218;
    end
    assign _4493 = _4491 == _290;
    assign _4494 = ~ _4493;
    assign _4488 = _265[210:210];
    assign _4495 = _4488 & _4494;
    assign _4498 = _4495 & _4497;
    assign _4526 = _4498 ? _4491 : _290;
    assign _4524 = _4518 ? _290 : _4511;
    assign _4527 = _4524 + _4526;
    assign _4541 = _4527 + _4540;
    assign _6900 = _287 ? _4541 : _4511;
    assign _6906 = _278 ? _6905 : _6900;
    assign _219 = _6906;
    always @(posedge _272) begin
        if (_270)
            _4511 <= _290;
        else
            _4511 <= _219;
    end
    assign _4513 = _4511 == _290;
    assign _4514 = ~ _4513;
    assign _4508 = _265[211:211];
    assign _4515 = _4508 & _4514;
    assign _4518 = _4515 & _4517;
    assign _4546 = _4518 ? _4511 : _290;
    assign _4544 = _4538 ? _290 : _4531;
    assign _4547 = _4544 + _4546;
    assign _4561 = _4547 + _4560;
    assign _6907 = _287 ? _4561 : _4531;
    assign _6913 = _278 ? _6912 : _6907;
    assign _220 = _6913;
    always @(posedge _272) begin
        if (_270)
            _4531 <= _290;
        else
            _4531 <= _220;
    end
    assign _4533 = _4531 == _290;
    assign _4534 = ~ _4533;
    assign _4528 = _265[212:212];
    assign _4535 = _4528 & _4534;
    assign _4538 = _4535 & _4537;
    assign _4566 = _4538 ? _4531 : _290;
    assign _4564 = _4558 ? _290 : _4551;
    assign _4567 = _4564 + _4566;
    assign _4581 = _4567 + _4580;
    assign _6914 = _287 ? _4581 : _4551;
    assign _6920 = _278 ? _6919 : _6914;
    assign _221 = _6920;
    always @(posedge _272) begin
        if (_270)
            _4551 <= _290;
        else
            _4551 <= _221;
    end
    assign _4553 = _4551 == _290;
    assign _4554 = ~ _4553;
    assign _4548 = _265[213:213];
    assign _4555 = _4548 & _4554;
    assign _4558 = _4555 & _4557;
    assign _4586 = _4558 ? _4551 : _290;
    assign _4584 = _4578 ? _290 : _4571;
    assign _4587 = _4584 + _4586;
    assign _4601 = _4587 + _4600;
    assign _6921 = _287 ? _4601 : _4571;
    assign _6927 = _278 ? _6926 : _6921;
    assign _222 = _6927;
    always @(posedge _272) begin
        if (_270)
            _4571 <= _290;
        else
            _4571 <= _222;
    end
    assign _4573 = _4571 == _290;
    assign _4574 = ~ _4573;
    assign _4568 = _265[214:214];
    assign _4575 = _4568 & _4574;
    assign _4578 = _4575 & _4577;
    assign _4606 = _4578 ? _4571 : _290;
    assign _4604 = _4598 ? _290 : _4591;
    assign _4607 = _4604 + _4606;
    assign _4621 = _4607 + _4620;
    assign _6928 = _287 ? _4621 : _4591;
    assign _6934 = _278 ? _6933 : _6928;
    assign _223 = _6934;
    always @(posedge _272) begin
        if (_270)
            _4591 <= _290;
        else
            _4591 <= _223;
    end
    assign _4593 = _4591 == _290;
    assign _4594 = ~ _4593;
    assign _4588 = _265[215:215];
    assign _4595 = _4588 & _4594;
    assign _4598 = _4595 & _4597;
    assign _4626 = _4598 ? _4591 : _290;
    assign _4624 = _4618 ? _290 : _4611;
    assign _4627 = _4624 + _4626;
    assign _4641 = _4627 + _4640;
    assign _6935 = _287 ? _4641 : _4611;
    assign _6941 = _278 ? _6940 : _6935;
    assign _224 = _6941;
    always @(posedge _272) begin
        if (_270)
            _4611 <= _290;
        else
            _4611 <= _224;
    end
    assign _4613 = _4611 == _290;
    assign _4614 = ~ _4613;
    assign _4608 = _265[216:216];
    assign _4615 = _4608 & _4614;
    assign _4618 = _4615 & _4617;
    assign _4646 = _4618 ? _4611 : _290;
    assign _4644 = _4638 ? _290 : _4631;
    assign _4647 = _4644 + _4646;
    assign _4661 = _4647 + _4660;
    assign _6942 = _287 ? _4661 : _4631;
    assign _6948 = _278 ? _6947 : _6942;
    assign _225 = _6948;
    always @(posedge _272) begin
        if (_270)
            _4631 <= _290;
        else
            _4631 <= _225;
    end
    assign _4633 = _4631 == _290;
    assign _4634 = ~ _4633;
    assign _4628 = _265[217:217];
    assign _4635 = _4628 & _4634;
    assign _4638 = _4635 & _4637;
    assign _4666 = _4638 ? _4631 : _290;
    assign _4664 = _4658 ? _290 : _4651;
    assign _4667 = _4664 + _4666;
    assign _4681 = _4667 + _4680;
    assign _6949 = _287 ? _4681 : _4651;
    assign _6955 = _278 ? _6954 : _6949;
    assign _226 = _6955;
    always @(posedge _272) begin
        if (_270)
            _4651 <= _290;
        else
            _4651 <= _226;
    end
    assign _4653 = _4651 == _290;
    assign _4654 = ~ _4653;
    assign _4648 = _265[218:218];
    assign _4655 = _4648 & _4654;
    assign _4658 = _4655 & _4657;
    assign _4686 = _4658 ? _4651 : _290;
    assign _4684 = _4678 ? _290 : _4671;
    assign _4687 = _4684 + _4686;
    assign _4701 = _4687 + _4700;
    assign _6956 = _287 ? _4701 : _4671;
    assign _6962 = _278 ? _6961 : _6956;
    assign _227 = _6962;
    always @(posedge _272) begin
        if (_270)
            _4671 <= _290;
        else
            _4671 <= _227;
    end
    assign _4673 = _4671 == _290;
    assign _4674 = ~ _4673;
    assign _4668 = _265[219:219];
    assign _4675 = _4668 & _4674;
    assign _4678 = _4675 & _4677;
    assign _4706 = _4678 ? _4671 : _290;
    assign _4704 = _4698 ? _290 : _4691;
    assign _4707 = _4704 + _4706;
    assign _4721 = _4707 + _4720;
    assign _6963 = _287 ? _4721 : _4691;
    assign _6969 = _278 ? _6968 : _6963;
    assign _228 = _6969;
    always @(posedge _272) begin
        if (_270)
            _4691 <= _290;
        else
            _4691 <= _228;
    end
    assign _4693 = _4691 == _290;
    assign _4694 = ~ _4693;
    assign _4688 = _265[220:220];
    assign _4695 = _4688 & _4694;
    assign _4698 = _4695 & _4697;
    assign _4726 = _4698 ? _4691 : _290;
    assign _4724 = _4718 ? _290 : _4711;
    assign _4727 = _4724 + _4726;
    assign _4741 = _4727 + _4740;
    assign _6970 = _287 ? _4741 : _4711;
    assign _6976 = _278 ? _6975 : _6970;
    assign _229 = _6976;
    always @(posedge _272) begin
        if (_270)
            _4711 <= _290;
        else
            _4711 <= _229;
    end
    assign _4713 = _4711 == _290;
    assign _4714 = ~ _4713;
    assign _4708 = _265[221:221];
    assign _4715 = _4708 & _4714;
    assign _4718 = _4715 & _4717;
    assign _4746 = _4718 ? _4711 : _290;
    assign _4744 = _4738 ? _290 : _4731;
    assign _4747 = _4744 + _4746;
    assign _4761 = _4747 + _4760;
    assign _6977 = _287 ? _4761 : _4731;
    assign _6983 = _278 ? _6982 : _6977;
    assign _230 = _6983;
    always @(posedge _272) begin
        if (_270)
            _4731 <= _290;
        else
            _4731 <= _230;
    end
    assign _4733 = _4731 == _290;
    assign _4734 = ~ _4733;
    assign _4728 = _265[222:222];
    assign _4735 = _4728 & _4734;
    assign _4738 = _4735 & _4737;
    assign _4766 = _4738 ? _4731 : _290;
    assign _4764 = _4758 ? _290 : _4751;
    assign _4767 = _4764 + _4766;
    assign _4781 = _4767 + _4780;
    assign _6984 = _287 ? _4781 : _4751;
    assign _6990 = _278 ? _6989 : _6984;
    assign _231 = _6990;
    always @(posedge _272) begin
        if (_270)
            _4751 <= _290;
        else
            _4751 <= _231;
    end
    assign _4753 = _4751 == _290;
    assign _4754 = ~ _4753;
    assign _4748 = _265[223:223];
    assign _4755 = _4748 & _4754;
    assign _4758 = _4755 & _4757;
    assign _4786 = _4758 ? _4751 : _290;
    assign _4784 = _4778 ? _290 : _4771;
    assign _4787 = _4784 + _4786;
    assign _4801 = _4787 + _4800;
    assign _6991 = _287 ? _4801 : _4771;
    assign _6997 = _278 ? _6996 : _6991;
    assign _232 = _6997;
    always @(posedge _272) begin
        if (_270)
            _4771 <= _290;
        else
            _4771 <= _232;
    end
    assign _4773 = _4771 == _290;
    assign _4774 = ~ _4773;
    assign _4768 = _265[224:224];
    assign _4775 = _4768 & _4774;
    assign _4778 = _4775 & _4777;
    assign _4806 = _4778 ? _4771 : _290;
    assign _4804 = _4798 ? _290 : _4791;
    assign _4807 = _4804 + _4806;
    assign _4821 = _4807 + _4820;
    assign _6998 = _287 ? _4821 : _4791;
    assign _7004 = _278 ? _7003 : _6998;
    assign _233 = _7004;
    always @(posedge _272) begin
        if (_270)
            _4791 <= _290;
        else
            _4791 <= _233;
    end
    assign _4793 = _4791 == _290;
    assign _4794 = ~ _4793;
    assign _4788 = _265[225:225];
    assign _4795 = _4788 & _4794;
    assign _4798 = _4795 & _4797;
    assign _4826 = _4798 ? _4791 : _290;
    assign _4824 = _4818 ? _290 : _4811;
    assign _4827 = _4824 + _4826;
    assign _4841 = _4827 + _4840;
    assign _7005 = _287 ? _4841 : _4811;
    assign _7011 = _278 ? _7010 : _7005;
    assign _234 = _7011;
    always @(posedge _272) begin
        if (_270)
            _4811 <= _290;
        else
            _4811 <= _234;
    end
    assign _4813 = _4811 == _290;
    assign _4814 = ~ _4813;
    assign _4808 = _265[226:226];
    assign _4815 = _4808 & _4814;
    assign _4818 = _4815 & _4817;
    assign _4846 = _4818 ? _4811 : _290;
    assign _4844 = _4838 ? _290 : _4831;
    assign _4847 = _4844 + _4846;
    assign _4861 = _4847 + _4860;
    assign _7012 = _287 ? _4861 : _4831;
    assign _7018 = _278 ? _7017 : _7012;
    assign _235 = _7018;
    always @(posedge _272) begin
        if (_270)
            _4831 <= _290;
        else
            _4831 <= _235;
    end
    assign _4833 = _4831 == _290;
    assign _4834 = ~ _4833;
    assign _4828 = _265[227:227];
    assign _4835 = _4828 & _4834;
    assign _4838 = _4835 & _4837;
    assign _4866 = _4838 ? _4831 : _290;
    assign _4864 = _4858 ? _290 : _4851;
    assign _4867 = _4864 + _4866;
    assign _4881 = _4867 + _4880;
    assign _7019 = _287 ? _4881 : _4851;
    assign _7025 = _278 ? _7024 : _7019;
    assign _236 = _7025;
    always @(posedge _272) begin
        if (_270)
            _4851 <= _290;
        else
            _4851 <= _236;
    end
    assign _4853 = _4851 == _290;
    assign _4854 = ~ _4853;
    assign _4848 = _265[228:228];
    assign _4855 = _4848 & _4854;
    assign _4858 = _4855 & _4857;
    assign _4886 = _4858 ? _4851 : _290;
    assign _4884 = _4878 ? _290 : _4871;
    assign _4887 = _4884 + _4886;
    assign _4901 = _4887 + _4900;
    assign _7026 = _287 ? _4901 : _4871;
    assign _7032 = _278 ? _7031 : _7026;
    assign _237 = _7032;
    always @(posedge _272) begin
        if (_270)
            _4871 <= _290;
        else
            _4871 <= _237;
    end
    assign _4873 = _4871 == _290;
    assign _4874 = ~ _4873;
    assign _4868 = _265[229:229];
    assign _4875 = _4868 & _4874;
    assign _4878 = _4875 & _4877;
    assign _4906 = _4878 ? _4871 : _290;
    assign _4904 = _4898 ? _290 : _4891;
    assign _4907 = _4904 + _4906;
    assign _4921 = _4907 + _4920;
    assign _7033 = _287 ? _4921 : _4891;
    assign _7039 = _278 ? _7038 : _7033;
    assign _238 = _7039;
    always @(posedge _272) begin
        if (_270)
            _4891 <= _290;
        else
            _4891 <= _238;
    end
    assign _4893 = _4891 == _290;
    assign _4894 = ~ _4893;
    assign _4888 = _265[230:230];
    assign _4895 = _4888 & _4894;
    assign _4898 = _4895 & _4897;
    assign _4926 = _4898 ? _4891 : _290;
    assign _4924 = _4918 ? _290 : _4911;
    assign _4927 = _4924 + _4926;
    assign _4941 = _4927 + _4940;
    assign _7040 = _287 ? _4941 : _4911;
    assign _7046 = _278 ? _7045 : _7040;
    assign _239 = _7046;
    always @(posedge _272) begin
        if (_270)
            _4911 <= _290;
        else
            _4911 <= _239;
    end
    assign _4913 = _4911 == _290;
    assign _4914 = ~ _4913;
    assign _4908 = _265[231:231];
    assign _4915 = _4908 & _4914;
    assign _4918 = _4915 & _4917;
    assign _4946 = _4918 ? _4911 : _290;
    assign _4944 = _4938 ? _290 : _4931;
    assign _4947 = _4944 + _4946;
    assign _4961 = _4947 + _4960;
    assign _7047 = _287 ? _4961 : _4931;
    assign _7053 = _278 ? _7052 : _7047;
    assign _240 = _7053;
    always @(posedge _272) begin
        if (_270)
            _4931 <= _290;
        else
            _4931 <= _240;
    end
    assign _4933 = _4931 == _290;
    assign _4934 = ~ _4933;
    assign _4928 = _265[232:232];
    assign _4935 = _4928 & _4934;
    assign _4938 = _4935 & _4937;
    assign _4966 = _4938 ? _4931 : _290;
    assign _4964 = _4958 ? _290 : _4951;
    assign _4967 = _4964 + _4966;
    assign _4981 = _4967 + _4980;
    assign _7054 = _287 ? _4981 : _4951;
    assign _7060 = _278 ? _7059 : _7054;
    assign _241 = _7060;
    always @(posedge _272) begin
        if (_270)
            _4951 <= _290;
        else
            _4951 <= _241;
    end
    assign _4953 = _4951 == _290;
    assign _4954 = ~ _4953;
    assign _4948 = _265[233:233];
    assign _4955 = _4948 & _4954;
    assign _4958 = _4955 & _4957;
    assign _4986 = _4958 ? _4951 : _290;
    assign _4984 = _4978 ? _290 : _4971;
    assign _4987 = _4984 + _4986;
    assign _5001 = _4987 + _5000;
    assign _7061 = _287 ? _5001 : _4971;
    assign _7067 = _278 ? _7066 : _7061;
    assign _242 = _7067;
    always @(posedge _272) begin
        if (_270)
            _4971 <= _290;
        else
            _4971 <= _242;
    end
    assign _4973 = _4971 == _290;
    assign _4974 = ~ _4973;
    assign _4968 = _265[234:234];
    assign _4975 = _4968 & _4974;
    assign _4978 = _4975 & _4977;
    assign _5006 = _4978 ? _4971 : _290;
    assign _5004 = _4998 ? _290 : _4991;
    assign _5007 = _5004 + _5006;
    assign _5021 = _5007 + _5020;
    assign _7068 = _287 ? _5021 : _4991;
    assign _7074 = _278 ? _7073 : _7068;
    assign _243 = _7074;
    always @(posedge _272) begin
        if (_270)
            _4991 <= _290;
        else
            _4991 <= _243;
    end
    assign _4993 = _4991 == _290;
    assign _4994 = ~ _4993;
    assign _4988 = _265[235:235];
    assign _4995 = _4988 & _4994;
    assign _4998 = _4995 & _4997;
    assign _5026 = _4998 ? _4991 : _290;
    assign _5024 = _5018 ? _290 : _5011;
    assign _5027 = _5024 + _5026;
    assign _5041 = _5027 + _5040;
    assign _7075 = _287 ? _5041 : _5011;
    assign _7081 = _278 ? _7080 : _7075;
    assign _244 = _7081;
    always @(posedge _272) begin
        if (_270)
            _5011 <= _290;
        else
            _5011 <= _244;
    end
    assign _5013 = _5011 == _290;
    assign _5014 = ~ _5013;
    assign _5008 = _265[236:236];
    assign _5015 = _5008 & _5014;
    assign _5018 = _5015 & _5017;
    assign _5046 = _5018 ? _5011 : _290;
    assign _5044 = _5038 ? _290 : _5031;
    assign _5047 = _5044 + _5046;
    assign _5061 = _5047 + _5060;
    assign _7082 = _287 ? _5061 : _5031;
    assign _7088 = _278 ? _7087 : _7082;
    assign _245 = _7088;
    always @(posedge _272) begin
        if (_270)
            _5031 <= _290;
        else
            _5031 <= _245;
    end
    assign _5033 = _5031 == _290;
    assign _5034 = ~ _5033;
    assign _5028 = _265[237:237];
    assign _5035 = _5028 & _5034;
    assign _5038 = _5035 & _5037;
    assign _5066 = _5038 ? _5031 : _290;
    assign _5064 = _5058 ? _290 : _5051;
    assign _5067 = _5064 + _5066;
    assign _5081 = _5067 + _5080;
    assign _7089 = _287 ? _5081 : _5051;
    assign _7095 = _278 ? _7094 : _7089;
    assign _246 = _7095;
    always @(posedge _272) begin
        if (_270)
            _5051 <= _290;
        else
            _5051 <= _246;
    end
    assign _5053 = _5051 == _290;
    assign _5054 = ~ _5053;
    assign _5048 = _265[238:238];
    assign _5055 = _5048 & _5054;
    assign _5058 = _5055 & _5057;
    assign _5086 = _5058 ? _5051 : _290;
    assign _5084 = _5078 ? _290 : _5071;
    assign _5087 = _5084 + _5086;
    assign _5101 = _5087 + _5100;
    assign _7096 = _287 ? _5101 : _5071;
    assign _7102 = _278 ? _7101 : _7096;
    assign _247 = _7102;
    always @(posedge _272) begin
        if (_270)
            _5071 <= _290;
        else
            _5071 <= _247;
    end
    assign _5073 = _5071 == _290;
    assign _5074 = ~ _5073;
    assign _5068 = _265[239:239];
    assign _5075 = _5068 & _5074;
    assign _5078 = _5075 & _5077;
    assign _5106 = _5078 ? _5071 : _290;
    assign _5104 = _5098 ? _290 : _5091;
    assign _5107 = _5104 + _5106;
    assign _5121 = _5107 + _5120;
    assign _7103 = _287 ? _5121 : _5091;
    assign _7109 = _278 ? _7108 : _7103;
    assign _248 = _7109;
    always @(posedge _272) begin
        if (_270)
            _5091 <= _290;
        else
            _5091 <= _248;
    end
    assign _5093 = _5091 == _290;
    assign _5094 = ~ _5093;
    assign _5088 = _265[240:240];
    assign _5095 = _5088 & _5094;
    assign _5098 = _5095 & _5097;
    assign _5126 = _5098 ? _5091 : _290;
    assign _5124 = _5118 ? _290 : _5111;
    assign _5127 = _5124 + _5126;
    assign _5141 = _5127 + _5140;
    assign _7110 = _287 ? _5141 : _5111;
    assign _7116 = _278 ? _7115 : _7110;
    assign _249 = _7116;
    always @(posedge _272) begin
        if (_270)
            _5111 <= _290;
        else
            _5111 <= _249;
    end
    assign _5113 = _5111 == _290;
    assign _5114 = ~ _5113;
    assign _5108 = _265[241:241];
    assign _5115 = _5108 & _5114;
    assign _5118 = _5115 & _5117;
    assign _5146 = _5118 ? _5111 : _290;
    assign _5144 = _5138 ? _290 : _5131;
    assign _5147 = _5144 + _5146;
    assign _5161 = _5147 + _5160;
    assign _7117 = _287 ? _5161 : _5131;
    assign _7123 = _278 ? _7122 : _7117;
    assign _250 = _7123;
    always @(posedge _272) begin
        if (_270)
            _5131 <= _290;
        else
            _5131 <= _250;
    end
    assign _5133 = _5131 == _290;
    assign _5134 = ~ _5133;
    assign _5128 = _265[242:242];
    assign _5135 = _5128 & _5134;
    assign _5138 = _5135 & _5137;
    assign _5166 = _5138 ? _5131 : _290;
    assign _5164 = _5158 ? _290 : _5151;
    assign _5167 = _5164 + _5166;
    assign _5181 = _5167 + _5180;
    assign _7124 = _287 ? _5181 : _5151;
    assign _7130 = _278 ? _7129 : _7124;
    assign _251 = _7130;
    always @(posedge _272) begin
        if (_270)
            _5151 <= _290;
        else
            _5151 <= _251;
    end
    assign _5153 = _5151 == _290;
    assign _5154 = ~ _5153;
    assign _5148 = _265[243:243];
    assign _5155 = _5148 & _5154;
    assign _5158 = _5155 & _5157;
    assign _5186 = _5158 ? _5151 : _290;
    assign _5184 = _5178 ? _290 : _5171;
    assign _5187 = _5184 + _5186;
    assign _5201 = _5187 + _5200;
    assign _7131 = _287 ? _5201 : _5171;
    assign _7137 = _278 ? _7136 : _7131;
    assign _252 = _7137;
    always @(posedge _272) begin
        if (_270)
            _5171 <= _290;
        else
            _5171 <= _252;
    end
    assign _5173 = _5171 == _290;
    assign _5174 = ~ _5173;
    assign _5168 = _265[244:244];
    assign _5175 = _5168 & _5174;
    assign _5178 = _5175 & _5177;
    assign _5206 = _5178 ? _5171 : _290;
    assign _5204 = _5198 ? _290 : _5191;
    assign _5207 = _5204 + _5206;
    assign _5221 = _5207 + _5220;
    assign _7138 = _287 ? _5221 : _5191;
    assign _7144 = _278 ? _7143 : _7138;
    assign _253 = _7144;
    always @(posedge _272) begin
        if (_270)
            _5191 <= _290;
        else
            _5191 <= _253;
    end
    assign _5193 = _5191 == _290;
    assign _5194 = ~ _5193;
    assign _5188 = _265[245:245];
    assign _5195 = _5188 & _5194;
    assign _5198 = _5195 & _5197;
    assign _5226 = _5198 ? _5191 : _290;
    assign _5224 = _5218 ? _290 : _5211;
    assign _5227 = _5224 + _5226;
    assign _5241 = _5227 + _5240;
    assign _7145 = _287 ? _5241 : _5211;
    assign _7151 = _278 ? _7150 : _7145;
    assign _254 = _7151;
    always @(posedge _272) begin
        if (_270)
            _5211 <= _290;
        else
            _5211 <= _254;
    end
    assign _5213 = _5211 == _290;
    assign _5214 = ~ _5213;
    assign _5208 = _265[246:246];
    assign _5215 = _5208 & _5214;
    assign _5218 = _5215 & _5217;
    assign _5246 = _5218 ? _5211 : _290;
    assign _5244 = _5238 ? _290 : _5231;
    assign _5247 = _5244 + _5246;
    assign _5261 = _5247 + _5260;
    assign _7152 = _287 ? _5261 : _5231;
    assign _7158 = _278 ? _7157 : _7152;
    assign _255 = _7158;
    always @(posedge _272) begin
        if (_270)
            _5231 <= _290;
        else
            _5231 <= _255;
    end
    assign _5233 = _5231 == _290;
    assign _5234 = ~ _5233;
    assign _5228 = _265[247:247];
    assign _5235 = _5228 & _5234;
    assign _5238 = _5235 & _5237;
    assign _5266 = _5238 ? _5231 : _290;
    assign _5264 = _5258 ? _290 : _5251;
    assign _5267 = _5264 + _5266;
    assign _5281 = _5267 + _5280;
    assign _7159 = _287 ? _5281 : _5251;
    assign _7165 = _278 ? _7164 : _7159;
    assign _256 = _7165;
    always @(posedge _272) begin
        if (_270)
            _5251 <= _290;
        else
            _5251 <= _256;
    end
    assign _5253 = _5251 == _290;
    assign _5254 = ~ _5253;
    assign _5248 = _265[248:248];
    assign _5255 = _5248 & _5254;
    assign _5258 = _5255 & _5257;
    assign _5286 = _5258 ? _5251 : _290;
    assign _5284 = _5278 ? _290 : _5271;
    assign _5287 = _5284 + _5286;
    assign _5301 = _5287 + _5300;
    assign _7166 = _287 ? _5301 : _5271;
    assign _7172 = _278 ? _7171 : _7166;
    assign _257 = _7172;
    always @(posedge _272) begin
        if (_270)
            _5271 <= _290;
        else
            _5271 <= _257;
    end
    assign _5273 = _5271 == _290;
    assign _5274 = ~ _5273;
    assign _5268 = _265[249:249];
    assign _5275 = _5268 & _5274;
    assign _5278 = _5275 & _5277;
    assign _5306 = _5278 ? _5271 : _290;
    assign _5304 = _5298 ? _290 : _5291;
    assign _5307 = _5304 + _5306;
    assign _5321 = _5307 + _5320;
    assign _7173 = _287 ? _5321 : _5291;
    assign _7179 = _278 ? _7178 : _7173;
    assign _258 = _7179;
    always @(posedge _272) begin
        if (_270)
            _5291 <= _290;
        else
            _5291 <= _258;
    end
    assign _5293 = _5291 == _290;
    assign _5294 = ~ _5293;
    assign _5288 = _265[250:250];
    assign _5295 = _5288 & _5294;
    assign _5298 = _5295 & _5297;
    assign _5326 = _5298 ? _5291 : _290;
    assign _5324 = _5318 ? _290 : _5311;
    assign _5327 = _5324 + _5326;
    assign _5341 = _5327 + _5340;
    assign _7180 = _287 ? _5341 : _5311;
    assign _7186 = _278 ? _7185 : _7180;
    assign _259 = _7186;
    always @(posedge _272) begin
        if (_270)
            _5311 <= _290;
        else
            _5311 <= _259;
    end
    assign _5313 = _5311 == _290;
    assign _5314 = ~ _5313;
    assign _5308 = _265[251:251];
    assign _5315 = _5308 & _5314;
    assign _5318 = _5315 & _5317;
    assign _5346 = _5318 ? _5311 : _290;
    assign _5344 = _5338 ? _290 : _5331;
    assign _5347 = _5344 + _5346;
    assign _5361 = _5347 + _5360;
    assign _7187 = _287 ? _5361 : _5331;
    assign _7193 = _278 ? _7192 : _7187;
    assign _260 = _7193;
    always @(posedge _272) begin
        if (_270)
            _5331 <= _290;
        else
            _5331 <= _260;
    end
    assign _5333 = _5331 == _290;
    assign _5334 = ~ _5333;
    assign _5328 = _265[252:252];
    assign _5335 = _5328 & _5334;
    assign _5338 = _5335 & _5337;
    assign _5366 = _5338 ? _5331 : _290;
    assign _5364 = _5358 ? _290 : _5351;
    assign _5367 = _5364 + _5366;
    assign _5381 = _5367 + _5380;
    assign _7194 = _287 ? _5381 : _5351;
    assign _7200 = _278 ? _7199 : _7194;
    assign _261 = _7200;
    always @(posedge _272) begin
        if (_270)
            _5351 <= _290;
        else
            _5351 <= _261;
    end
    assign _5353 = _5351 == _290;
    assign _5354 = ~ _5353;
    assign _5348 = _265[253:253];
    assign _5355 = _5348 & _5354;
    assign _5358 = _5355 & _5357;
    assign _5386 = _5358 ? _5351 : _290;
    assign _5384 = _5378 ? _290 : _5371;
    assign _5387 = _5384 + _5386;
    assign _5401 = _5387 + _5400;
    assign _7201 = _287 ? _5401 : _5371;
    assign _7207 = _278 ? _7206 : _7201;
    assign _262 = _7207;
    always @(posedge _272) begin
        if (_270)
            _5371 <= _290;
        else
            _5371 <= _262;
    end
    assign _5373 = _5371 == _290;
    assign _5374 = ~ _5373;
    assign _5368 = _265[254:254];
    assign _5375 = _5368 & _5374;
    assign _5378 = _5375 & _5377;
    assign _5406 = _5378 ? _5371 : _290;
    assign _5404 = _5398 ? _290 : _5391;
    assign _5407 = _5404 + _5406;
    assign _7208 = _287 ? _5407 : _5391;
    assign _7214 = _278 ? _7213 : _7208;
    assign _263 = _7214;
    always @(posedge _272) begin
        if (_270)
            _5391 <= _290;
        else
            _5391 <= _263;
    end
    assign _5393 = _5391 == _290;
    assign _5394 = ~ _5393;
    assign _265 = row_bits;
    assign _5388 = _265[255:255];
    assign _5395 = _5388 & _5394;
    assign _5398 = _5395 & _5397;
    assign _7220 = { _5398,
                     _5378,
                     _5358,
                     _5338,
                     _5318,
                     _5298,
                     _5278,
                     _5258,
                     _5238,
                     _5218,
                     _5198,
                     _5178,
                     _5158,
                     _5138,
                     _5118,
                     _5098,
                     _5078,
                     _5058,
                     _5038,
                     _5018,
                     _4998,
                     _4978,
                     _4958,
                     _4938,
                     _4918,
                     _4898,
                     _4878,
                     _4858,
                     _4838,
                     _4818,
                     _4798,
                     _4778,
                     _4758,
                     _4738,
                     _4718,
                     _4698,
                     _4678,
                     _4658,
                     _4638,
                     _4618,
                     _4598,
                     _4578,
                     _4558,
                     _4538,
                     _4518,
                     _4498,
                     _4478,
                     _4458,
                     _4438,
                     _4418,
                     _4398,
                     _4378,
                     _4358,
                     _4338,
                     _4318,
                     _4298,
                     _4278,
                     _4258,
                     _4238,
                     _4218,
                     _4198,
                     _4178,
                     _4158,
                     _4138,
                     _4118,
                     _4098,
                     _4078,
                     _4058,
                     _4038,
                     _4018,
                     _3998,
                     _3978,
                     _3958,
                     _3938,
                     _3918,
                     _3898,
                     _3878,
                     _3858,
                     _3838,
                     _3818,
                     _3798,
                     _3778,
                     _3758,
                     _3738,
                     _3718,
                     _3698,
                     _3678,
                     _3658,
                     _3638,
                     _3618,
                     _3598,
                     _3578,
                     _3558,
                     _3538,
                     _3518,
                     _3498,
                     _3478,
                     _3458,
                     _3438,
                     _3418,
                     _3398,
                     _3378,
                     _3358,
                     _3338,
                     _3318,
                     _3298,
                     _3278,
                     _3258,
                     _3238,
                     _3218,
                     _3198,
                     _3178,
                     _3158,
                     _3138,
                     _3118,
                     _3098,
                     _3078,
                     _3058,
                     _3038,
                     _3018,
                     _2998,
                     _2978,
                     _2958,
                     _2938,
                     _2918,
                     _2898,
                     _2878,
                     _2858,
                     _2838,
                     _2818,
                     _2798,
                     _2778,
                     _2758,
                     _2738,
                     _2718,
                     _2698,
                     _2678,
                     _2658,
                     _2638,
                     _2618,
                     _2598,
                     _2578,
                     _2558,
                     _2538,
                     _2518,
                     _2498,
                     _2478,
                     _2458,
                     _2438,
                     _2418,
                     _2398,
                     _2378,
                     _2358,
                     _2338,
                     _2318,
                     _2298,
                     _2278,
                     _2258,
                     _2238,
                     _2218,
                     _2198,
                     _2178,
                     _2158,
                     _2138,
                     _2118,
                     _2098,
                     _2078,
                     _2058,
                     _2038,
                     _2018,
                     _1998,
                     _1978,
                     _1958,
                     _1938,
                     _1918,
                     _1898,
                     _1878,
                     _1858,
                     _1838,
                     _1818,
                     _1798,
                     _1778,
                     _1758,
                     _1738,
                     _1718,
                     _1698,
                     _1678,
                     _1658,
                     _1638,
                     _1618,
                     _1598,
                     _1578,
                     _1558,
                     _1538,
                     _1518,
                     _1498,
                     _1478,
                     _1458,
                     _1438,
                     _1418,
                     _1398,
                     _1378,
                     _1358,
                     _1338,
                     _1318,
                     _1298,
                     _1278,
                     _1258,
                     _1238,
                     _1218,
                     _1198,
                     _1178,
                     _1158,
                     _1138,
                     _1118,
                     _1098,
                     _1078,
                     _1058,
                     _1038,
                     _1018,
                     _998,
                     _978,
                     _958,
                     _938,
                     _918,
                     _898,
                     _878,
                     _858,
                     _838,
                     _818,
                     _798,
                     _778,
                     _758,
                     _738,
                     _718,
                     _698,
                     _678,
                     _658,
                     _638,
                     _618,
                     _598,
                     _578,
                     _558,
                     _538,
                     _518,
                     _498,
                     _478,
                     _458,
                     _438,
                     _418,
                     _398,
                     _378,
                     _358,
                     _338,
                     _319,
                     _306 };
    assign _7221 = _7220[255:255];
    assign _7222 = { _8232,
                     _7221 };
    assign _7226 = _7222 + _7225;
    assign _7234 = _7226 + _7233;
    assign _7250 = _7234 + _7249;
    assign _7282 = _7250 + _7281;
    assign _7346 = _7282 + _7345;
    assign _7474 = _7346 + _7473;
    assign _7730 = _7474 + _7729;
    assign _8242 = _7730 + _8241;
    assign _7218 = 55'b0000000000000000000000000000000000000000000000000000000;
    assign _8243 = { _7218,
                     _8242 };
    assign _8244 = _7217 + _8243;
    assign _8245 = _287 ? _8244 : _7217;
    assign _8247 = _278 ? _290 : _8245;
    assign _266 = _8247;
    always @(posedge _272) begin
        if (_270)
            _7217 <= _290;
        else
            _7217 <= _266;
    end
    assign _8249 = _284 == _8248;
    assign vdd = 1'b1;
    assign _282 = 2'b00;
    assign _270 = clear;
    assign _272 = clock;
    assign _8248 = 2'b01;
    assign _274 = row_last;
    assign _276 = row_valid;
    assign _287 = _286 & _276;
    assign _8250 = _287 & _274;
    assign _8251 = _8250 ? _8248 : _284;
    assign _278 = load;
    assign _8252 = _278 ? _282 : _8251;
    assign _279 = _8252;
    always @(posedge _272) begin
        if (_270)
            _284 <= _282;
        else
            _284 <= _279;
    end
    assign _286 = _284 == _282;
    assign ready = _286;
    assign done_ = _8249;
    assign part1_result = _7217;
    assign part2_result = _291;
    assign state = _284;

endmodule
