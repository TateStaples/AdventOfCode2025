module day9_opt_b (
    y,
    x,
    clear,
    clock,
    tile_last,
    tile_valid,
    load,
    ready,
    done_,
    part1_result,
    part2_result,
    state
);

    input [63:0] y;
    input [63:0] x;
    input clear;
    input clock;
    input tile_last;
    input tile_valid;
    input load;
    output ready;
    output done_;
    output [63:0] part1_result;
    output [63:0] part2_result;
    output [1:0] state;

    wire [63:0] _1055;
    wire [63:0] _10319;
    wire _10317;
    wire [63:0] _10321;
    wire [63:0] _10311;
    wire [63:0] _10309;
    wire [63:0] _10308;
    reg [63:0] _10305;
    wire [8:0] _1063;
    wire _1064;
    wire _1065;
    wire [63:0] _1069;
    wire [63:0] _1071;
    wire [63:0] _3;
    reg [63:0] _1068;
    wire [8:0] _1072;
    wire _1073;
    wire _1074;
    wire [63:0] _1078;
    wire [63:0] _1080;
    wire [63:0] _4;
    reg [63:0] _1077;
    wire [8:0] _1081;
    wire _1082;
    wire _1083;
    wire [63:0] _1087;
    wire [63:0] _1089;
    wire [63:0] _5;
    reg [63:0] _1086;
    wire [8:0] _1090;
    wire _1091;
    wire _1092;
    wire [63:0] _1096;
    wire [63:0] _1098;
    wire [63:0] _6;
    reg [63:0] _1095;
    wire [8:0] _1099;
    wire _1100;
    wire _1101;
    wire [63:0] _1105;
    wire [63:0] _1107;
    wire [63:0] _7;
    reg [63:0] _1104;
    wire [8:0] _1108;
    wire _1109;
    wire _1110;
    wire [63:0] _1114;
    wire [63:0] _1116;
    wire [63:0] _8;
    reg [63:0] _1113;
    wire [8:0] _1117;
    wire _1118;
    wire _1119;
    wire [63:0] _1123;
    wire [63:0] _1125;
    wire [63:0] _9;
    reg [63:0] _1122;
    wire [8:0] _1126;
    wire _1127;
    wire _1128;
    wire [63:0] _1132;
    wire [63:0] _1134;
    wire [63:0] _10;
    reg [63:0] _1131;
    wire [8:0] _1135;
    wire _1136;
    wire _1137;
    wire [63:0] _1141;
    wire [63:0] _1143;
    wire [63:0] _11;
    reg [63:0] _1140;
    wire [8:0] _1144;
    wire _1145;
    wire _1146;
    wire [63:0] _1150;
    wire [63:0] _1152;
    wire [63:0] _12;
    reg [63:0] _1149;
    wire [8:0] _1153;
    wire _1154;
    wire _1155;
    wire [63:0] _1159;
    wire [63:0] _1161;
    wire [63:0] _13;
    reg [63:0] _1158;
    wire [8:0] _1162;
    wire _1163;
    wire _1164;
    wire [63:0] _1168;
    wire [63:0] _1170;
    wire [63:0] _14;
    reg [63:0] _1167;
    wire [8:0] _1171;
    wire _1172;
    wire _1173;
    wire [63:0] _1177;
    wire [63:0] _1179;
    wire [63:0] _15;
    reg [63:0] _1176;
    wire [8:0] _1180;
    wire _1181;
    wire _1182;
    wire [63:0] _1186;
    wire [63:0] _1188;
    wire [63:0] _16;
    reg [63:0] _1185;
    wire [8:0] _1189;
    wire _1190;
    wire _1191;
    wire [63:0] _1195;
    wire [63:0] _1197;
    wire [63:0] _17;
    reg [63:0] _1194;
    wire [8:0] _1198;
    wire _1199;
    wire _1200;
    wire [63:0] _1204;
    wire [63:0] _1206;
    wire [63:0] _18;
    reg [63:0] _1203;
    wire [8:0] _1207;
    wire _1208;
    wire _1209;
    wire [63:0] _1213;
    wire [63:0] _1215;
    wire [63:0] _19;
    reg [63:0] _1212;
    wire [8:0] _1216;
    wire _1217;
    wire _1218;
    wire [63:0] _1222;
    wire [63:0] _1224;
    wire [63:0] _20;
    reg [63:0] _1221;
    wire [8:0] _1225;
    wire _1226;
    wire _1227;
    wire [63:0] _1231;
    wire [63:0] _1233;
    wire [63:0] _21;
    reg [63:0] _1230;
    wire [8:0] _1234;
    wire _1235;
    wire _1236;
    wire [63:0] _1240;
    wire [63:0] _1242;
    wire [63:0] _22;
    reg [63:0] _1239;
    wire [8:0] _1243;
    wire _1244;
    wire _1245;
    wire [63:0] _1249;
    wire [63:0] _1251;
    wire [63:0] _23;
    reg [63:0] _1248;
    wire [8:0] _1252;
    wire _1253;
    wire _1254;
    wire [63:0] _1258;
    wire [63:0] _1260;
    wire [63:0] _24;
    reg [63:0] _1257;
    wire [8:0] _1261;
    wire _1262;
    wire _1263;
    wire [63:0] _1267;
    wire [63:0] _1269;
    wire [63:0] _25;
    reg [63:0] _1266;
    wire [8:0] _1270;
    wire _1271;
    wire _1272;
    wire [63:0] _1276;
    wire [63:0] _1278;
    wire [63:0] _26;
    reg [63:0] _1275;
    wire [8:0] _1279;
    wire _1280;
    wire _1281;
    wire [63:0] _1285;
    wire [63:0] _1287;
    wire [63:0] _27;
    reg [63:0] _1284;
    wire [8:0] _1288;
    wire _1289;
    wire _1290;
    wire [63:0] _1294;
    wire [63:0] _1296;
    wire [63:0] _28;
    reg [63:0] _1293;
    wire [8:0] _1297;
    wire _1298;
    wire _1299;
    wire [63:0] _1303;
    wire [63:0] _1305;
    wire [63:0] _29;
    reg [63:0] _1302;
    wire [8:0] _1306;
    wire _1307;
    wire _1308;
    wire [63:0] _1312;
    wire [63:0] _1314;
    wire [63:0] _30;
    reg [63:0] _1311;
    wire [8:0] _1315;
    wire _1316;
    wire _1317;
    wire [63:0] _1321;
    wire [63:0] _1323;
    wire [63:0] _31;
    reg [63:0] _1320;
    wire [8:0] _1324;
    wire _1325;
    wire _1326;
    wire [63:0] _1330;
    wire [63:0] _1332;
    wire [63:0] _32;
    reg [63:0] _1329;
    wire [8:0] _1333;
    wire _1334;
    wire _1335;
    wire [63:0] _1339;
    wire [63:0] _1341;
    wire [63:0] _33;
    reg [63:0] _1338;
    wire [8:0] _1342;
    wire _1343;
    wire _1344;
    wire [63:0] _1348;
    wire [63:0] _1350;
    wire [63:0] _34;
    reg [63:0] _1347;
    wire [8:0] _1351;
    wire _1352;
    wire _1353;
    wire [63:0] _1357;
    wire [63:0] _1359;
    wire [63:0] _35;
    reg [63:0] _1356;
    wire [8:0] _1360;
    wire _1361;
    wire _1362;
    wire [63:0] _1366;
    wire [63:0] _1368;
    wire [63:0] _36;
    reg [63:0] _1365;
    wire [8:0] _1369;
    wire _1370;
    wire _1371;
    wire [63:0] _1375;
    wire [63:0] _1377;
    wire [63:0] _37;
    reg [63:0] _1374;
    wire [8:0] _1378;
    wire _1379;
    wire _1380;
    wire [63:0] _1384;
    wire [63:0] _1386;
    wire [63:0] _38;
    reg [63:0] _1383;
    wire [8:0] _1387;
    wire _1388;
    wire _1389;
    wire [63:0] _1393;
    wire [63:0] _1395;
    wire [63:0] _39;
    reg [63:0] _1392;
    wire [8:0] _1396;
    wire _1397;
    wire _1398;
    wire [63:0] _1402;
    wire [63:0] _1404;
    wire [63:0] _40;
    reg [63:0] _1401;
    wire [8:0] _1405;
    wire _1406;
    wire _1407;
    wire [63:0] _1411;
    wire [63:0] _1413;
    wire [63:0] _41;
    reg [63:0] _1410;
    wire [8:0] _1414;
    wire _1415;
    wire _1416;
    wire [63:0] _1420;
    wire [63:0] _1422;
    wire [63:0] _42;
    reg [63:0] _1419;
    wire [8:0] _1423;
    wire _1424;
    wire _1425;
    wire [63:0] _1429;
    wire [63:0] _1431;
    wire [63:0] _43;
    reg [63:0] _1428;
    wire [8:0] _1432;
    wire _1433;
    wire _1434;
    wire [63:0] _1438;
    wire [63:0] _1440;
    wire [63:0] _44;
    reg [63:0] _1437;
    wire [8:0] _1441;
    wire _1442;
    wire _1443;
    wire [63:0] _1447;
    wire [63:0] _1449;
    wire [63:0] _45;
    reg [63:0] _1446;
    wire [8:0] _1450;
    wire _1451;
    wire _1452;
    wire [63:0] _1456;
    wire [63:0] _1458;
    wire [63:0] _46;
    reg [63:0] _1455;
    wire [8:0] _1459;
    wire _1460;
    wire _1461;
    wire [63:0] _1465;
    wire [63:0] _1467;
    wire [63:0] _47;
    reg [63:0] _1464;
    wire [8:0] _1468;
    wire _1469;
    wire _1470;
    wire [63:0] _1474;
    wire [63:0] _1476;
    wire [63:0] _48;
    reg [63:0] _1473;
    wire [8:0] _1477;
    wire _1478;
    wire _1479;
    wire [63:0] _1483;
    wire [63:0] _1485;
    wire [63:0] _49;
    reg [63:0] _1482;
    wire [8:0] _1486;
    wire _1487;
    wire _1488;
    wire [63:0] _1492;
    wire [63:0] _1494;
    wire [63:0] _50;
    reg [63:0] _1491;
    wire [8:0] _1495;
    wire _1496;
    wire _1497;
    wire [63:0] _1501;
    wire [63:0] _1503;
    wire [63:0] _51;
    reg [63:0] _1500;
    wire [8:0] _1504;
    wire _1505;
    wire _1506;
    wire [63:0] _1510;
    wire [63:0] _1512;
    wire [63:0] _52;
    reg [63:0] _1509;
    wire [8:0] _1513;
    wire _1514;
    wire _1515;
    wire [63:0] _1519;
    wire [63:0] _1521;
    wire [63:0] _53;
    reg [63:0] _1518;
    wire [8:0] _1522;
    wire _1523;
    wire _1524;
    wire [63:0] _1528;
    wire [63:0] _1530;
    wire [63:0] _54;
    reg [63:0] _1527;
    wire [8:0] _1531;
    wire _1532;
    wire _1533;
    wire [63:0] _1537;
    wire [63:0] _1539;
    wire [63:0] _55;
    reg [63:0] _1536;
    wire [8:0] _1540;
    wire _1541;
    wire _1542;
    wire [63:0] _1546;
    wire [63:0] _1548;
    wire [63:0] _56;
    reg [63:0] _1545;
    wire [8:0] _1549;
    wire _1550;
    wire _1551;
    wire [63:0] _1555;
    wire [63:0] _1557;
    wire [63:0] _57;
    reg [63:0] _1554;
    wire [8:0] _1558;
    wire _1559;
    wire _1560;
    wire [63:0] _1564;
    wire [63:0] _1566;
    wire [63:0] _58;
    reg [63:0] _1563;
    wire [8:0] _1567;
    wire _1568;
    wire _1569;
    wire [63:0] _1573;
    wire [63:0] _1575;
    wire [63:0] _59;
    reg [63:0] _1572;
    wire [8:0] _1576;
    wire _1577;
    wire _1578;
    wire [63:0] _1582;
    wire [63:0] _1584;
    wire [63:0] _60;
    reg [63:0] _1581;
    wire [8:0] _1585;
    wire _1586;
    wire _1587;
    wire [63:0] _1591;
    wire [63:0] _1593;
    wire [63:0] _61;
    reg [63:0] _1590;
    wire [8:0] _1594;
    wire _1595;
    wire _1596;
    wire [63:0] _1600;
    wire [63:0] _1602;
    wire [63:0] _62;
    reg [63:0] _1599;
    wire [8:0] _1603;
    wire _1604;
    wire _1605;
    wire [63:0] _1609;
    wire [63:0] _1611;
    wire [63:0] _63;
    reg [63:0] _1608;
    wire [8:0] _1612;
    wire _1613;
    wire _1614;
    wire [63:0] _1618;
    wire [63:0] _1620;
    wire [63:0] _64;
    reg [63:0] _1617;
    wire [8:0] _1621;
    wire _1622;
    wire _1623;
    wire [63:0] _1627;
    wire [63:0] _1629;
    wire [63:0] _65;
    reg [63:0] _1626;
    wire [8:0] _1630;
    wire _1631;
    wire _1632;
    wire [63:0] _1636;
    wire [63:0] _1638;
    wire [63:0] _66;
    reg [63:0] _1635;
    wire [8:0] _1639;
    wire _1640;
    wire _1641;
    wire [63:0] _1645;
    wire [63:0] _1647;
    wire [63:0] _67;
    reg [63:0] _1644;
    wire [8:0] _1648;
    wire _1649;
    wire _1650;
    wire [63:0] _1654;
    wire [63:0] _1656;
    wire [63:0] _68;
    reg [63:0] _1653;
    wire [8:0] _1657;
    wire _1658;
    wire _1659;
    wire [63:0] _1663;
    wire [63:0] _1665;
    wire [63:0] _69;
    reg [63:0] _1662;
    wire [8:0] _1666;
    wire _1667;
    wire _1668;
    wire [63:0] _1672;
    wire [63:0] _1674;
    wire [63:0] _70;
    reg [63:0] _1671;
    wire [8:0] _1675;
    wire _1676;
    wire _1677;
    wire [63:0] _1681;
    wire [63:0] _1683;
    wire [63:0] _71;
    reg [63:0] _1680;
    wire [8:0] _1684;
    wire _1685;
    wire _1686;
    wire [63:0] _1690;
    wire [63:0] _1692;
    wire [63:0] _72;
    reg [63:0] _1689;
    wire [8:0] _1693;
    wire _1694;
    wire _1695;
    wire [63:0] _1699;
    wire [63:0] _1701;
    wire [63:0] _73;
    reg [63:0] _1698;
    wire [8:0] _1702;
    wire _1703;
    wire _1704;
    wire [63:0] _1708;
    wire [63:0] _1710;
    wire [63:0] _74;
    reg [63:0] _1707;
    wire [8:0] _1711;
    wire _1712;
    wire _1713;
    wire [63:0] _1717;
    wire [63:0] _1719;
    wire [63:0] _75;
    reg [63:0] _1716;
    wire [8:0] _1720;
    wire _1721;
    wire _1722;
    wire [63:0] _1726;
    wire [63:0] _1728;
    wire [63:0] _76;
    reg [63:0] _1725;
    wire [8:0] _1729;
    wire _1730;
    wire _1731;
    wire [63:0] _1735;
    wire [63:0] _1737;
    wire [63:0] _77;
    reg [63:0] _1734;
    wire [8:0] _1738;
    wire _1739;
    wire _1740;
    wire [63:0] _1744;
    wire [63:0] _1746;
    wire [63:0] _78;
    reg [63:0] _1743;
    wire [8:0] _1747;
    wire _1748;
    wire _1749;
    wire [63:0] _1753;
    wire [63:0] _1755;
    wire [63:0] _79;
    reg [63:0] _1752;
    wire [8:0] _1756;
    wire _1757;
    wire _1758;
    wire [63:0] _1762;
    wire [63:0] _1764;
    wire [63:0] _80;
    reg [63:0] _1761;
    wire [8:0] _1765;
    wire _1766;
    wire _1767;
    wire [63:0] _1771;
    wire [63:0] _1773;
    wire [63:0] _81;
    reg [63:0] _1770;
    wire [8:0] _1774;
    wire _1775;
    wire _1776;
    wire [63:0] _1780;
    wire [63:0] _1782;
    wire [63:0] _82;
    reg [63:0] _1779;
    wire [8:0] _1783;
    wire _1784;
    wire _1785;
    wire [63:0] _1789;
    wire [63:0] _1791;
    wire [63:0] _83;
    reg [63:0] _1788;
    wire [8:0] _1792;
    wire _1793;
    wire _1794;
    wire [63:0] _1798;
    wire [63:0] _1800;
    wire [63:0] _84;
    reg [63:0] _1797;
    wire [8:0] _1801;
    wire _1802;
    wire _1803;
    wire [63:0] _1807;
    wire [63:0] _1809;
    wire [63:0] _85;
    reg [63:0] _1806;
    wire [8:0] _1810;
    wire _1811;
    wire _1812;
    wire [63:0] _1816;
    wire [63:0] _1818;
    wire [63:0] _86;
    reg [63:0] _1815;
    wire [8:0] _1819;
    wire _1820;
    wire _1821;
    wire [63:0] _1825;
    wire [63:0] _1827;
    wire [63:0] _87;
    reg [63:0] _1824;
    wire [8:0] _1828;
    wire _1829;
    wire _1830;
    wire [63:0] _1834;
    wire [63:0] _1836;
    wire [63:0] _88;
    reg [63:0] _1833;
    wire [8:0] _1837;
    wire _1838;
    wire _1839;
    wire [63:0] _1843;
    wire [63:0] _1845;
    wire [63:0] _89;
    reg [63:0] _1842;
    wire [8:0] _1846;
    wire _1847;
    wire _1848;
    wire [63:0] _1852;
    wire [63:0] _1854;
    wire [63:0] _90;
    reg [63:0] _1851;
    wire [8:0] _1855;
    wire _1856;
    wire _1857;
    wire [63:0] _1861;
    wire [63:0] _1863;
    wire [63:0] _91;
    reg [63:0] _1860;
    wire [8:0] _1864;
    wire _1865;
    wire _1866;
    wire [63:0] _1870;
    wire [63:0] _1872;
    wire [63:0] _92;
    reg [63:0] _1869;
    wire [8:0] _1873;
    wire _1874;
    wire _1875;
    wire [63:0] _1879;
    wire [63:0] _1881;
    wire [63:0] _93;
    reg [63:0] _1878;
    wire [8:0] _1882;
    wire _1883;
    wire _1884;
    wire [63:0] _1888;
    wire [63:0] _1890;
    wire [63:0] _94;
    reg [63:0] _1887;
    wire [8:0] _1891;
    wire _1892;
    wire _1893;
    wire [63:0] _1897;
    wire [63:0] _1899;
    wire [63:0] _95;
    reg [63:0] _1896;
    wire [8:0] _1900;
    wire _1901;
    wire _1902;
    wire [63:0] _1906;
    wire [63:0] _1908;
    wire [63:0] _96;
    reg [63:0] _1905;
    wire [8:0] _1909;
    wire _1910;
    wire _1911;
    wire [63:0] _1915;
    wire [63:0] _1917;
    wire [63:0] _97;
    reg [63:0] _1914;
    wire [8:0] _1918;
    wire _1919;
    wire _1920;
    wire [63:0] _1924;
    wire [63:0] _1926;
    wire [63:0] _98;
    reg [63:0] _1923;
    wire [8:0] _1927;
    wire _1928;
    wire _1929;
    wire [63:0] _1933;
    wire [63:0] _1935;
    wire [63:0] _99;
    reg [63:0] _1932;
    wire [8:0] _1936;
    wire _1937;
    wire _1938;
    wire [63:0] _1942;
    wire [63:0] _1944;
    wire [63:0] _100;
    reg [63:0] _1941;
    wire [8:0] _1945;
    wire _1946;
    wire _1947;
    wire [63:0] _1951;
    wire [63:0] _1953;
    wire [63:0] _101;
    reg [63:0] _1950;
    wire [8:0] _1954;
    wire _1955;
    wire _1956;
    wire [63:0] _1960;
    wire [63:0] _1962;
    wire [63:0] _102;
    reg [63:0] _1959;
    wire [8:0] _1963;
    wire _1964;
    wire _1965;
    wire [63:0] _1969;
    wire [63:0] _1971;
    wire [63:0] _103;
    reg [63:0] _1968;
    wire [8:0] _1972;
    wire _1973;
    wire _1974;
    wire [63:0] _1978;
    wire [63:0] _1980;
    wire [63:0] _104;
    reg [63:0] _1977;
    wire [8:0] _1981;
    wire _1982;
    wire _1983;
    wire [63:0] _1987;
    wire [63:0] _1989;
    wire [63:0] _105;
    reg [63:0] _1986;
    wire [8:0] _1990;
    wire _1991;
    wire _1992;
    wire [63:0] _1996;
    wire [63:0] _1998;
    wire [63:0] _106;
    reg [63:0] _1995;
    wire [8:0] _1999;
    wire _2000;
    wire _2001;
    wire [63:0] _2005;
    wire [63:0] _2007;
    wire [63:0] _107;
    reg [63:0] _2004;
    wire [8:0] _2008;
    wire _2009;
    wire _2010;
    wire [63:0] _2014;
    wire [63:0] _2016;
    wire [63:0] _108;
    reg [63:0] _2013;
    wire [8:0] _2017;
    wire _2018;
    wire _2019;
    wire [63:0] _2023;
    wire [63:0] _2025;
    wire [63:0] _109;
    reg [63:0] _2022;
    wire [8:0] _2026;
    wire _2027;
    wire _2028;
    wire [63:0] _2032;
    wire [63:0] _2034;
    wire [63:0] _110;
    reg [63:0] _2031;
    wire [8:0] _2035;
    wire _2036;
    wire _2037;
    wire [63:0] _2041;
    wire [63:0] _2043;
    wire [63:0] _111;
    reg [63:0] _2040;
    wire [8:0] _2044;
    wire _2045;
    wire _2046;
    wire [63:0] _2050;
    wire [63:0] _2052;
    wire [63:0] _112;
    reg [63:0] _2049;
    wire [8:0] _2053;
    wire _2054;
    wire _2055;
    wire [63:0] _2059;
    wire [63:0] _2061;
    wire [63:0] _113;
    reg [63:0] _2058;
    wire [8:0] _2062;
    wire _2063;
    wire _2064;
    wire [63:0] _2068;
    wire [63:0] _2070;
    wire [63:0] _114;
    reg [63:0] _2067;
    wire [8:0] _2071;
    wire _2072;
    wire _2073;
    wire [63:0] _2077;
    wire [63:0] _2079;
    wire [63:0] _115;
    reg [63:0] _2076;
    wire [8:0] _2080;
    wire _2081;
    wire _2082;
    wire [63:0] _2086;
    wire [63:0] _2088;
    wire [63:0] _116;
    reg [63:0] _2085;
    wire [8:0] _2089;
    wire _2090;
    wire _2091;
    wire [63:0] _2095;
    wire [63:0] _2097;
    wire [63:0] _117;
    reg [63:0] _2094;
    wire [8:0] _2098;
    wire _2099;
    wire _2100;
    wire [63:0] _2104;
    wire [63:0] _2106;
    wire [63:0] _118;
    reg [63:0] _2103;
    wire [8:0] _2107;
    wire _2108;
    wire _2109;
    wire [63:0] _2113;
    wire [63:0] _2115;
    wire [63:0] _119;
    reg [63:0] _2112;
    wire [8:0] _2116;
    wire _2117;
    wire _2118;
    wire [63:0] _2122;
    wire [63:0] _2124;
    wire [63:0] _120;
    reg [63:0] _2121;
    wire [8:0] _2125;
    wire _2126;
    wire _2127;
    wire [63:0] _2131;
    wire [63:0] _2133;
    wire [63:0] _121;
    reg [63:0] _2130;
    wire [8:0] _2134;
    wire _2135;
    wire _2136;
    wire [63:0] _2140;
    wire [63:0] _2142;
    wire [63:0] _122;
    reg [63:0] _2139;
    wire [8:0] _2143;
    wire _2144;
    wire _2145;
    wire [63:0] _2149;
    wire [63:0] _2151;
    wire [63:0] _123;
    reg [63:0] _2148;
    wire [8:0] _2152;
    wire _2153;
    wire _2154;
    wire [63:0] _2158;
    wire [63:0] _2160;
    wire [63:0] _124;
    reg [63:0] _2157;
    wire [8:0] _2161;
    wire _2162;
    wire _2163;
    wire [63:0] _2167;
    wire [63:0] _2169;
    wire [63:0] _125;
    reg [63:0] _2166;
    wire [8:0] _2170;
    wire _2171;
    wire _2172;
    wire [63:0] _2176;
    wire [63:0] _2178;
    wire [63:0] _126;
    reg [63:0] _2175;
    wire [8:0] _2179;
    wire _2180;
    wire _2181;
    wire [63:0] _2185;
    wire [63:0] _2187;
    wire [63:0] _127;
    reg [63:0] _2184;
    wire [8:0] _2188;
    wire _2189;
    wire _2190;
    wire [63:0] _2194;
    wire [63:0] _2196;
    wire [63:0] _128;
    reg [63:0] _2193;
    wire [8:0] _2197;
    wire _2198;
    wire _2199;
    wire [63:0] _2203;
    wire [63:0] _2205;
    wire [63:0] _129;
    reg [63:0] _2202;
    wire [8:0] _2206;
    wire _2207;
    wire _2208;
    wire [63:0] _2212;
    wire [63:0] _2214;
    wire [63:0] _130;
    reg [63:0] _2211;
    wire [8:0] _2215;
    wire _2216;
    wire _2217;
    wire [63:0] _2221;
    wire [63:0] _2223;
    wire [63:0] _131;
    reg [63:0] _2220;
    wire [8:0] _2224;
    wire _2225;
    wire _2226;
    wire [63:0] _2230;
    wire [63:0] _2232;
    wire [63:0] _132;
    reg [63:0] _2229;
    wire [8:0] _2233;
    wire _2234;
    wire _2235;
    wire [63:0] _2239;
    wire [63:0] _2241;
    wire [63:0] _133;
    reg [63:0] _2238;
    wire [8:0] _2242;
    wire _2243;
    wire _2244;
    wire [63:0] _2248;
    wire [63:0] _2250;
    wire [63:0] _134;
    reg [63:0] _2247;
    wire [8:0] _2251;
    wire _2252;
    wire _2253;
    wire [63:0] _2257;
    wire [63:0] _2259;
    wire [63:0] _135;
    reg [63:0] _2256;
    wire [8:0] _2260;
    wire _2261;
    wire _2262;
    wire [63:0] _2266;
    wire [63:0] _2268;
    wire [63:0] _136;
    reg [63:0] _2265;
    wire [8:0] _2269;
    wire _2270;
    wire _2271;
    wire [63:0] _2275;
    wire [63:0] _2277;
    wire [63:0] _137;
    reg [63:0] _2274;
    wire [8:0] _2278;
    wire _2279;
    wire _2280;
    wire [63:0] _2284;
    wire [63:0] _2286;
    wire [63:0] _138;
    reg [63:0] _2283;
    wire [8:0] _2287;
    wire _2288;
    wire _2289;
    wire [63:0] _2293;
    wire [63:0] _2295;
    wire [63:0] _139;
    reg [63:0] _2292;
    wire [8:0] _2296;
    wire _2297;
    wire _2298;
    wire [63:0] _2302;
    wire [63:0] _2304;
    wire [63:0] _140;
    reg [63:0] _2301;
    wire [8:0] _2305;
    wire _2306;
    wire _2307;
    wire [63:0] _2311;
    wire [63:0] _2313;
    wire [63:0] _141;
    reg [63:0] _2310;
    wire [8:0] _2314;
    wire _2315;
    wire _2316;
    wire [63:0] _2320;
    wire [63:0] _2322;
    wire [63:0] _142;
    reg [63:0] _2319;
    wire [8:0] _2323;
    wire _2324;
    wire _2325;
    wire [63:0] _2329;
    wire [63:0] _2331;
    wire [63:0] _143;
    reg [63:0] _2328;
    wire [8:0] _2332;
    wire _2333;
    wire _2334;
    wire [63:0] _2338;
    wire [63:0] _2340;
    wire [63:0] _144;
    reg [63:0] _2337;
    wire [8:0] _2341;
    wire _2342;
    wire _2343;
    wire [63:0] _2347;
    wire [63:0] _2349;
    wire [63:0] _145;
    reg [63:0] _2346;
    wire [8:0] _2350;
    wire _2351;
    wire _2352;
    wire [63:0] _2356;
    wire [63:0] _2358;
    wire [63:0] _146;
    reg [63:0] _2355;
    wire [8:0] _2359;
    wire _2360;
    wire _2361;
    wire [63:0] _2365;
    wire [63:0] _2367;
    wire [63:0] _147;
    reg [63:0] _2364;
    wire [8:0] _2368;
    wire _2369;
    wire _2370;
    wire [63:0] _2374;
    wire [63:0] _2376;
    wire [63:0] _148;
    reg [63:0] _2373;
    wire [8:0] _2377;
    wire _2378;
    wire _2379;
    wire [63:0] _2383;
    wire [63:0] _2385;
    wire [63:0] _149;
    reg [63:0] _2382;
    wire [8:0] _2386;
    wire _2387;
    wire _2388;
    wire [63:0] _2392;
    wire [63:0] _2394;
    wire [63:0] _150;
    reg [63:0] _2391;
    wire [8:0] _2395;
    wire _2396;
    wire _2397;
    wire [63:0] _2401;
    wire [63:0] _2403;
    wire [63:0] _151;
    reg [63:0] _2400;
    wire [8:0] _2404;
    wire _2405;
    wire _2406;
    wire [63:0] _2410;
    wire [63:0] _2412;
    wire [63:0] _152;
    reg [63:0] _2409;
    wire [8:0] _2413;
    wire _2414;
    wire _2415;
    wire [63:0] _2419;
    wire [63:0] _2421;
    wire [63:0] _153;
    reg [63:0] _2418;
    wire [8:0] _2422;
    wire _2423;
    wire _2424;
    wire [63:0] _2428;
    wire [63:0] _2430;
    wire [63:0] _154;
    reg [63:0] _2427;
    wire [8:0] _2431;
    wire _2432;
    wire _2433;
    wire [63:0] _2437;
    wire [63:0] _2439;
    wire [63:0] _155;
    reg [63:0] _2436;
    wire [8:0] _2440;
    wire _2441;
    wire _2442;
    wire [63:0] _2446;
    wire [63:0] _2448;
    wire [63:0] _156;
    reg [63:0] _2445;
    wire [8:0] _2449;
    wire _2450;
    wire _2451;
    wire [63:0] _2455;
    wire [63:0] _2457;
    wire [63:0] _157;
    reg [63:0] _2454;
    wire [8:0] _2458;
    wire _2459;
    wire _2460;
    wire [63:0] _2464;
    wire [63:0] _2466;
    wire [63:0] _158;
    reg [63:0] _2463;
    wire [8:0] _2467;
    wire _2468;
    wire _2469;
    wire [63:0] _2473;
    wire [63:0] _2475;
    wire [63:0] _159;
    reg [63:0] _2472;
    wire [8:0] _2476;
    wire _2477;
    wire _2478;
    wire [63:0] _2482;
    wire [63:0] _2484;
    wire [63:0] _160;
    reg [63:0] _2481;
    wire [8:0] _2485;
    wire _2486;
    wire _2487;
    wire [63:0] _2491;
    wire [63:0] _2493;
    wire [63:0] _161;
    reg [63:0] _2490;
    wire [8:0] _2494;
    wire _2495;
    wire _2496;
    wire [63:0] _2500;
    wire [63:0] _2502;
    wire [63:0] _162;
    reg [63:0] _2499;
    wire [8:0] _2503;
    wire _2504;
    wire _2505;
    wire [63:0] _2509;
    wire [63:0] _2511;
    wire [63:0] _163;
    reg [63:0] _2508;
    wire [8:0] _2512;
    wire _2513;
    wire _2514;
    wire [63:0] _2518;
    wire [63:0] _2520;
    wire [63:0] _164;
    reg [63:0] _2517;
    wire [8:0] _2521;
    wire _2522;
    wire _2523;
    wire [63:0] _2527;
    wire [63:0] _2529;
    wire [63:0] _165;
    reg [63:0] _2526;
    wire [8:0] _2530;
    wire _2531;
    wire _2532;
    wire [63:0] _2536;
    wire [63:0] _2538;
    wire [63:0] _166;
    reg [63:0] _2535;
    wire [8:0] _2539;
    wire _2540;
    wire _2541;
    wire [63:0] _2545;
    wire [63:0] _2547;
    wire [63:0] _167;
    reg [63:0] _2544;
    wire [8:0] _2548;
    wire _2549;
    wire _2550;
    wire [63:0] _2554;
    wire [63:0] _2556;
    wire [63:0] _168;
    reg [63:0] _2553;
    wire [8:0] _2557;
    wire _2558;
    wire _2559;
    wire [63:0] _2563;
    wire [63:0] _2565;
    wire [63:0] _169;
    reg [63:0] _2562;
    wire [8:0] _2566;
    wire _2567;
    wire _2568;
    wire [63:0] _2572;
    wire [63:0] _2574;
    wire [63:0] _170;
    reg [63:0] _2571;
    wire [8:0] _2575;
    wire _2576;
    wire _2577;
    wire [63:0] _2581;
    wire [63:0] _2583;
    wire [63:0] _171;
    reg [63:0] _2580;
    wire [8:0] _2584;
    wire _2585;
    wire _2586;
    wire [63:0] _2590;
    wire [63:0] _2592;
    wire [63:0] _172;
    reg [63:0] _2589;
    wire [8:0] _2593;
    wire _2594;
    wire _2595;
    wire [63:0] _2599;
    wire [63:0] _2601;
    wire [63:0] _173;
    reg [63:0] _2598;
    wire [8:0] _2602;
    wire _2603;
    wire _2604;
    wire [63:0] _2608;
    wire [63:0] _2610;
    wire [63:0] _174;
    reg [63:0] _2607;
    wire [8:0] _2611;
    wire _2612;
    wire _2613;
    wire [63:0] _2617;
    wire [63:0] _2619;
    wire [63:0] _175;
    reg [63:0] _2616;
    wire [8:0] _2620;
    wire _2621;
    wire _2622;
    wire [63:0] _2626;
    wire [63:0] _2628;
    wire [63:0] _176;
    reg [63:0] _2625;
    wire [8:0] _2629;
    wire _2630;
    wire _2631;
    wire [63:0] _2635;
    wire [63:0] _2637;
    wire [63:0] _177;
    reg [63:0] _2634;
    wire [8:0] _2638;
    wire _2639;
    wire _2640;
    wire [63:0] _2644;
    wire [63:0] _2646;
    wire [63:0] _178;
    reg [63:0] _2643;
    wire [8:0] _2647;
    wire _2648;
    wire _2649;
    wire [63:0] _2653;
    wire [63:0] _2655;
    wire [63:0] _179;
    reg [63:0] _2652;
    wire [8:0] _2656;
    wire _2657;
    wire _2658;
    wire [63:0] _2662;
    wire [63:0] _2664;
    wire [63:0] _180;
    reg [63:0] _2661;
    wire [8:0] _2665;
    wire _2666;
    wire _2667;
    wire [63:0] _2671;
    wire [63:0] _2673;
    wire [63:0] _181;
    reg [63:0] _2670;
    wire [8:0] _2674;
    wire _2675;
    wire _2676;
    wire [63:0] _2680;
    wire [63:0] _2682;
    wire [63:0] _182;
    reg [63:0] _2679;
    wire [8:0] _2683;
    wire _2684;
    wire _2685;
    wire [63:0] _2689;
    wire [63:0] _2691;
    wire [63:0] _183;
    reg [63:0] _2688;
    wire [8:0] _2692;
    wire _2693;
    wire _2694;
    wire [63:0] _2698;
    wire [63:0] _2700;
    wire [63:0] _184;
    reg [63:0] _2697;
    wire [8:0] _2701;
    wire _2702;
    wire _2703;
    wire [63:0] _2707;
    wire [63:0] _2709;
    wire [63:0] _185;
    reg [63:0] _2706;
    wire [8:0] _2710;
    wire _2711;
    wire _2712;
    wire [63:0] _2716;
    wire [63:0] _2718;
    wire [63:0] _186;
    reg [63:0] _2715;
    wire [8:0] _2719;
    wire _2720;
    wire _2721;
    wire [63:0] _2725;
    wire [63:0] _2727;
    wire [63:0] _187;
    reg [63:0] _2724;
    wire [8:0] _2728;
    wire _2729;
    wire _2730;
    wire [63:0] _2734;
    wire [63:0] _2736;
    wire [63:0] _188;
    reg [63:0] _2733;
    wire [8:0] _2737;
    wire _2738;
    wire _2739;
    wire [63:0] _2743;
    wire [63:0] _2745;
    wire [63:0] _189;
    reg [63:0] _2742;
    wire [8:0] _2746;
    wire _2747;
    wire _2748;
    wire [63:0] _2752;
    wire [63:0] _2754;
    wire [63:0] _190;
    reg [63:0] _2751;
    wire [8:0] _2755;
    wire _2756;
    wire _2757;
    wire [63:0] _2761;
    wire [63:0] _2763;
    wire [63:0] _191;
    reg [63:0] _2760;
    wire [8:0] _2764;
    wire _2765;
    wire _2766;
    wire [63:0] _2770;
    wire [63:0] _2772;
    wire [63:0] _192;
    reg [63:0] _2769;
    wire [8:0] _2773;
    wire _2774;
    wire _2775;
    wire [63:0] _2779;
    wire [63:0] _2781;
    wire [63:0] _193;
    reg [63:0] _2778;
    wire [8:0] _2782;
    wire _2783;
    wire _2784;
    wire [63:0] _2788;
    wire [63:0] _2790;
    wire [63:0] _194;
    reg [63:0] _2787;
    wire [8:0] _2791;
    wire _2792;
    wire _2793;
    wire [63:0] _2797;
    wire [63:0] _2799;
    wire [63:0] _195;
    reg [63:0] _2796;
    wire [8:0] _2800;
    wire _2801;
    wire _2802;
    wire [63:0] _2806;
    wire [63:0] _2808;
    wire [63:0] _196;
    reg [63:0] _2805;
    wire [8:0] _2809;
    wire _2810;
    wire _2811;
    wire [63:0] _2815;
    wire [63:0] _2817;
    wire [63:0] _197;
    reg [63:0] _2814;
    wire [8:0] _2818;
    wire _2819;
    wire _2820;
    wire [63:0] _2824;
    wire [63:0] _2826;
    wire [63:0] _198;
    reg [63:0] _2823;
    wire [8:0] _2827;
    wire _2828;
    wire _2829;
    wire [63:0] _2833;
    wire [63:0] _2835;
    wire [63:0] _199;
    reg [63:0] _2832;
    wire [8:0] _2836;
    wire _2837;
    wire _2838;
    wire [63:0] _2842;
    wire [63:0] _2844;
    wire [63:0] _200;
    reg [63:0] _2841;
    wire [8:0] _2845;
    wire _2846;
    wire _2847;
    wire [63:0] _2851;
    wire [63:0] _2853;
    wire [63:0] _201;
    reg [63:0] _2850;
    wire [8:0] _2854;
    wire _2855;
    wire _2856;
    wire [63:0] _2860;
    wire [63:0] _2862;
    wire [63:0] _202;
    reg [63:0] _2859;
    wire [8:0] _2863;
    wire _2864;
    wire _2865;
    wire [63:0] _2869;
    wire [63:0] _2871;
    wire [63:0] _203;
    reg [63:0] _2868;
    wire [8:0] _2872;
    wire _2873;
    wire _2874;
    wire [63:0] _2878;
    wire [63:0] _2880;
    wire [63:0] _204;
    reg [63:0] _2877;
    wire [8:0] _2881;
    wire _2882;
    wire _2883;
    wire [63:0] _2887;
    wire [63:0] _2889;
    wire [63:0] _205;
    reg [63:0] _2886;
    wire [8:0] _2890;
    wire _2891;
    wire _2892;
    wire [63:0] _2896;
    wire [63:0] _2898;
    wire [63:0] _206;
    reg [63:0] _2895;
    wire [8:0] _2899;
    wire _2900;
    wire _2901;
    wire [63:0] _2905;
    wire [63:0] _2907;
    wire [63:0] _207;
    reg [63:0] _2904;
    wire [8:0] _2908;
    wire _2909;
    wire _2910;
    wire [63:0] _2914;
    wire [63:0] _2916;
    wire [63:0] _208;
    reg [63:0] _2913;
    wire [8:0] _2917;
    wire _2918;
    wire _2919;
    wire [63:0] _2923;
    wire [63:0] _2925;
    wire [63:0] _209;
    reg [63:0] _2922;
    wire [8:0] _2926;
    wire _2927;
    wire _2928;
    wire [63:0] _2932;
    wire [63:0] _2934;
    wire [63:0] _210;
    reg [63:0] _2931;
    wire [8:0] _2935;
    wire _2936;
    wire _2937;
    wire [63:0] _2941;
    wire [63:0] _2943;
    wire [63:0] _211;
    reg [63:0] _2940;
    wire [8:0] _2944;
    wire _2945;
    wire _2946;
    wire [63:0] _2950;
    wire [63:0] _2952;
    wire [63:0] _212;
    reg [63:0] _2949;
    wire [8:0] _2953;
    wire _2954;
    wire _2955;
    wire [63:0] _2959;
    wire [63:0] _2961;
    wire [63:0] _213;
    reg [63:0] _2958;
    wire [8:0] _2962;
    wire _2963;
    wire _2964;
    wire [63:0] _2968;
    wire [63:0] _2970;
    wire [63:0] _214;
    reg [63:0] _2967;
    wire [8:0] _2971;
    wire _2972;
    wire _2973;
    wire [63:0] _2977;
    wire [63:0] _2979;
    wire [63:0] _215;
    reg [63:0] _2976;
    wire [8:0] _2980;
    wire _2981;
    wire _2982;
    wire [63:0] _2986;
    wire [63:0] _2988;
    wire [63:0] _216;
    reg [63:0] _2985;
    wire [8:0] _2989;
    wire _2990;
    wire _2991;
    wire [63:0] _2995;
    wire [63:0] _2997;
    wire [63:0] _217;
    reg [63:0] _2994;
    wire [8:0] _2998;
    wire _2999;
    wire _3000;
    wire [63:0] _3004;
    wire [63:0] _3006;
    wire [63:0] _218;
    reg [63:0] _3003;
    wire [8:0] _3007;
    wire _3008;
    wire _3009;
    wire [63:0] _3013;
    wire [63:0] _3015;
    wire [63:0] _219;
    reg [63:0] _3012;
    wire [8:0] _3016;
    wire _3017;
    wire _3018;
    wire [63:0] _3022;
    wire [63:0] _3024;
    wire [63:0] _220;
    reg [63:0] _3021;
    wire [8:0] _3025;
    wire _3026;
    wire _3027;
    wire [63:0] _3031;
    wire [63:0] _3033;
    wire [63:0] _221;
    reg [63:0] _3030;
    wire [8:0] _3034;
    wire _3035;
    wire _3036;
    wire [63:0] _3040;
    wire [63:0] _3042;
    wire [63:0] _222;
    reg [63:0] _3039;
    wire [8:0] _3043;
    wire _3044;
    wire _3045;
    wire [63:0] _3049;
    wire [63:0] _3051;
    wire [63:0] _223;
    reg [63:0] _3048;
    wire [8:0] _3052;
    wire _3053;
    wire _3054;
    wire [63:0] _3058;
    wire [63:0] _3060;
    wire [63:0] _224;
    reg [63:0] _3057;
    wire [8:0] _3061;
    wire _3062;
    wire _3063;
    wire [63:0] _3067;
    wire [63:0] _3069;
    wire [63:0] _225;
    reg [63:0] _3066;
    wire [8:0] _3070;
    wire _3071;
    wire _3072;
    wire [63:0] _3076;
    wire [63:0] _3078;
    wire [63:0] _226;
    reg [63:0] _3075;
    wire [8:0] _3079;
    wire _3080;
    wire _3081;
    wire [63:0] _3085;
    wire [63:0] _3087;
    wire [63:0] _227;
    reg [63:0] _3084;
    wire [8:0] _3088;
    wire _3089;
    wire _3090;
    wire [63:0] _3094;
    wire [63:0] _3096;
    wire [63:0] _228;
    reg [63:0] _3093;
    wire [8:0] _3097;
    wire _3098;
    wire _3099;
    wire [63:0] _3103;
    wire [63:0] _3105;
    wire [63:0] _229;
    reg [63:0] _3102;
    wire [8:0] _3106;
    wire _3107;
    wire _3108;
    wire [63:0] _3112;
    wire [63:0] _3114;
    wire [63:0] _230;
    reg [63:0] _3111;
    wire [8:0] _3115;
    wire _3116;
    wire _3117;
    wire [63:0] _3121;
    wire [63:0] _3123;
    wire [63:0] _231;
    reg [63:0] _3120;
    wire [8:0] _3124;
    wire _3125;
    wire _3126;
    wire [63:0] _3130;
    wire [63:0] _3132;
    wire [63:0] _232;
    reg [63:0] _3129;
    wire [8:0] _3133;
    wire _3134;
    wire _3135;
    wire [63:0] _3139;
    wire [63:0] _3141;
    wire [63:0] _233;
    reg [63:0] _3138;
    wire [8:0] _3142;
    wire _3143;
    wire _3144;
    wire [63:0] _3148;
    wire [63:0] _3150;
    wire [63:0] _234;
    reg [63:0] _3147;
    wire [8:0] _3151;
    wire _3152;
    wire _3153;
    wire [63:0] _3157;
    wire [63:0] _3159;
    wire [63:0] _235;
    reg [63:0] _3156;
    wire [8:0] _3160;
    wire _3161;
    wire _3162;
    wire [63:0] _3166;
    wire [63:0] _3168;
    wire [63:0] _236;
    reg [63:0] _3165;
    wire [8:0] _3169;
    wire _3170;
    wire _3171;
    wire [63:0] _3175;
    wire [63:0] _3177;
    wire [63:0] _237;
    reg [63:0] _3174;
    wire [8:0] _3178;
    wire _3179;
    wire _3180;
    wire [63:0] _3184;
    wire [63:0] _3186;
    wire [63:0] _238;
    reg [63:0] _3183;
    wire [8:0] _3187;
    wire _3188;
    wire _3189;
    wire [63:0] _3193;
    wire [63:0] _3195;
    wire [63:0] _239;
    reg [63:0] _3192;
    wire [8:0] _3196;
    wire _3197;
    wire _3198;
    wire [63:0] _3202;
    wire [63:0] _3204;
    wire [63:0] _240;
    reg [63:0] _3201;
    wire [8:0] _3205;
    wire _3206;
    wire _3207;
    wire [63:0] _3211;
    wire [63:0] _3213;
    wire [63:0] _241;
    reg [63:0] _3210;
    wire [8:0] _3214;
    wire _3215;
    wire _3216;
    wire [63:0] _3220;
    wire [63:0] _3222;
    wire [63:0] _242;
    reg [63:0] _3219;
    wire [8:0] _3223;
    wire _3224;
    wire _3225;
    wire [63:0] _3229;
    wire [63:0] _3231;
    wire [63:0] _243;
    reg [63:0] _3228;
    wire [8:0] _3232;
    wire _3233;
    wire _3234;
    wire [63:0] _3238;
    wire [63:0] _3240;
    wire [63:0] _244;
    reg [63:0] _3237;
    wire [8:0] _3241;
    wire _3242;
    wire _3243;
    wire [63:0] _3247;
    wire [63:0] _3249;
    wire [63:0] _245;
    reg [63:0] _3246;
    wire [8:0] _3250;
    wire _3251;
    wire _3252;
    wire [63:0] _3256;
    wire [63:0] _3258;
    wire [63:0] _246;
    reg [63:0] _3255;
    wire [8:0] _3259;
    wire _3260;
    wire _3261;
    wire [63:0] _3265;
    wire [63:0] _3267;
    wire [63:0] _247;
    reg [63:0] _3264;
    wire [8:0] _3268;
    wire _3269;
    wire _3270;
    wire [63:0] _3274;
    wire [63:0] _3276;
    wire [63:0] _248;
    reg [63:0] _3273;
    wire [8:0] _3277;
    wire _3278;
    wire _3279;
    wire [63:0] _3283;
    wire [63:0] _3285;
    wire [63:0] _249;
    reg [63:0] _3282;
    wire [8:0] _3286;
    wire _3287;
    wire _3288;
    wire [63:0] _3292;
    wire [63:0] _3294;
    wire [63:0] _250;
    reg [63:0] _3291;
    wire [8:0] _3295;
    wire _3296;
    wire _3297;
    wire [63:0] _3301;
    wire [63:0] _3303;
    wire [63:0] _251;
    reg [63:0] _3300;
    wire [8:0] _3304;
    wire _3305;
    wire _3306;
    wire [63:0] _3310;
    wire [63:0] _3312;
    wire [63:0] _252;
    reg [63:0] _3309;
    wire [8:0] _3313;
    wire _3314;
    wire _3315;
    wire [63:0] _3319;
    wire [63:0] _3321;
    wire [63:0] _253;
    reg [63:0] _3318;
    wire [8:0] _3322;
    wire _3323;
    wire _3324;
    wire [63:0] _3328;
    wire [63:0] _3330;
    wire [63:0] _254;
    reg [63:0] _3327;
    wire [8:0] _3331;
    wire _3332;
    wire _3333;
    wire [63:0] _3337;
    wire [63:0] _3339;
    wire [63:0] _255;
    reg [63:0] _3336;
    wire [8:0] _3340;
    wire _3341;
    wire _3342;
    wire [63:0] _3346;
    wire [63:0] _3348;
    wire [63:0] _256;
    reg [63:0] _3345;
    wire [8:0] _3349;
    wire _3350;
    wire _3351;
    wire [63:0] _3355;
    wire [63:0] _3357;
    wire [63:0] _257;
    reg [63:0] _3354;
    wire [8:0] _3358;
    wire _3359;
    wire _3360;
    wire [63:0] _3364;
    wire [63:0] _3366;
    wire [63:0] _258;
    reg [63:0] _3363;
    wire [8:0] _3367;
    wire _3368;
    wire _3369;
    wire [63:0] _3373;
    wire [63:0] _3375;
    wire [63:0] _259;
    reg [63:0] _3372;
    wire [8:0] _3376;
    wire _3377;
    wire _3378;
    wire [63:0] _3382;
    wire [63:0] _3384;
    wire [63:0] _260;
    reg [63:0] _3381;
    wire [8:0] _3385;
    wire _3386;
    wire _3387;
    wire [63:0] _3391;
    wire [63:0] _3393;
    wire [63:0] _261;
    reg [63:0] _3390;
    wire [8:0] _3394;
    wire _3395;
    wire _3396;
    wire [63:0] _3400;
    wire [63:0] _3402;
    wire [63:0] _262;
    reg [63:0] _3399;
    wire [8:0] _3403;
    wire _3404;
    wire _3405;
    wire [63:0] _3409;
    wire [63:0] _3411;
    wire [63:0] _263;
    reg [63:0] _3408;
    wire [8:0] _3412;
    wire _3413;
    wire _3414;
    wire [63:0] _3418;
    wire [63:0] _3420;
    wire [63:0] _264;
    reg [63:0] _3417;
    wire [8:0] _3421;
    wire _3422;
    wire _3423;
    wire [63:0] _3427;
    wire [63:0] _3429;
    wire [63:0] _265;
    reg [63:0] _3426;
    wire [8:0] _3430;
    wire _3431;
    wire _3432;
    wire [63:0] _3436;
    wire [63:0] _3438;
    wire [63:0] _266;
    reg [63:0] _3435;
    wire [8:0] _3439;
    wire _3440;
    wire _3441;
    wire [63:0] _3445;
    wire [63:0] _3447;
    wire [63:0] _267;
    reg [63:0] _3444;
    wire [8:0] _3448;
    wire _3449;
    wire _3450;
    wire [63:0] _3454;
    wire [63:0] _3456;
    wire [63:0] _268;
    reg [63:0] _3453;
    wire [8:0] _3457;
    wire _3458;
    wire _3459;
    wire [63:0] _3463;
    wire [63:0] _3465;
    wire [63:0] _269;
    reg [63:0] _3462;
    wire [8:0] _3466;
    wire _3467;
    wire _3468;
    wire [63:0] _3472;
    wire [63:0] _3474;
    wire [63:0] _270;
    reg [63:0] _3471;
    wire [8:0] _3475;
    wire _3476;
    wire _3477;
    wire [63:0] _3481;
    wire [63:0] _3483;
    wire [63:0] _271;
    reg [63:0] _3480;
    wire [8:0] _3484;
    wire _3485;
    wire _3486;
    wire [63:0] _3490;
    wire [63:0] _3492;
    wire [63:0] _272;
    reg [63:0] _3489;
    wire [8:0] _3493;
    wire _3494;
    wire _3495;
    wire [63:0] _3499;
    wire [63:0] _3501;
    wire [63:0] _273;
    reg [63:0] _3498;
    wire [8:0] _3502;
    wire _3503;
    wire _3504;
    wire [63:0] _3508;
    wire [63:0] _3510;
    wire [63:0] _274;
    reg [63:0] _3507;
    wire [8:0] _3511;
    wire _3512;
    wire _3513;
    wire [63:0] _3517;
    wire [63:0] _3519;
    wire [63:0] _275;
    reg [63:0] _3516;
    wire [8:0] _3520;
    wire _3521;
    wire _3522;
    wire [63:0] _3526;
    wire [63:0] _3528;
    wire [63:0] _276;
    reg [63:0] _3525;
    wire [8:0] _3529;
    wire _3530;
    wire _3531;
    wire [63:0] _3535;
    wire [63:0] _3537;
    wire [63:0] _277;
    reg [63:0] _3534;
    wire [8:0] _3538;
    wire _3539;
    wire _3540;
    wire [63:0] _3544;
    wire [63:0] _3546;
    wire [63:0] _278;
    reg [63:0] _3543;
    wire [8:0] _3547;
    wire _3548;
    wire _3549;
    wire [63:0] _3553;
    wire [63:0] _3555;
    wire [63:0] _279;
    reg [63:0] _3552;
    wire [8:0] _3556;
    wire _3557;
    wire _3558;
    wire [63:0] _3562;
    wire [63:0] _3564;
    wire [63:0] _280;
    reg [63:0] _3561;
    wire [8:0] _3565;
    wire _3566;
    wire _3567;
    wire [63:0] _3571;
    wire [63:0] _3573;
    wire [63:0] _281;
    reg [63:0] _3570;
    wire [8:0] _3574;
    wire _3575;
    wire _3576;
    wire [63:0] _3580;
    wire [63:0] _3582;
    wire [63:0] _282;
    reg [63:0] _3579;
    wire [8:0] _3583;
    wire _3584;
    wire _3585;
    wire [63:0] _3589;
    wire [63:0] _3591;
    wire [63:0] _283;
    reg [63:0] _3588;
    wire [8:0] _3592;
    wire _3593;
    wire _3594;
    wire [63:0] _3598;
    wire [63:0] _3600;
    wire [63:0] _284;
    reg [63:0] _3597;
    wire [8:0] _3601;
    wire _3602;
    wire _3603;
    wire [63:0] _3607;
    wire [63:0] _3609;
    wire [63:0] _285;
    reg [63:0] _3606;
    wire [8:0] _3610;
    wire _3611;
    wire _3612;
    wire [63:0] _3616;
    wire [63:0] _3618;
    wire [63:0] _286;
    reg [63:0] _3615;
    wire [8:0] _3619;
    wire _3620;
    wire _3621;
    wire [63:0] _3625;
    wire [63:0] _3627;
    wire [63:0] _287;
    reg [63:0] _3624;
    wire [8:0] _3628;
    wire _3629;
    wire _3630;
    wire [63:0] _3634;
    wire [63:0] _3636;
    wire [63:0] _288;
    reg [63:0] _3633;
    wire [8:0] _3637;
    wire _3638;
    wire _3639;
    wire [63:0] _3643;
    wire [63:0] _3645;
    wire [63:0] _289;
    reg [63:0] _3642;
    wire [8:0] _3646;
    wire _3647;
    wire _3648;
    wire [63:0] _3652;
    wire [63:0] _3654;
    wire [63:0] _290;
    reg [63:0] _3651;
    wire [8:0] _3655;
    wire _3656;
    wire _3657;
    wire [63:0] _3661;
    wire [63:0] _3663;
    wire [63:0] _291;
    reg [63:0] _3660;
    wire [8:0] _3664;
    wire _3665;
    wire _3666;
    wire [63:0] _3670;
    wire [63:0] _3672;
    wire [63:0] _292;
    reg [63:0] _3669;
    wire [8:0] _3673;
    wire _3674;
    wire _3675;
    wire [63:0] _3679;
    wire [63:0] _3681;
    wire [63:0] _293;
    reg [63:0] _3678;
    wire [8:0] _3682;
    wire _3683;
    wire _3684;
    wire [63:0] _3688;
    wire [63:0] _3690;
    wire [63:0] _294;
    reg [63:0] _3687;
    wire [8:0] _3691;
    wire _3692;
    wire _3693;
    wire [63:0] _3697;
    wire [63:0] _3699;
    wire [63:0] _295;
    reg [63:0] _3696;
    wire [8:0] _3700;
    wire _3701;
    wire _3702;
    wire [63:0] _3706;
    wire [63:0] _3708;
    wire [63:0] _296;
    reg [63:0] _3705;
    wire [8:0] _3709;
    wire _3710;
    wire _3711;
    wire [63:0] _3715;
    wire [63:0] _3717;
    wire [63:0] _297;
    reg [63:0] _3714;
    wire [8:0] _3718;
    wire _3719;
    wire _3720;
    wire [63:0] _3724;
    wire [63:0] _3726;
    wire [63:0] _298;
    reg [63:0] _3723;
    wire [8:0] _3727;
    wire _3728;
    wire _3729;
    wire [63:0] _3733;
    wire [63:0] _3735;
    wire [63:0] _299;
    reg [63:0] _3732;
    wire [8:0] _3736;
    wire _3737;
    wire _3738;
    wire [63:0] _3742;
    wire [63:0] _3744;
    wire [63:0] _300;
    reg [63:0] _3741;
    wire [8:0] _3745;
    wire _3746;
    wire _3747;
    wire [63:0] _3751;
    wire [63:0] _3753;
    wire [63:0] _301;
    reg [63:0] _3750;
    wire [8:0] _3754;
    wire _3755;
    wire _3756;
    wire [63:0] _3760;
    wire [63:0] _3762;
    wire [63:0] _302;
    reg [63:0] _3759;
    wire [8:0] _3763;
    wire _3764;
    wire _3765;
    wire [63:0] _3769;
    wire [63:0] _3771;
    wire [63:0] _303;
    reg [63:0] _3768;
    wire [8:0] _3772;
    wire _3773;
    wire _3774;
    wire [63:0] _3778;
    wire [63:0] _3780;
    wire [63:0] _304;
    reg [63:0] _3777;
    wire [8:0] _3781;
    wire _3782;
    wire _3783;
    wire [63:0] _3787;
    wire [63:0] _3789;
    wire [63:0] _305;
    reg [63:0] _3786;
    wire [8:0] _3790;
    wire _3791;
    wire _3792;
    wire [63:0] _3796;
    wire [63:0] _3798;
    wire [63:0] _306;
    reg [63:0] _3795;
    wire [8:0] _3799;
    wire _3800;
    wire _3801;
    wire [63:0] _3805;
    wire [63:0] _3807;
    wire [63:0] _307;
    reg [63:0] _3804;
    wire [8:0] _3808;
    wire _3809;
    wire _3810;
    wire [63:0] _3814;
    wire [63:0] _3816;
    wire [63:0] _308;
    reg [63:0] _3813;
    wire [8:0] _3817;
    wire _3818;
    wire _3819;
    wire [63:0] _3823;
    wire [63:0] _3825;
    wire [63:0] _309;
    reg [63:0] _3822;
    wire [8:0] _3826;
    wire _3827;
    wire _3828;
    wire [63:0] _3832;
    wire [63:0] _3834;
    wire [63:0] _310;
    reg [63:0] _3831;
    wire [8:0] _3835;
    wire _3836;
    wire _3837;
    wire [63:0] _3841;
    wire [63:0] _3843;
    wire [63:0] _311;
    reg [63:0] _3840;
    wire [8:0] _3844;
    wire _3845;
    wire _3846;
    wire [63:0] _3850;
    wire [63:0] _3852;
    wire [63:0] _312;
    reg [63:0] _3849;
    wire [8:0] _3853;
    wire _3854;
    wire _3855;
    wire [63:0] _3859;
    wire [63:0] _3861;
    wire [63:0] _313;
    reg [63:0] _3858;
    wire [8:0] _3862;
    wire _3863;
    wire _3864;
    wire [63:0] _3868;
    wire [63:0] _3870;
    wire [63:0] _314;
    reg [63:0] _3867;
    wire [8:0] _3871;
    wire _3872;
    wire _3873;
    wire [63:0] _3877;
    wire [63:0] _3879;
    wire [63:0] _315;
    reg [63:0] _3876;
    wire [8:0] _3880;
    wire _3881;
    wire _3882;
    wire [63:0] _3886;
    wire [63:0] _3888;
    wire [63:0] _316;
    reg [63:0] _3885;
    wire [8:0] _3889;
    wire _3890;
    wire _3891;
    wire [63:0] _3895;
    wire [63:0] _3897;
    wire [63:0] _317;
    reg [63:0] _3894;
    wire [8:0] _3898;
    wire _3899;
    wire _3900;
    wire [63:0] _3904;
    wire [63:0] _3906;
    wire [63:0] _318;
    reg [63:0] _3903;
    wire [8:0] _3907;
    wire _3908;
    wire _3909;
    wire [63:0] _3913;
    wire [63:0] _3915;
    wire [63:0] _319;
    reg [63:0] _3912;
    wire [8:0] _3916;
    wire _3917;
    wire _3918;
    wire [63:0] _3922;
    wire [63:0] _3924;
    wire [63:0] _320;
    reg [63:0] _3921;
    wire [8:0] _3925;
    wire _3926;
    wire _3927;
    wire [63:0] _3931;
    wire [63:0] _3933;
    wire [63:0] _321;
    reg [63:0] _3930;
    wire [8:0] _3934;
    wire _3935;
    wire _3936;
    wire [63:0] _3940;
    wire [63:0] _3942;
    wire [63:0] _322;
    reg [63:0] _3939;
    wire [8:0] _3943;
    wire _3944;
    wire _3945;
    wire [63:0] _3949;
    wire [63:0] _3951;
    wire [63:0] _323;
    reg [63:0] _3948;
    wire [8:0] _3952;
    wire _3953;
    wire _3954;
    wire [63:0] _3958;
    wire [63:0] _3960;
    wire [63:0] _324;
    reg [63:0] _3957;
    wire [8:0] _3961;
    wire _3962;
    wire _3963;
    wire [63:0] _3967;
    wire [63:0] _3969;
    wire [63:0] _325;
    reg [63:0] _3966;
    wire [8:0] _3970;
    wire _3971;
    wire _3972;
    wire [63:0] _3976;
    wire [63:0] _3978;
    wire [63:0] _326;
    reg [63:0] _3975;
    wire [8:0] _3979;
    wire _3980;
    wire _3981;
    wire [63:0] _3985;
    wire [63:0] _3987;
    wire [63:0] _327;
    reg [63:0] _3984;
    wire [8:0] _3988;
    wire _3989;
    wire _3990;
    wire [63:0] _3994;
    wire [63:0] _3996;
    wire [63:0] _328;
    reg [63:0] _3993;
    wire [8:0] _3997;
    wire _3998;
    wire _3999;
    wire [63:0] _4003;
    wire [63:0] _4005;
    wire [63:0] _329;
    reg [63:0] _4002;
    wire [8:0] _4006;
    wire _4007;
    wire _4008;
    wire [63:0] _4012;
    wire [63:0] _4014;
    wire [63:0] _330;
    reg [63:0] _4011;
    wire [8:0] _4015;
    wire _4016;
    wire _4017;
    wire [63:0] _4021;
    wire [63:0] _4023;
    wire [63:0] _331;
    reg [63:0] _4020;
    wire [8:0] _4024;
    wire _4025;
    wire _4026;
    wire [63:0] _4030;
    wire [63:0] _4032;
    wire [63:0] _332;
    reg [63:0] _4029;
    wire [8:0] _4033;
    wire _4034;
    wire _4035;
    wire [63:0] _4039;
    wire [63:0] _4041;
    wire [63:0] _333;
    reg [63:0] _4038;
    wire [8:0] _4042;
    wire _4043;
    wire _4044;
    wire [63:0] _4048;
    wire [63:0] _4050;
    wire [63:0] _334;
    reg [63:0] _4047;
    wire [8:0] _4051;
    wire _4052;
    wire _4053;
    wire [63:0] _4057;
    wire [63:0] _4059;
    wire [63:0] _335;
    reg [63:0] _4056;
    wire [8:0] _4060;
    wire _4061;
    wire _4062;
    wire [63:0] _4066;
    wire [63:0] _4068;
    wire [63:0] _336;
    reg [63:0] _4065;
    wire [8:0] _4069;
    wire _4070;
    wire _4071;
    wire [63:0] _4075;
    wire [63:0] _4077;
    wire [63:0] _337;
    reg [63:0] _4074;
    wire [8:0] _4078;
    wire _4079;
    wire _4080;
    wire [63:0] _4084;
    wire [63:0] _4086;
    wire [63:0] _338;
    reg [63:0] _4083;
    wire [8:0] _4087;
    wire _4088;
    wire _4089;
    wire [63:0] _4093;
    wire [63:0] _4095;
    wire [63:0] _339;
    reg [63:0] _4092;
    wire [8:0] _4096;
    wire _4097;
    wire _4098;
    wire [63:0] _4102;
    wire [63:0] _4104;
    wire [63:0] _340;
    reg [63:0] _4101;
    wire [8:0] _4105;
    wire _4106;
    wire _4107;
    wire [63:0] _4111;
    wire [63:0] _4113;
    wire [63:0] _341;
    reg [63:0] _4110;
    wire [8:0] _4114;
    wire _4115;
    wire _4116;
    wire [63:0] _4120;
    wire [63:0] _4122;
    wire [63:0] _342;
    reg [63:0] _4119;
    wire [8:0] _4123;
    wire _4124;
    wire _4125;
    wire [63:0] _4129;
    wire [63:0] _4131;
    wire [63:0] _343;
    reg [63:0] _4128;
    wire [8:0] _4132;
    wire _4133;
    wire _4134;
    wire [63:0] _4138;
    wire [63:0] _4140;
    wire [63:0] _344;
    reg [63:0] _4137;
    wire [8:0] _4141;
    wire _4142;
    wire _4143;
    wire [63:0] _4147;
    wire [63:0] _4149;
    wire [63:0] _345;
    reg [63:0] _4146;
    wire [8:0] _4150;
    wire _4151;
    wire _4152;
    wire [63:0] _4156;
    wire [63:0] _4158;
    wire [63:0] _346;
    reg [63:0] _4155;
    wire [8:0] _4159;
    wire _4160;
    wire _4161;
    wire [63:0] _4165;
    wire [63:0] _4167;
    wire [63:0] _347;
    reg [63:0] _4164;
    wire [8:0] _4168;
    wire _4169;
    wire _4170;
    wire [63:0] _4174;
    wire [63:0] _4176;
    wire [63:0] _348;
    reg [63:0] _4173;
    wire [8:0] _4177;
    wire _4178;
    wire _4179;
    wire [63:0] _4183;
    wire [63:0] _4185;
    wire [63:0] _349;
    reg [63:0] _4182;
    wire [8:0] _4186;
    wire _4187;
    wire _4188;
    wire [63:0] _4192;
    wire [63:0] _4194;
    wire [63:0] _350;
    reg [63:0] _4191;
    wire [8:0] _4195;
    wire _4196;
    wire _4197;
    wire [63:0] _4201;
    wire [63:0] _4203;
    wire [63:0] _351;
    reg [63:0] _4200;
    wire [8:0] _4204;
    wire _4205;
    wire _4206;
    wire [63:0] _4210;
    wire [63:0] _4212;
    wire [63:0] _352;
    reg [63:0] _4209;
    wire [8:0] _4213;
    wire _4214;
    wire _4215;
    wire [63:0] _4219;
    wire [63:0] _4221;
    wire [63:0] _353;
    reg [63:0] _4218;
    wire [8:0] _4222;
    wire _4223;
    wire _4224;
    wire [63:0] _4228;
    wire [63:0] _4230;
    wire [63:0] _354;
    reg [63:0] _4227;
    wire [8:0] _4231;
    wire _4232;
    wire _4233;
    wire [63:0] _4237;
    wire [63:0] _4239;
    wire [63:0] _355;
    reg [63:0] _4236;
    wire [8:0] _4240;
    wire _4241;
    wire _4242;
    wire [63:0] _4246;
    wire [63:0] _4248;
    wire [63:0] _356;
    reg [63:0] _4245;
    wire [8:0] _4249;
    wire _4250;
    wire _4251;
    wire [63:0] _4255;
    wire [63:0] _4257;
    wire [63:0] _357;
    reg [63:0] _4254;
    wire [8:0] _4258;
    wire _4259;
    wire _4260;
    wire [63:0] _4264;
    wire [63:0] _4266;
    wire [63:0] _358;
    reg [63:0] _4263;
    wire [8:0] _4267;
    wire _4268;
    wire _4269;
    wire [63:0] _4273;
    wire [63:0] _4275;
    wire [63:0] _359;
    reg [63:0] _4272;
    wire [8:0] _4276;
    wire _4277;
    wire _4278;
    wire [63:0] _4282;
    wire [63:0] _4284;
    wire [63:0] _360;
    reg [63:0] _4281;
    wire [8:0] _4285;
    wire _4286;
    wire _4287;
    wire [63:0] _4291;
    wire [63:0] _4293;
    wire [63:0] _361;
    reg [63:0] _4290;
    wire [8:0] _4294;
    wire _4295;
    wire _4296;
    wire [63:0] _4300;
    wire [63:0] _4302;
    wire [63:0] _362;
    reg [63:0] _4299;
    wire [8:0] _4303;
    wire _4304;
    wire _4305;
    wire [63:0] _4309;
    wire [63:0] _4311;
    wire [63:0] _363;
    reg [63:0] _4308;
    wire [8:0] _4312;
    wire _4313;
    wire _4314;
    wire [63:0] _4318;
    wire [63:0] _4320;
    wire [63:0] _364;
    reg [63:0] _4317;
    wire [8:0] _4321;
    wire _4322;
    wire _4323;
    wire [63:0] _4327;
    wire [63:0] _4329;
    wire [63:0] _365;
    reg [63:0] _4326;
    wire [8:0] _4330;
    wire _4331;
    wire _4332;
    wire [63:0] _4336;
    wire [63:0] _4338;
    wire [63:0] _366;
    reg [63:0] _4335;
    wire [8:0] _4339;
    wire _4340;
    wire _4341;
    wire [63:0] _4345;
    wire [63:0] _4347;
    wire [63:0] _367;
    reg [63:0] _4344;
    wire [8:0] _4348;
    wire _4349;
    wire _4350;
    wire [63:0] _4354;
    wire [63:0] _4356;
    wire [63:0] _368;
    reg [63:0] _4353;
    wire [8:0] _4357;
    wire _4358;
    wire _4359;
    wire [63:0] _4363;
    wire [63:0] _4365;
    wire [63:0] _369;
    reg [63:0] _4362;
    wire [8:0] _4366;
    wire _4367;
    wire _4368;
    wire [63:0] _4372;
    wire [63:0] _4374;
    wire [63:0] _370;
    reg [63:0] _4371;
    wire [8:0] _4375;
    wire _4376;
    wire _4377;
    wire [63:0] _4381;
    wire [63:0] _4383;
    wire [63:0] _371;
    reg [63:0] _4380;
    wire [8:0] _4384;
    wire _4385;
    wire _4386;
    wire [63:0] _4390;
    wire [63:0] _4392;
    wire [63:0] _372;
    reg [63:0] _4389;
    wire [8:0] _4393;
    wire _4394;
    wire _4395;
    wire [63:0] _4399;
    wire [63:0] _4401;
    wire [63:0] _373;
    reg [63:0] _4398;
    wire [8:0] _4402;
    wire _4403;
    wire _4404;
    wire [63:0] _4408;
    wire [63:0] _4410;
    wire [63:0] _374;
    reg [63:0] _4407;
    wire [8:0] _4411;
    wire _4412;
    wire _4413;
    wire [63:0] _4417;
    wire [63:0] _4419;
    wire [63:0] _375;
    reg [63:0] _4416;
    wire [8:0] _4420;
    wire _4421;
    wire _4422;
    wire [63:0] _4426;
    wire [63:0] _4428;
    wire [63:0] _376;
    reg [63:0] _4425;
    wire [8:0] _4429;
    wire _4430;
    wire _4431;
    wire [63:0] _4435;
    wire [63:0] _4437;
    wire [63:0] _377;
    reg [63:0] _4434;
    wire [8:0] _4438;
    wire _4439;
    wire _4440;
    wire [63:0] _4444;
    wire [63:0] _4446;
    wire [63:0] _378;
    reg [63:0] _4443;
    wire [8:0] _4447;
    wire _4448;
    wire _4449;
    wire [63:0] _4453;
    wire [63:0] _4455;
    wire [63:0] _379;
    reg [63:0] _4452;
    wire [8:0] _4456;
    wire _4457;
    wire _4458;
    wire [63:0] _4462;
    wire [63:0] _4464;
    wire [63:0] _380;
    reg [63:0] _4461;
    wire [8:0] _4465;
    wire _4466;
    wire _4467;
    wire [63:0] _4471;
    wire [63:0] _4473;
    wire [63:0] _381;
    reg [63:0] _4470;
    wire [8:0] _4474;
    wire _4475;
    wire _4476;
    wire [63:0] _4480;
    wire [63:0] _4482;
    wire [63:0] _382;
    reg [63:0] _4479;
    wire [8:0] _4483;
    wire _4484;
    wire _4485;
    wire [63:0] _4489;
    wire [63:0] _4491;
    wire [63:0] _383;
    reg [63:0] _4488;
    wire [8:0] _4492;
    wire _4493;
    wire _4494;
    wire [63:0] _4498;
    wire [63:0] _4500;
    wire [63:0] _384;
    reg [63:0] _4497;
    wire [8:0] _4501;
    wire _4502;
    wire _4503;
    wire [63:0] _4507;
    wire [63:0] _4509;
    wire [63:0] _385;
    reg [63:0] _4506;
    wire [8:0] _4510;
    wire _4511;
    wire _4512;
    wire [63:0] _4516;
    wire [63:0] _4518;
    wire [63:0] _386;
    reg [63:0] _4515;
    wire [8:0] _4519;
    wire _4520;
    wire _4521;
    wire [63:0] _4525;
    wire [63:0] _4527;
    wire [63:0] _387;
    reg [63:0] _4524;
    wire [8:0] _4528;
    wire _4529;
    wire _4530;
    wire [63:0] _4534;
    wire [63:0] _4536;
    wire [63:0] _388;
    reg [63:0] _4533;
    wire [8:0] _4537;
    wire _4538;
    wire _4539;
    wire [63:0] _4543;
    wire [63:0] _4545;
    wire [63:0] _389;
    reg [63:0] _4542;
    wire [8:0] _4546;
    wire _4547;
    wire _4548;
    wire [63:0] _4552;
    wire [63:0] _4554;
    wire [63:0] _390;
    reg [63:0] _4551;
    wire [8:0] _4555;
    wire _4556;
    wire _4557;
    wire [63:0] _4561;
    wire [63:0] _4563;
    wire [63:0] _391;
    reg [63:0] _4560;
    wire [8:0] _4564;
    wire _4565;
    wire _4566;
    wire [63:0] _4570;
    wire [63:0] _4572;
    wire [63:0] _392;
    reg [63:0] _4569;
    wire [8:0] _4573;
    wire _4574;
    wire _4575;
    wire [63:0] _4579;
    wire [63:0] _4581;
    wire [63:0] _393;
    reg [63:0] _4578;
    wire [8:0] _4582;
    wire _4583;
    wire _4584;
    wire [63:0] _4588;
    wire [63:0] _4590;
    wire [63:0] _394;
    reg [63:0] _4587;
    wire [8:0] _4591;
    wire _4592;
    wire _4593;
    wire [63:0] _4597;
    wire [63:0] _4599;
    wire [63:0] _395;
    reg [63:0] _4596;
    wire [8:0] _4600;
    wire _4601;
    wire _4602;
    wire [63:0] _4606;
    wire [63:0] _4608;
    wire [63:0] _396;
    reg [63:0] _4605;
    wire [8:0] _4609;
    wire _4610;
    wire _4611;
    wire [63:0] _4615;
    wire [63:0] _4617;
    wire [63:0] _397;
    reg [63:0] _4614;
    wire [8:0] _4618;
    wire _4619;
    wire _4620;
    wire [63:0] _4624;
    wire [63:0] _4626;
    wire [63:0] _398;
    reg [63:0] _4623;
    wire [8:0] _4627;
    wire _4628;
    wire _4629;
    wire [63:0] _4633;
    wire [63:0] _4635;
    wire [63:0] _399;
    reg [63:0] _4632;
    wire [8:0] _4636;
    wire _4637;
    wire _4638;
    wire [63:0] _4642;
    wire [63:0] _4644;
    wire [63:0] _400;
    reg [63:0] _4641;
    wire [8:0] _4645;
    wire _4646;
    wire _4647;
    wire [63:0] _4651;
    wire [63:0] _4653;
    wire [63:0] _401;
    reg [63:0] _4650;
    wire [8:0] _4654;
    wire _4655;
    wire _4656;
    wire [63:0] _4660;
    wire [63:0] _4662;
    wire [63:0] _402;
    reg [63:0] _4659;
    wire [8:0] _4663;
    wire _4664;
    wire _4665;
    wire [63:0] _4669;
    wire [63:0] _4671;
    wire [63:0] _403;
    reg [63:0] _4668;
    wire [8:0] _4672;
    wire _4673;
    wire _4674;
    wire [63:0] _4678;
    wire [63:0] _4680;
    wire [63:0] _404;
    reg [63:0] _4677;
    wire [8:0] _4681;
    wire _4682;
    wire _4683;
    wire [63:0] _4687;
    wire [63:0] _4689;
    wire [63:0] _405;
    reg [63:0] _4686;
    wire [8:0] _4690;
    wire _4691;
    wire _4692;
    wire [63:0] _4696;
    wire [63:0] _4698;
    wire [63:0] _406;
    reg [63:0] _4695;
    wire [8:0] _4699;
    wire _4700;
    wire _4701;
    wire [63:0] _4705;
    wire [63:0] _4707;
    wire [63:0] _407;
    reg [63:0] _4704;
    wire [8:0] _4708;
    wire _4709;
    wire _4710;
    wire [63:0] _4714;
    wire [63:0] _4716;
    wire [63:0] _408;
    reg [63:0] _4713;
    wire [8:0] _4717;
    wire _4718;
    wire _4719;
    wire [63:0] _4723;
    wire [63:0] _4725;
    wire [63:0] _409;
    reg [63:0] _4722;
    wire [8:0] _4726;
    wire _4727;
    wire _4728;
    wire [63:0] _4732;
    wire [63:0] _4734;
    wire [63:0] _410;
    reg [63:0] _4731;
    wire [8:0] _4735;
    wire _4736;
    wire _4737;
    wire [63:0] _4741;
    wire [63:0] _4743;
    wire [63:0] _411;
    reg [63:0] _4740;
    wire [8:0] _4744;
    wire _4745;
    wire _4746;
    wire [63:0] _4750;
    wire [63:0] _4752;
    wire [63:0] _412;
    reg [63:0] _4749;
    wire [8:0] _4753;
    wire _4754;
    wire _4755;
    wire [63:0] _4759;
    wire [63:0] _4761;
    wire [63:0] _413;
    reg [63:0] _4758;
    wire [8:0] _4762;
    wire _4763;
    wire _4764;
    wire [63:0] _4768;
    wire [63:0] _4770;
    wire [63:0] _414;
    reg [63:0] _4767;
    wire [8:0] _4771;
    wire _4772;
    wire _4773;
    wire [63:0] _4777;
    wire [63:0] _4779;
    wire [63:0] _415;
    reg [63:0] _4776;
    wire [8:0] _4780;
    wire _4781;
    wire _4782;
    wire [63:0] _4786;
    wire [63:0] _4788;
    wire [63:0] _416;
    reg [63:0] _4785;
    wire [8:0] _4789;
    wire _4790;
    wire _4791;
    wire [63:0] _4795;
    wire [63:0] _4797;
    wire [63:0] _417;
    reg [63:0] _4794;
    wire [8:0] _4798;
    wire _4799;
    wire _4800;
    wire [63:0] _4804;
    wire [63:0] _4806;
    wire [63:0] _418;
    reg [63:0] _4803;
    wire [8:0] _4807;
    wire _4808;
    wire _4809;
    wire [63:0] _4813;
    wire [63:0] _4815;
    wire [63:0] _419;
    reg [63:0] _4812;
    wire [8:0] _4816;
    wire _4817;
    wire _4818;
    wire [63:0] _4822;
    wire [63:0] _4824;
    wire [63:0] _420;
    reg [63:0] _4821;
    wire [8:0] _4825;
    wire _4826;
    wire _4827;
    wire [63:0] _4831;
    wire [63:0] _4833;
    wire [63:0] _421;
    reg [63:0] _4830;
    wire [8:0] _4834;
    wire _4835;
    wire _4836;
    wire [63:0] _4840;
    wire [63:0] _4842;
    wire [63:0] _422;
    reg [63:0] _4839;
    wire [8:0] _4843;
    wire _4844;
    wire _4845;
    wire [63:0] _4849;
    wire [63:0] _4851;
    wire [63:0] _423;
    reg [63:0] _4848;
    wire [8:0] _4852;
    wire _4853;
    wire _4854;
    wire [63:0] _4858;
    wire [63:0] _4860;
    wire [63:0] _424;
    reg [63:0] _4857;
    wire [8:0] _4861;
    wire _4862;
    wire _4863;
    wire [63:0] _4867;
    wire [63:0] _4869;
    wire [63:0] _425;
    reg [63:0] _4866;
    wire [8:0] _4870;
    wire _4871;
    wire _4872;
    wire [63:0] _4876;
    wire [63:0] _4878;
    wire [63:0] _426;
    reg [63:0] _4875;
    wire [8:0] _4879;
    wire _4880;
    wire _4881;
    wire [63:0] _4885;
    wire [63:0] _4887;
    wire [63:0] _427;
    reg [63:0] _4884;
    wire [8:0] _4888;
    wire _4889;
    wire _4890;
    wire [63:0] _4894;
    wire [63:0] _4896;
    wire [63:0] _428;
    reg [63:0] _4893;
    wire [8:0] _4897;
    wire _4898;
    wire _4899;
    wire [63:0] _4903;
    wire [63:0] _4905;
    wire [63:0] _429;
    reg [63:0] _4902;
    wire [8:0] _4906;
    wire _4907;
    wire _4908;
    wire [63:0] _4912;
    wire [63:0] _4914;
    wire [63:0] _430;
    reg [63:0] _4911;
    wire [8:0] _4915;
    wire _4916;
    wire _4917;
    wire [63:0] _4921;
    wire [63:0] _4923;
    wire [63:0] _431;
    reg [63:0] _4920;
    wire [8:0] _4924;
    wire _4925;
    wire _4926;
    wire [63:0] _4930;
    wire [63:0] _4932;
    wire [63:0] _432;
    reg [63:0] _4929;
    wire [8:0] _4933;
    wire _4934;
    wire _4935;
    wire [63:0] _4939;
    wire [63:0] _4941;
    wire [63:0] _433;
    reg [63:0] _4938;
    wire [8:0] _4942;
    wire _4943;
    wire _4944;
    wire [63:0] _4948;
    wire [63:0] _4950;
    wire [63:0] _434;
    reg [63:0] _4947;
    wire [8:0] _4951;
    wire _4952;
    wire _4953;
    wire [63:0] _4957;
    wire [63:0] _4959;
    wire [63:0] _435;
    reg [63:0] _4956;
    wire [8:0] _4960;
    wire _4961;
    wire _4962;
    wire [63:0] _4966;
    wire [63:0] _4968;
    wire [63:0] _436;
    reg [63:0] _4965;
    wire [8:0] _4969;
    wire _4970;
    wire _4971;
    wire [63:0] _4975;
    wire [63:0] _4977;
    wire [63:0] _437;
    reg [63:0] _4974;
    wire [8:0] _4978;
    wire _4979;
    wire _4980;
    wire [63:0] _4984;
    wire [63:0] _4986;
    wire [63:0] _438;
    reg [63:0] _4983;
    wire [8:0] _4987;
    wire _4988;
    wire _4989;
    wire [63:0] _4993;
    wire [63:0] _4995;
    wire [63:0] _439;
    reg [63:0] _4992;
    wire [8:0] _4996;
    wire _4997;
    wire _4998;
    wire [63:0] _5002;
    wire [63:0] _5004;
    wire [63:0] _440;
    reg [63:0] _5001;
    wire [8:0] _5005;
    wire _5006;
    wire _5007;
    wire [63:0] _5011;
    wire [63:0] _5013;
    wire [63:0] _441;
    reg [63:0] _5010;
    wire [8:0] _5014;
    wire _5015;
    wire _5016;
    wire [63:0] _5020;
    wire [63:0] _5022;
    wire [63:0] _442;
    reg [63:0] _5019;
    wire [8:0] _5023;
    wire _5024;
    wire _5025;
    wire [63:0] _5029;
    wire [63:0] _5031;
    wire [63:0] _443;
    reg [63:0] _5028;
    wire [8:0] _5032;
    wire _5033;
    wire _5034;
    wire [63:0] _5038;
    wire [63:0] _5040;
    wire [63:0] _444;
    reg [63:0] _5037;
    wire [8:0] _5041;
    wire _5042;
    wire _5043;
    wire [63:0] _5047;
    wire [63:0] _5049;
    wire [63:0] _445;
    reg [63:0] _5046;
    wire [8:0] _5050;
    wire _5051;
    wire _5052;
    wire [63:0] _5056;
    wire [63:0] _5058;
    wire [63:0] _446;
    reg [63:0] _5055;
    wire [8:0] _5059;
    wire _5060;
    wire _5061;
    wire [63:0] _5065;
    wire [63:0] _5067;
    wire [63:0] _447;
    reg [63:0] _5064;
    wire [8:0] _5068;
    wire _5069;
    wire _5070;
    wire [63:0] _5074;
    wire [63:0] _5076;
    wire [63:0] _448;
    reg [63:0] _5073;
    wire [8:0] _5077;
    wire _5078;
    wire _5079;
    wire [63:0] _5083;
    wire [63:0] _5085;
    wire [63:0] _449;
    reg [63:0] _5082;
    wire [8:0] _5086;
    wire _5087;
    wire _5088;
    wire [63:0] _5092;
    wire [63:0] _5094;
    wire [63:0] _450;
    reg [63:0] _5091;
    wire [8:0] _5095;
    wire _5096;
    wire _5097;
    wire [63:0] _5101;
    wire [63:0] _5103;
    wire [63:0] _451;
    reg [63:0] _5100;
    wire [8:0] _5104;
    wire _5105;
    wire _5106;
    wire [63:0] _5110;
    wire [63:0] _5112;
    wire [63:0] _452;
    reg [63:0] _5109;
    wire [8:0] _5113;
    wire _5114;
    wire _5115;
    wire [63:0] _5119;
    wire [63:0] _5121;
    wire [63:0] _453;
    reg [63:0] _5118;
    wire [8:0] _5122;
    wire _5123;
    wire _5124;
    wire [63:0] _5128;
    wire [63:0] _5130;
    wire [63:0] _454;
    reg [63:0] _5127;
    wire [8:0] _5131;
    wire _5132;
    wire _5133;
    wire [63:0] _5137;
    wire [63:0] _5139;
    wire [63:0] _455;
    reg [63:0] _5136;
    wire [8:0] _5140;
    wire _5141;
    wire _5142;
    wire [63:0] _5146;
    wire [63:0] _5148;
    wire [63:0] _456;
    reg [63:0] _5145;
    wire [8:0] _5149;
    wire _5150;
    wire _5151;
    wire [63:0] _5155;
    wire [63:0] _5157;
    wire [63:0] _457;
    reg [63:0] _5154;
    wire [8:0] _5158;
    wire _5159;
    wire _5160;
    wire [63:0] _5164;
    wire [63:0] _5166;
    wire [63:0] _458;
    reg [63:0] _5163;
    wire [8:0] _5167;
    wire _5168;
    wire _5169;
    wire [63:0] _5173;
    wire [63:0] _5175;
    wire [63:0] _459;
    reg [63:0] _5172;
    wire [8:0] _5176;
    wire _5177;
    wire _5178;
    wire [63:0] _5182;
    wire [63:0] _5184;
    wire [63:0] _460;
    reg [63:0] _5181;
    wire [8:0] _5185;
    wire _5186;
    wire _5187;
    wire [63:0] _5191;
    wire [63:0] _5193;
    wire [63:0] _461;
    reg [63:0] _5190;
    wire [8:0] _5194;
    wire _5195;
    wire _5196;
    wire [63:0] _5200;
    wire [63:0] _5202;
    wire [63:0] _462;
    reg [63:0] _5199;
    wire [8:0] _5203;
    wire _5204;
    wire _5205;
    wire [63:0] _5209;
    wire [63:0] _5211;
    wire [63:0] _463;
    reg [63:0] _5208;
    wire [8:0] _5212;
    wire _5213;
    wire _5214;
    wire [63:0] _5218;
    wire [63:0] _5220;
    wire [63:0] _464;
    reg [63:0] _5217;
    wire [8:0] _5221;
    wire _5222;
    wire _5223;
    wire [63:0] _5227;
    wire [63:0] _5229;
    wire [63:0] _465;
    reg [63:0] _5226;
    wire [8:0] _5230;
    wire _5231;
    wire _5232;
    wire [63:0] _5236;
    wire [63:0] _5238;
    wire [63:0] _466;
    reg [63:0] _5235;
    wire [8:0] _5239;
    wire _5240;
    wire _5241;
    wire [63:0] _5245;
    wire [63:0] _5247;
    wire [63:0] _467;
    reg [63:0] _5244;
    wire [8:0] _5248;
    wire _5249;
    wire _5250;
    wire [63:0] _5254;
    wire [63:0] _5256;
    wire [63:0] _468;
    reg [63:0] _5253;
    wire [8:0] _5257;
    wire _5258;
    wire _5259;
    wire [63:0] _5263;
    wire [63:0] _5265;
    wire [63:0] _469;
    reg [63:0] _5262;
    wire [8:0] _5266;
    wire _5267;
    wire _5268;
    wire [63:0] _5272;
    wire [63:0] _5274;
    wire [63:0] _470;
    reg [63:0] _5271;
    wire [8:0] _5275;
    wire _5276;
    wire _5277;
    wire [63:0] _5281;
    wire [63:0] _5283;
    wire [63:0] _471;
    reg [63:0] _5280;
    wire [8:0] _5284;
    wire _5285;
    wire _5286;
    wire [63:0] _5290;
    wire [63:0] _5292;
    wire [63:0] _472;
    reg [63:0] _5289;
    wire [8:0] _5293;
    wire _5294;
    wire _5295;
    wire [63:0] _5299;
    wire [63:0] _5301;
    wire [63:0] _473;
    reg [63:0] _5298;
    wire [8:0] _5302;
    wire _5303;
    wire _5304;
    wire [63:0] _5308;
    wire [63:0] _5310;
    wire [63:0] _474;
    reg [63:0] _5307;
    wire [8:0] _5311;
    wire _5312;
    wire _5313;
    wire [63:0] _5317;
    wire [63:0] _5319;
    wire [63:0] _475;
    reg [63:0] _5316;
    wire [8:0] _5320;
    wire _5321;
    wire _5322;
    wire [63:0] _5326;
    wire [63:0] _5328;
    wire [63:0] _476;
    reg [63:0] _5325;
    wire [8:0] _5329;
    wire _5330;
    wire _5331;
    wire [63:0] _5335;
    wire [63:0] _5337;
    wire [63:0] _477;
    reg [63:0] _5334;
    wire [8:0] _5338;
    wire _5339;
    wire _5340;
    wire [63:0] _5344;
    wire [63:0] _5346;
    wire [63:0] _478;
    reg [63:0] _5343;
    wire [8:0] _5347;
    wire _5348;
    wire _5349;
    wire [63:0] _5353;
    wire [63:0] _5355;
    wire [63:0] _479;
    reg [63:0] _5352;
    wire [8:0] _5356;
    wire _5357;
    wire _5358;
    wire [63:0] _5362;
    wire [63:0] _5364;
    wire [63:0] _480;
    reg [63:0] _5361;
    wire [8:0] _5365;
    wire _5366;
    wire _5367;
    wire [63:0] _5371;
    wire [63:0] _5373;
    wire [63:0] _481;
    reg [63:0] _5370;
    wire [8:0] _5374;
    wire _5375;
    wire _5376;
    wire [63:0] _5380;
    wire [63:0] _5382;
    wire [63:0] _482;
    reg [63:0] _5379;
    wire [8:0] _5383;
    wire _5384;
    wire _5385;
    wire [63:0] _5389;
    wire [63:0] _5391;
    wire [63:0] _483;
    reg [63:0] _5388;
    wire [8:0] _5392;
    wire _5393;
    wire _5394;
    wire [63:0] _5398;
    wire [63:0] _5400;
    wire [63:0] _484;
    reg [63:0] _5397;
    wire [8:0] _5401;
    wire _5402;
    wire _5403;
    wire [63:0] _5407;
    wire [63:0] _5409;
    wire [63:0] _485;
    reg [63:0] _5406;
    wire [8:0] _5410;
    wire _5411;
    wire _5412;
    wire [63:0] _5416;
    wire [63:0] _5418;
    wire [63:0] _486;
    reg [63:0] _5415;
    wire [8:0] _5419;
    wire _5420;
    wire _5421;
    wire [63:0] _5425;
    wire [63:0] _5427;
    wire [63:0] _487;
    reg [63:0] _5424;
    wire [8:0] _5428;
    wire _5429;
    wire _5430;
    wire [63:0] _5434;
    wire [63:0] _5436;
    wire [63:0] _488;
    reg [63:0] _5433;
    wire [8:0] _5437;
    wire _5438;
    wire _5439;
    wire [63:0] _5443;
    wire [63:0] _5445;
    wire [63:0] _489;
    reg [63:0] _5442;
    wire [8:0] _5446;
    wire _5447;
    wire _5448;
    wire [63:0] _5452;
    wire [63:0] _5454;
    wire [63:0] _490;
    reg [63:0] _5451;
    wire [8:0] _5455;
    wire _5456;
    wire _5457;
    wire [63:0] _5461;
    wire [63:0] _5463;
    wire [63:0] _491;
    reg [63:0] _5460;
    wire [8:0] _5464;
    wire _5465;
    wire _5466;
    wire [63:0] _5470;
    wire [63:0] _5472;
    wire [63:0] _492;
    reg [63:0] _5469;
    wire [8:0] _5473;
    wire _5474;
    wire _5475;
    wire [63:0] _5479;
    wire [63:0] _5481;
    wire [63:0] _493;
    reg [63:0] _5478;
    wire [8:0] _5482;
    wire _5483;
    wire _5484;
    wire [63:0] _5488;
    wire [63:0] _5490;
    wire [63:0] _494;
    reg [63:0] _5487;
    wire [8:0] _5491;
    wire _5492;
    wire _5493;
    wire [63:0] _5497;
    wire [63:0] _5499;
    wire [63:0] _495;
    reg [63:0] _5496;
    wire [8:0] _5500;
    wire _5501;
    wire _5502;
    wire [63:0] _5506;
    wire [63:0] _5508;
    wire [63:0] _496;
    reg [63:0] _5505;
    wire [8:0] _5509;
    wire _5510;
    wire _5511;
    wire [63:0] _5515;
    wire [63:0] _5517;
    wire [63:0] _497;
    reg [63:0] _5514;
    wire [8:0] _5518;
    wire _5519;
    wire _5520;
    wire [63:0] _5524;
    wire [63:0] _5526;
    wire [63:0] _498;
    reg [63:0] _5523;
    wire [8:0] _5527;
    wire _5528;
    wire _5529;
    wire [63:0] _5533;
    wire [63:0] _5535;
    wire [63:0] _499;
    reg [63:0] _5532;
    wire [8:0] _5536;
    wire _5537;
    wire _5538;
    wire [63:0] _5542;
    wire [63:0] _5544;
    wire [63:0] _500;
    reg [63:0] _5541;
    wire [8:0] _5545;
    wire _5546;
    wire _5547;
    wire [63:0] _5551;
    wire [63:0] _5553;
    wire [63:0] _501;
    reg [63:0] _5550;
    wire [8:0] _5554;
    wire _5555;
    wire _5556;
    wire [63:0] _5560;
    wire [63:0] _5562;
    wire [63:0] _502;
    reg [63:0] _5559;
    wire [8:0] _5563;
    wire _5564;
    wire _5565;
    wire [63:0] _5569;
    wire [63:0] _5571;
    wire [63:0] _503;
    reg [63:0] _5568;
    wire [8:0] _5572;
    wire _5573;
    wire _5574;
    wire [63:0] _5578;
    wire [63:0] _5580;
    wire [63:0] _504;
    reg [63:0] _5577;
    wire [8:0] _5581;
    wire _5582;
    wire _5583;
    wire [63:0] _5587;
    wire [63:0] _5589;
    wire [63:0] _505;
    reg [63:0] _5586;
    wire [8:0] _5590;
    wire _5591;
    wire _5592;
    wire [63:0] _5596;
    wire [63:0] _5598;
    wire [63:0] _506;
    reg [63:0] _5595;
    wire [8:0] _5599;
    wire _5600;
    wire _5601;
    wire [63:0] _5605;
    wire [63:0] _5607;
    wire [63:0] _507;
    reg [63:0] _5604;
    wire [8:0] _5608;
    wire _5609;
    wire _5610;
    wire [63:0] _5614;
    wire [63:0] _5616;
    wire [63:0] _508;
    reg [63:0] _5613;
    wire [8:0] _5617;
    wire _5618;
    wire _5619;
    wire [63:0] _5623;
    wire [63:0] _5625;
    wire [63:0] _509;
    reg [63:0] _5622;
    wire [8:0] _5626;
    wire _5627;
    wire _5628;
    wire [63:0] _5632;
    wire [63:0] _5634;
    wire [63:0] _510;
    reg [63:0] _5631;
    wire [8:0] _5635;
    wire _5636;
    wire _5637;
    wire [63:0] _5641;
    wire [63:0] _5643;
    wire [63:0] _511;
    reg [63:0] _5640;
    wire [8:0] _5644;
    wire _5645;
    wire _5646;
    wire [63:0] _5650;
    wire [63:0] _5652;
    wire [63:0] _512;
    reg [63:0] _5649;
    wire [8:0] _5653;
    wire _5654;
    wire _5655;
    wire [63:0] _5659;
    wire [63:0] _5661;
    wire [63:0] _513;
    reg [63:0] _5658;
    wire [63:0] _515;
    wire [8:0] _5662;
    wire _5663;
    wire _5664;
    wire [63:0] _5668;
    wire [63:0] _5670;
    wire [63:0] _516;
    reg [63:0] _5667;
    reg [63:0] _10304;
    wire _10306;
    wire _10307;
    wire [63:0] _10310;
    wire [63:0] _10312;
    wire [63:0] _10300;
    wire [63:0] _10299;
    reg [63:0] _10296;
    wire _5672;
    wire _5673;
    wire [63:0] _5677;
    wire [63:0] _5679;
    wire [63:0] _517;
    reg [63:0] _5676;
    wire _5681;
    wire _5682;
    wire [63:0] _5686;
    wire [63:0] _5688;
    wire [63:0] _518;
    reg [63:0] _5685;
    wire _5690;
    wire _5691;
    wire [63:0] _5695;
    wire [63:0] _5697;
    wire [63:0] _519;
    reg [63:0] _5694;
    wire _5699;
    wire _5700;
    wire [63:0] _5704;
    wire [63:0] _5706;
    wire [63:0] _520;
    reg [63:0] _5703;
    wire _5708;
    wire _5709;
    wire [63:0] _5713;
    wire [63:0] _5715;
    wire [63:0] _521;
    reg [63:0] _5712;
    wire _5717;
    wire _5718;
    wire [63:0] _5722;
    wire [63:0] _5724;
    wire [63:0] _522;
    reg [63:0] _5721;
    wire _5726;
    wire _5727;
    wire [63:0] _5731;
    wire [63:0] _5733;
    wire [63:0] _523;
    reg [63:0] _5730;
    wire _5735;
    wire _5736;
    wire [63:0] _5740;
    wire [63:0] _5742;
    wire [63:0] _524;
    reg [63:0] _5739;
    wire _5744;
    wire _5745;
    wire [63:0] _5749;
    wire [63:0] _5751;
    wire [63:0] _525;
    reg [63:0] _5748;
    wire _5753;
    wire _5754;
    wire [63:0] _5758;
    wire [63:0] _5760;
    wire [63:0] _526;
    reg [63:0] _5757;
    wire _5762;
    wire _5763;
    wire [63:0] _5767;
    wire [63:0] _5769;
    wire [63:0] _527;
    reg [63:0] _5766;
    wire _5771;
    wire _5772;
    wire [63:0] _5776;
    wire [63:0] _5778;
    wire [63:0] _528;
    reg [63:0] _5775;
    wire _5780;
    wire _5781;
    wire [63:0] _5785;
    wire [63:0] _5787;
    wire [63:0] _529;
    reg [63:0] _5784;
    wire _5789;
    wire _5790;
    wire [63:0] _5794;
    wire [63:0] _5796;
    wire [63:0] _530;
    reg [63:0] _5793;
    wire _5798;
    wire _5799;
    wire [63:0] _5803;
    wire [63:0] _5805;
    wire [63:0] _531;
    reg [63:0] _5802;
    wire _5807;
    wire _5808;
    wire [63:0] _5812;
    wire [63:0] _5814;
    wire [63:0] _532;
    reg [63:0] _5811;
    wire _5816;
    wire _5817;
    wire [63:0] _5821;
    wire [63:0] _5823;
    wire [63:0] _533;
    reg [63:0] _5820;
    wire _5825;
    wire _5826;
    wire [63:0] _5830;
    wire [63:0] _5832;
    wire [63:0] _534;
    reg [63:0] _5829;
    wire _5834;
    wire _5835;
    wire [63:0] _5839;
    wire [63:0] _5841;
    wire [63:0] _535;
    reg [63:0] _5838;
    wire _5843;
    wire _5844;
    wire [63:0] _5848;
    wire [63:0] _5850;
    wire [63:0] _536;
    reg [63:0] _5847;
    wire _5852;
    wire _5853;
    wire [63:0] _5857;
    wire [63:0] _5859;
    wire [63:0] _537;
    reg [63:0] _5856;
    wire _5861;
    wire _5862;
    wire [63:0] _5866;
    wire [63:0] _5868;
    wire [63:0] _538;
    reg [63:0] _5865;
    wire _5870;
    wire _5871;
    wire [63:0] _5875;
    wire [63:0] _5877;
    wire [63:0] _539;
    reg [63:0] _5874;
    wire _5879;
    wire _5880;
    wire [63:0] _5884;
    wire [63:0] _5886;
    wire [63:0] _540;
    reg [63:0] _5883;
    wire _5888;
    wire _5889;
    wire [63:0] _5893;
    wire [63:0] _5895;
    wire [63:0] _541;
    reg [63:0] _5892;
    wire _5897;
    wire _5898;
    wire [63:0] _5902;
    wire [63:0] _5904;
    wire [63:0] _542;
    reg [63:0] _5901;
    wire _5906;
    wire _5907;
    wire [63:0] _5911;
    wire [63:0] _5913;
    wire [63:0] _543;
    reg [63:0] _5910;
    wire _5915;
    wire _5916;
    wire [63:0] _5920;
    wire [63:0] _5922;
    wire [63:0] _544;
    reg [63:0] _5919;
    wire _5924;
    wire _5925;
    wire [63:0] _5929;
    wire [63:0] _5931;
    wire [63:0] _545;
    reg [63:0] _5928;
    wire _5933;
    wire _5934;
    wire [63:0] _5938;
    wire [63:0] _5940;
    wire [63:0] _546;
    reg [63:0] _5937;
    wire _5942;
    wire _5943;
    wire [63:0] _5947;
    wire [63:0] _5949;
    wire [63:0] _547;
    reg [63:0] _5946;
    wire _5951;
    wire _5952;
    wire [63:0] _5956;
    wire [63:0] _5958;
    wire [63:0] _548;
    reg [63:0] _5955;
    wire _5960;
    wire _5961;
    wire [63:0] _5965;
    wire [63:0] _5967;
    wire [63:0] _549;
    reg [63:0] _5964;
    wire _5969;
    wire _5970;
    wire [63:0] _5974;
    wire [63:0] _5976;
    wire [63:0] _550;
    reg [63:0] _5973;
    wire _5978;
    wire _5979;
    wire [63:0] _5983;
    wire [63:0] _5985;
    wire [63:0] _551;
    reg [63:0] _5982;
    wire _5987;
    wire _5988;
    wire [63:0] _5992;
    wire [63:0] _5994;
    wire [63:0] _552;
    reg [63:0] _5991;
    wire _5996;
    wire _5997;
    wire [63:0] _6001;
    wire [63:0] _6003;
    wire [63:0] _553;
    reg [63:0] _6000;
    wire _6005;
    wire _6006;
    wire [63:0] _6010;
    wire [63:0] _6012;
    wire [63:0] _554;
    reg [63:0] _6009;
    wire _6014;
    wire _6015;
    wire [63:0] _6019;
    wire [63:0] _6021;
    wire [63:0] _555;
    reg [63:0] _6018;
    wire _6023;
    wire _6024;
    wire [63:0] _6028;
    wire [63:0] _6030;
    wire [63:0] _556;
    reg [63:0] _6027;
    wire _6032;
    wire _6033;
    wire [63:0] _6037;
    wire [63:0] _6039;
    wire [63:0] _557;
    reg [63:0] _6036;
    wire _6041;
    wire _6042;
    wire [63:0] _6046;
    wire [63:0] _6048;
    wire [63:0] _558;
    reg [63:0] _6045;
    wire _6050;
    wire _6051;
    wire [63:0] _6055;
    wire [63:0] _6057;
    wire [63:0] _559;
    reg [63:0] _6054;
    wire _6059;
    wire _6060;
    wire [63:0] _6064;
    wire [63:0] _6066;
    wire [63:0] _560;
    reg [63:0] _6063;
    wire _6068;
    wire _6069;
    wire [63:0] _6073;
    wire [63:0] _6075;
    wire [63:0] _561;
    reg [63:0] _6072;
    wire _6077;
    wire _6078;
    wire [63:0] _6082;
    wire [63:0] _6084;
    wire [63:0] _562;
    reg [63:0] _6081;
    wire _6086;
    wire _6087;
    wire [63:0] _6091;
    wire [63:0] _6093;
    wire [63:0] _563;
    reg [63:0] _6090;
    wire _6095;
    wire _6096;
    wire [63:0] _6100;
    wire [63:0] _6102;
    wire [63:0] _564;
    reg [63:0] _6099;
    wire _6104;
    wire _6105;
    wire [63:0] _6109;
    wire [63:0] _6111;
    wire [63:0] _565;
    reg [63:0] _6108;
    wire _6113;
    wire _6114;
    wire [63:0] _6118;
    wire [63:0] _6120;
    wire [63:0] _566;
    reg [63:0] _6117;
    wire _6122;
    wire _6123;
    wire [63:0] _6127;
    wire [63:0] _6129;
    wire [63:0] _567;
    reg [63:0] _6126;
    wire _6131;
    wire _6132;
    wire [63:0] _6136;
    wire [63:0] _6138;
    wire [63:0] _568;
    reg [63:0] _6135;
    wire _6140;
    wire _6141;
    wire [63:0] _6145;
    wire [63:0] _6147;
    wire [63:0] _569;
    reg [63:0] _6144;
    wire _6149;
    wire _6150;
    wire [63:0] _6154;
    wire [63:0] _6156;
    wire [63:0] _570;
    reg [63:0] _6153;
    wire _6158;
    wire _6159;
    wire [63:0] _6163;
    wire [63:0] _6165;
    wire [63:0] _571;
    reg [63:0] _6162;
    wire _6167;
    wire _6168;
    wire [63:0] _6172;
    wire [63:0] _6174;
    wire [63:0] _572;
    reg [63:0] _6171;
    wire _6176;
    wire _6177;
    wire [63:0] _6181;
    wire [63:0] _6183;
    wire [63:0] _573;
    reg [63:0] _6180;
    wire _6185;
    wire _6186;
    wire [63:0] _6190;
    wire [63:0] _6192;
    wire [63:0] _574;
    reg [63:0] _6189;
    wire _6194;
    wire _6195;
    wire [63:0] _6199;
    wire [63:0] _6201;
    wire [63:0] _575;
    reg [63:0] _6198;
    wire _6203;
    wire _6204;
    wire [63:0] _6208;
    wire [63:0] _6210;
    wire [63:0] _576;
    reg [63:0] _6207;
    wire _6212;
    wire _6213;
    wire [63:0] _6217;
    wire [63:0] _6219;
    wire [63:0] _577;
    reg [63:0] _6216;
    wire _6221;
    wire _6222;
    wire [63:0] _6226;
    wire [63:0] _6228;
    wire [63:0] _578;
    reg [63:0] _6225;
    wire _6230;
    wire _6231;
    wire [63:0] _6235;
    wire [63:0] _6237;
    wire [63:0] _579;
    reg [63:0] _6234;
    wire _6239;
    wire _6240;
    wire [63:0] _6244;
    wire [63:0] _6246;
    wire [63:0] _580;
    reg [63:0] _6243;
    wire _6248;
    wire _6249;
    wire [63:0] _6253;
    wire [63:0] _6255;
    wire [63:0] _581;
    reg [63:0] _6252;
    wire _6257;
    wire _6258;
    wire [63:0] _6262;
    wire [63:0] _6264;
    wire [63:0] _582;
    reg [63:0] _6261;
    wire _6266;
    wire _6267;
    wire [63:0] _6271;
    wire [63:0] _6273;
    wire [63:0] _583;
    reg [63:0] _6270;
    wire _6275;
    wire _6276;
    wire [63:0] _6280;
    wire [63:0] _6282;
    wire [63:0] _584;
    reg [63:0] _6279;
    wire _6284;
    wire _6285;
    wire [63:0] _6289;
    wire [63:0] _6291;
    wire [63:0] _585;
    reg [63:0] _6288;
    wire _6293;
    wire _6294;
    wire [63:0] _6298;
    wire [63:0] _6300;
    wire [63:0] _586;
    reg [63:0] _6297;
    wire _6302;
    wire _6303;
    wire [63:0] _6307;
    wire [63:0] _6309;
    wire [63:0] _587;
    reg [63:0] _6306;
    wire _6311;
    wire _6312;
    wire [63:0] _6316;
    wire [63:0] _6318;
    wire [63:0] _588;
    reg [63:0] _6315;
    wire _6320;
    wire _6321;
    wire [63:0] _6325;
    wire [63:0] _6327;
    wire [63:0] _589;
    reg [63:0] _6324;
    wire _6329;
    wire _6330;
    wire [63:0] _6334;
    wire [63:0] _6336;
    wire [63:0] _590;
    reg [63:0] _6333;
    wire _6338;
    wire _6339;
    wire [63:0] _6343;
    wire [63:0] _6345;
    wire [63:0] _591;
    reg [63:0] _6342;
    wire _6347;
    wire _6348;
    wire [63:0] _6352;
    wire [63:0] _6354;
    wire [63:0] _592;
    reg [63:0] _6351;
    wire _6356;
    wire _6357;
    wire [63:0] _6361;
    wire [63:0] _6363;
    wire [63:0] _593;
    reg [63:0] _6360;
    wire _6365;
    wire _6366;
    wire [63:0] _6370;
    wire [63:0] _6372;
    wire [63:0] _594;
    reg [63:0] _6369;
    wire _6374;
    wire _6375;
    wire [63:0] _6379;
    wire [63:0] _6381;
    wire [63:0] _595;
    reg [63:0] _6378;
    wire _6383;
    wire _6384;
    wire [63:0] _6388;
    wire [63:0] _6390;
    wire [63:0] _596;
    reg [63:0] _6387;
    wire _6392;
    wire _6393;
    wire [63:0] _6397;
    wire [63:0] _6399;
    wire [63:0] _597;
    reg [63:0] _6396;
    wire _6401;
    wire _6402;
    wire [63:0] _6406;
    wire [63:0] _6408;
    wire [63:0] _598;
    reg [63:0] _6405;
    wire _6410;
    wire _6411;
    wire [63:0] _6415;
    wire [63:0] _6417;
    wire [63:0] _599;
    reg [63:0] _6414;
    wire _6419;
    wire _6420;
    wire [63:0] _6424;
    wire [63:0] _6426;
    wire [63:0] _600;
    reg [63:0] _6423;
    wire _6428;
    wire _6429;
    wire [63:0] _6433;
    wire [63:0] _6435;
    wire [63:0] _601;
    reg [63:0] _6432;
    wire _6437;
    wire _6438;
    wire [63:0] _6442;
    wire [63:0] _6444;
    wire [63:0] _602;
    reg [63:0] _6441;
    wire _6446;
    wire _6447;
    wire [63:0] _6451;
    wire [63:0] _6453;
    wire [63:0] _603;
    reg [63:0] _6450;
    wire _6455;
    wire _6456;
    wire [63:0] _6460;
    wire [63:0] _6462;
    wire [63:0] _604;
    reg [63:0] _6459;
    wire _6464;
    wire _6465;
    wire [63:0] _6469;
    wire [63:0] _6471;
    wire [63:0] _605;
    reg [63:0] _6468;
    wire _6473;
    wire _6474;
    wire [63:0] _6478;
    wire [63:0] _6480;
    wire [63:0] _606;
    reg [63:0] _6477;
    wire _6482;
    wire _6483;
    wire [63:0] _6487;
    wire [63:0] _6489;
    wire [63:0] _607;
    reg [63:0] _6486;
    wire _6491;
    wire _6492;
    wire [63:0] _6496;
    wire [63:0] _6498;
    wire [63:0] _608;
    reg [63:0] _6495;
    wire _6500;
    wire _6501;
    wire [63:0] _6505;
    wire [63:0] _6507;
    wire [63:0] _609;
    reg [63:0] _6504;
    wire _6509;
    wire _6510;
    wire [63:0] _6514;
    wire [63:0] _6516;
    wire [63:0] _610;
    reg [63:0] _6513;
    wire _6518;
    wire _6519;
    wire [63:0] _6523;
    wire [63:0] _6525;
    wire [63:0] _611;
    reg [63:0] _6522;
    wire _6527;
    wire _6528;
    wire [63:0] _6532;
    wire [63:0] _6534;
    wire [63:0] _612;
    reg [63:0] _6531;
    wire _6536;
    wire _6537;
    wire [63:0] _6541;
    wire [63:0] _6543;
    wire [63:0] _613;
    reg [63:0] _6540;
    wire _6545;
    wire _6546;
    wire [63:0] _6550;
    wire [63:0] _6552;
    wire [63:0] _614;
    reg [63:0] _6549;
    wire _6554;
    wire _6555;
    wire [63:0] _6559;
    wire [63:0] _6561;
    wire [63:0] _615;
    reg [63:0] _6558;
    wire _6563;
    wire _6564;
    wire [63:0] _6568;
    wire [63:0] _6570;
    wire [63:0] _616;
    reg [63:0] _6567;
    wire _6572;
    wire _6573;
    wire [63:0] _6577;
    wire [63:0] _6579;
    wire [63:0] _617;
    reg [63:0] _6576;
    wire _6581;
    wire _6582;
    wire [63:0] _6586;
    wire [63:0] _6588;
    wire [63:0] _618;
    reg [63:0] _6585;
    wire _6590;
    wire _6591;
    wire [63:0] _6595;
    wire [63:0] _6597;
    wire [63:0] _619;
    reg [63:0] _6594;
    wire _6599;
    wire _6600;
    wire [63:0] _6604;
    wire [63:0] _6606;
    wire [63:0] _620;
    reg [63:0] _6603;
    wire _6608;
    wire _6609;
    wire [63:0] _6613;
    wire [63:0] _6615;
    wire [63:0] _621;
    reg [63:0] _6612;
    wire _6617;
    wire _6618;
    wire [63:0] _6622;
    wire [63:0] _6624;
    wire [63:0] _622;
    reg [63:0] _6621;
    wire _6626;
    wire _6627;
    wire [63:0] _6631;
    wire [63:0] _6633;
    wire [63:0] _623;
    reg [63:0] _6630;
    wire _6635;
    wire _6636;
    wire [63:0] _6640;
    wire [63:0] _6642;
    wire [63:0] _624;
    reg [63:0] _6639;
    wire _6644;
    wire _6645;
    wire [63:0] _6649;
    wire [63:0] _6651;
    wire [63:0] _625;
    reg [63:0] _6648;
    wire _6653;
    wire _6654;
    wire [63:0] _6658;
    wire [63:0] _6660;
    wire [63:0] _626;
    reg [63:0] _6657;
    wire _6662;
    wire _6663;
    wire [63:0] _6667;
    wire [63:0] _6669;
    wire [63:0] _627;
    reg [63:0] _6666;
    wire _6671;
    wire _6672;
    wire [63:0] _6676;
    wire [63:0] _6678;
    wire [63:0] _628;
    reg [63:0] _6675;
    wire _6680;
    wire _6681;
    wire [63:0] _6685;
    wire [63:0] _6687;
    wire [63:0] _629;
    reg [63:0] _6684;
    wire _6689;
    wire _6690;
    wire [63:0] _6694;
    wire [63:0] _6696;
    wire [63:0] _630;
    reg [63:0] _6693;
    wire _6698;
    wire _6699;
    wire [63:0] _6703;
    wire [63:0] _6705;
    wire [63:0] _631;
    reg [63:0] _6702;
    wire _6707;
    wire _6708;
    wire [63:0] _6712;
    wire [63:0] _6714;
    wire [63:0] _632;
    reg [63:0] _6711;
    wire _6716;
    wire _6717;
    wire [63:0] _6721;
    wire [63:0] _6723;
    wire [63:0] _633;
    reg [63:0] _6720;
    wire _6725;
    wire _6726;
    wire [63:0] _6730;
    wire [63:0] _6732;
    wire [63:0] _634;
    reg [63:0] _6729;
    wire _6734;
    wire _6735;
    wire [63:0] _6739;
    wire [63:0] _6741;
    wire [63:0] _635;
    reg [63:0] _6738;
    wire _6743;
    wire _6744;
    wire [63:0] _6748;
    wire [63:0] _6750;
    wire [63:0] _636;
    reg [63:0] _6747;
    wire _6752;
    wire _6753;
    wire [63:0] _6757;
    wire [63:0] _6759;
    wire [63:0] _637;
    reg [63:0] _6756;
    wire _6761;
    wire _6762;
    wire [63:0] _6766;
    wire [63:0] _6768;
    wire [63:0] _638;
    reg [63:0] _6765;
    wire _6770;
    wire _6771;
    wire [63:0] _6775;
    wire [63:0] _6777;
    wire [63:0] _639;
    reg [63:0] _6774;
    wire _6779;
    wire _6780;
    wire [63:0] _6784;
    wire [63:0] _6786;
    wire [63:0] _640;
    reg [63:0] _6783;
    wire _6788;
    wire _6789;
    wire [63:0] _6793;
    wire [63:0] _6795;
    wire [63:0] _641;
    reg [63:0] _6792;
    wire _6797;
    wire _6798;
    wire [63:0] _6802;
    wire [63:0] _6804;
    wire [63:0] _642;
    reg [63:0] _6801;
    wire _6806;
    wire _6807;
    wire [63:0] _6811;
    wire [63:0] _6813;
    wire [63:0] _643;
    reg [63:0] _6810;
    wire _6815;
    wire _6816;
    wire [63:0] _6820;
    wire [63:0] _6822;
    wire [63:0] _644;
    reg [63:0] _6819;
    wire _6824;
    wire _6825;
    wire [63:0] _6829;
    wire [63:0] _6831;
    wire [63:0] _645;
    reg [63:0] _6828;
    wire _6833;
    wire _6834;
    wire [63:0] _6838;
    wire [63:0] _6840;
    wire [63:0] _646;
    reg [63:0] _6837;
    wire _6842;
    wire _6843;
    wire [63:0] _6847;
    wire [63:0] _6849;
    wire [63:0] _647;
    reg [63:0] _6846;
    wire _6851;
    wire _6852;
    wire [63:0] _6856;
    wire [63:0] _6858;
    wire [63:0] _648;
    reg [63:0] _6855;
    wire _6860;
    wire _6861;
    wire [63:0] _6865;
    wire [63:0] _6867;
    wire [63:0] _649;
    reg [63:0] _6864;
    wire _6869;
    wire _6870;
    wire [63:0] _6874;
    wire [63:0] _6876;
    wire [63:0] _650;
    reg [63:0] _6873;
    wire _6878;
    wire _6879;
    wire [63:0] _6883;
    wire [63:0] _6885;
    wire [63:0] _651;
    reg [63:0] _6882;
    wire _6887;
    wire _6888;
    wire [63:0] _6892;
    wire [63:0] _6894;
    wire [63:0] _652;
    reg [63:0] _6891;
    wire _6896;
    wire _6897;
    wire [63:0] _6901;
    wire [63:0] _6903;
    wire [63:0] _653;
    reg [63:0] _6900;
    wire _6905;
    wire _6906;
    wire [63:0] _6910;
    wire [63:0] _6912;
    wire [63:0] _654;
    reg [63:0] _6909;
    wire _6914;
    wire _6915;
    wire [63:0] _6919;
    wire [63:0] _6921;
    wire [63:0] _655;
    reg [63:0] _6918;
    wire _6923;
    wire _6924;
    wire [63:0] _6928;
    wire [63:0] _6930;
    wire [63:0] _656;
    reg [63:0] _6927;
    wire _6932;
    wire _6933;
    wire [63:0] _6937;
    wire [63:0] _6939;
    wire [63:0] _657;
    reg [63:0] _6936;
    wire _6941;
    wire _6942;
    wire [63:0] _6946;
    wire [63:0] _6948;
    wire [63:0] _658;
    reg [63:0] _6945;
    wire _6950;
    wire _6951;
    wire [63:0] _6955;
    wire [63:0] _6957;
    wire [63:0] _659;
    reg [63:0] _6954;
    wire _6959;
    wire _6960;
    wire [63:0] _6964;
    wire [63:0] _6966;
    wire [63:0] _660;
    reg [63:0] _6963;
    wire _6968;
    wire _6969;
    wire [63:0] _6973;
    wire [63:0] _6975;
    wire [63:0] _661;
    reg [63:0] _6972;
    wire _6977;
    wire _6978;
    wire [63:0] _6982;
    wire [63:0] _6984;
    wire [63:0] _662;
    reg [63:0] _6981;
    wire _6986;
    wire _6987;
    wire [63:0] _6991;
    wire [63:0] _6993;
    wire [63:0] _663;
    reg [63:0] _6990;
    wire _6995;
    wire _6996;
    wire [63:0] _7000;
    wire [63:0] _7002;
    wire [63:0] _664;
    reg [63:0] _6999;
    wire _7004;
    wire _7005;
    wire [63:0] _7009;
    wire [63:0] _7011;
    wire [63:0] _665;
    reg [63:0] _7008;
    wire _7013;
    wire _7014;
    wire [63:0] _7018;
    wire [63:0] _7020;
    wire [63:0] _666;
    reg [63:0] _7017;
    wire _7022;
    wire _7023;
    wire [63:0] _7027;
    wire [63:0] _7029;
    wire [63:0] _667;
    reg [63:0] _7026;
    wire _7031;
    wire _7032;
    wire [63:0] _7036;
    wire [63:0] _7038;
    wire [63:0] _668;
    reg [63:0] _7035;
    wire _7040;
    wire _7041;
    wire [63:0] _7045;
    wire [63:0] _7047;
    wire [63:0] _669;
    reg [63:0] _7044;
    wire _7049;
    wire _7050;
    wire [63:0] _7054;
    wire [63:0] _7056;
    wire [63:0] _670;
    reg [63:0] _7053;
    wire _7058;
    wire _7059;
    wire [63:0] _7063;
    wire [63:0] _7065;
    wire [63:0] _671;
    reg [63:0] _7062;
    wire _7067;
    wire _7068;
    wire [63:0] _7072;
    wire [63:0] _7074;
    wire [63:0] _672;
    reg [63:0] _7071;
    wire _7076;
    wire _7077;
    wire [63:0] _7081;
    wire [63:0] _7083;
    wire [63:0] _673;
    reg [63:0] _7080;
    wire _7085;
    wire _7086;
    wire [63:0] _7090;
    wire [63:0] _7092;
    wire [63:0] _674;
    reg [63:0] _7089;
    wire _7094;
    wire _7095;
    wire [63:0] _7099;
    wire [63:0] _7101;
    wire [63:0] _675;
    reg [63:0] _7098;
    wire _7103;
    wire _7104;
    wire [63:0] _7108;
    wire [63:0] _7110;
    wire [63:0] _676;
    reg [63:0] _7107;
    wire _7112;
    wire _7113;
    wire [63:0] _7117;
    wire [63:0] _7119;
    wire [63:0] _677;
    reg [63:0] _7116;
    wire _7121;
    wire _7122;
    wire [63:0] _7126;
    wire [63:0] _7128;
    wire [63:0] _678;
    reg [63:0] _7125;
    wire _7130;
    wire _7131;
    wire [63:0] _7135;
    wire [63:0] _7137;
    wire [63:0] _679;
    reg [63:0] _7134;
    wire _7139;
    wire _7140;
    wire [63:0] _7144;
    wire [63:0] _7146;
    wire [63:0] _680;
    reg [63:0] _7143;
    wire _7148;
    wire _7149;
    wire [63:0] _7153;
    wire [63:0] _7155;
    wire [63:0] _681;
    reg [63:0] _7152;
    wire _7157;
    wire _7158;
    wire [63:0] _7162;
    wire [63:0] _7164;
    wire [63:0] _682;
    reg [63:0] _7161;
    wire _7166;
    wire _7167;
    wire [63:0] _7171;
    wire [63:0] _7173;
    wire [63:0] _683;
    reg [63:0] _7170;
    wire _7175;
    wire _7176;
    wire [63:0] _7180;
    wire [63:0] _7182;
    wire [63:0] _684;
    reg [63:0] _7179;
    wire _7184;
    wire _7185;
    wire [63:0] _7189;
    wire [63:0] _7191;
    wire [63:0] _685;
    reg [63:0] _7188;
    wire _7193;
    wire _7194;
    wire [63:0] _7198;
    wire [63:0] _7200;
    wire [63:0] _686;
    reg [63:0] _7197;
    wire _7202;
    wire _7203;
    wire [63:0] _7207;
    wire [63:0] _7209;
    wire [63:0] _687;
    reg [63:0] _7206;
    wire _7211;
    wire _7212;
    wire [63:0] _7216;
    wire [63:0] _7218;
    wire [63:0] _688;
    reg [63:0] _7215;
    wire _7220;
    wire _7221;
    wire [63:0] _7225;
    wire [63:0] _7227;
    wire [63:0] _689;
    reg [63:0] _7224;
    wire _7229;
    wire _7230;
    wire [63:0] _7234;
    wire [63:0] _7236;
    wire [63:0] _690;
    reg [63:0] _7233;
    wire _7238;
    wire _7239;
    wire [63:0] _7243;
    wire [63:0] _7245;
    wire [63:0] _691;
    reg [63:0] _7242;
    wire _7247;
    wire _7248;
    wire [63:0] _7252;
    wire [63:0] _7254;
    wire [63:0] _692;
    reg [63:0] _7251;
    wire _7256;
    wire _7257;
    wire [63:0] _7261;
    wire [63:0] _7263;
    wire [63:0] _693;
    reg [63:0] _7260;
    wire _7265;
    wire _7266;
    wire [63:0] _7270;
    wire [63:0] _7272;
    wire [63:0] _694;
    reg [63:0] _7269;
    wire _7274;
    wire _7275;
    wire [63:0] _7279;
    wire [63:0] _7281;
    wire [63:0] _695;
    reg [63:0] _7278;
    wire _7283;
    wire _7284;
    wire [63:0] _7288;
    wire [63:0] _7290;
    wire [63:0] _696;
    reg [63:0] _7287;
    wire _7292;
    wire _7293;
    wire [63:0] _7297;
    wire [63:0] _7299;
    wire [63:0] _697;
    reg [63:0] _7296;
    wire _7301;
    wire _7302;
    wire [63:0] _7306;
    wire [63:0] _7308;
    wire [63:0] _698;
    reg [63:0] _7305;
    wire _7310;
    wire _7311;
    wire [63:0] _7315;
    wire [63:0] _7317;
    wire [63:0] _699;
    reg [63:0] _7314;
    wire _7319;
    wire _7320;
    wire [63:0] _7324;
    wire [63:0] _7326;
    wire [63:0] _700;
    reg [63:0] _7323;
    wire _7328;
    wire _7329;
    wire [63:0] _7333;
    wire [63:0] _7335;
    wire [63:0] _701;
    reg [63:0] _7332;
    wire _7337;
    wire _7338;
    wire [63:0] _7342;
    wire [63:0] _7344;
    wire [63:0] _702;
    reg [63:0] _7341;
    wire _7346;
    wire _7347;
    wire [63:0] _7351;
    wire [63:0] _7353;
    wire [63:0] _703;
    reg [63:0] _7350;
    wire _7355;
    wire _7356;
    wire [63:0] _7360;
    wire [63:0] _7362;
    wire [63:0] _704;
    reg [63:0] _7359;
    wire _7364;
    wire _7365;
    wire [63:0] _7369;
    wire [63:0] _7371;
    wire [63:0] _705;
    reg [63:0] _7368;
    wire _7373;
    wire _7374;
    wire [63:0] _7378;
    wire [63:0] _7380;
    wire [63:0] _706;
    reg [63:0] _7377;
    wire _7382;
    wire _7383;
    wire [63:0] _7387;
    wire [63:0] _7389;
    wire [63:0] _707;
    reg [63:0] _7386;
    wire _7391;
    wire _7392;
    wire [63:0] _7396;
    wire [63:0] _7398;
    wire [63:0] _708;
    reg [63:0] _7395;
    wire _7400;
    wire _7401;
    wire [63:0] _7405;
    wire [63:0] _7407;
    wire [63:0] _709;
    reg [63:0] _7404;
    wire _7409;
    wire _7410;
    wire [63:0] _7414;
    wire [63:0] _7416;
    wire [63:0] _710;
    reg [63:0] _7413;
    wire _7418;
    wire _7419;
    wire [63:0] _7423;
    wire [63:0] _7425;
    wire [63:0] _711;
    reg [63:0] _7422;
    wire _7427;
    wire _7428;
    wire [63:0] _7432;
    wire [63:0] _7434;
    wire [63:0] _712;
    reg [63:0] _7431;
    wire _7436;
    wire _7437;
    wire [63:0] _7441;
    wire [63:0] _7443;
    wire [63:0] _713;
    reg [63:0] _7440;
    wire _7445;
    wire _7446;
    wire [63:0] _7450;
    wire [63:0] _7452;
    wire [63:0] _714;
    reg [63:0] _7449;
    wire _7454;
    wire _7455;
    wire [63:0] _7459;
    wire [63:0] _7461;
    wire [63:0] _715;
    reg [63:0] _7458;
    wire _7463;
    wire _7464;
    wire [63:0] _7468;
    wire [63:0] _7470;
    wire [63:0] _716;
    reg [63:0] _7467;
    wire _7472;
    wire _7473;
    wire [63:0] _7477;
    wire [63:0] _7479;
    wire [63:0] _717;
    reg [63:0] _7476;
    wire _7481;
    wire _7482;
    wire [63:0] _7486;
    wire [63:0] _7488;
    wire [63:0] _718;
    reg [63:0] _7485;
    wire _7490;
    wire _7491;
    wire [63:0] _7495;
    wire [63:0] _7497;
    wire [63:0] _719;
    reg [63:0] _7494;
    wire _7499;
    wire _7500;
    wire [63:0] _7504;
    wire [63:0] _7506;
    wire [63:0] _720;
    reg [63:0] _7503;
    wire _7508;
    wire _7509;
    wire [63:0] _7513;
    wire [63:0] _7515;
    wire [63:0] _721;
    reg [63:0] _7512;
    wire _7517;
    wire _7518;
    wire [63:0] _7522;
    wire [63:0] _7524;
    wire [63:0] _722;
    reg [63:0] _7521;
    wire _7526;
    wire _7527;
    wire [63:0] _7531;
    wire [63:0] _7533;
    wire [63:0] _723;
    reg [63:0] _7530;
    wire _7535;
    wire _7536;
    wire [63:0] _7540;
    wire [63:0] _7542;
    wire [63:0] _724;
    reg [63:0] _7539;
    wire _7544;
    wire _7545;
    wire [63:0] _7549;
    wire [63:0] _7551;
    wire [63:0] _725;
    reg [63:0] _7548;
    wire _7553;
    wire _7554;
    wire [63:0] _7558;
    wire [63:0] _7560;
    wire [63:0] _726;
    reg [63:0] _7557;
    wire _7562;
    wire _7563;
    wire [63:0] _7567;
    wire [63:0] _7569;
    wire [63:0] _727;
    reg [63:0] _7566;
    wire _7571;
    wire _7572;
    wire [63:0] _7576;
    wire [63:0] _7578;
    wire [63:0] _728;
    reg [63:0] _7575;
    wire _7580;
    wire _7581;
    wire [63:0] _7585;
    wire [63:0] _7587;
    wire [63:0] _729;
    reg [63:0] _7584;
    wire _7589;
    wire _7590;
    wire [63:0] _7594;
    wire [63:0] _7596;
    wire [63:0] _730;
    reg [63:0] _7593;
    wire _7598;
    wire _7599;
    wire [63:0] _7603;
    wire [63:0] _7605;
    wire [63:0] _731;
    reg [63:0] _7602;
    wire _7607;
    wire _7608;
    wire [63:0] _7612;
    wire [63:0] _7614;
    wire [63:0] _732;
    reg [63:0] _7611;
    wire _7616;
    wire _7617;
    wire [63:0] _7621;
    wire [63:0] _7623;
    wire [63:0] _733;
    reg [63:0] _7620;
    wire _7625;
    wire _7626;
    wire [63:0] _7630;
    wire [63:0] _7632;
    wire [63:0] _734;
    reg [63:0] _7629;
    wire _7634;
    wire _7635;
    wire [63:0] _7639;
    wire [63:0] _7641;
    wire [63:0] _735;
    reg [63:0] _7638;
    wire _7643;
    wire _7644;
    wire [63:0] _7648;
    wire [63:0] _7650;
    wire [63:0] _736;
    reg [63:0] _7647;
    wire _7652;
    wire _7653;
    wire [63:0] _7657;
    wire [63:0] _7659;
    wire [63:0] _737;
    reg [63:0] _7656;
    wire _7661;
    wire _7662;
    wire [63:0] _7666;
    wire [63:0] _7668;
    wire [63:0] _738;
    reg [63:0] _7665;
    wire _7670;
    wire _7671;
    wire [63:0] _7675;
    wire [63:0] _7677;
    wire [63:0] _739;
    reg [63:0] _7674;
    wire _7679;
    wire _7680;
    wire [63:0] _7684;
    wire [63:0] _7686;
    wire [63:0] _740;
    reg [63:0] _7683;
    wire _7688;
    wire _7689;
    wire [63:0] _7693;
    wire [63:0] _7695;
    wire [63:0] _741;
    reg [63:0] _7692;
    wire _7697;
    wire _7698;
    wire [63:0] _7702;
    wire [63:0] _7704;
    wire [63:0] _742;
    reg [63:0] _7701;
    wire _7706;
    wire _7707;
    wire [63:0] _7711;
    wire [63:0] _7713;
    wire [63:0] _743;
    reg [63:0] _7710;
    wire _7715;
    wire _7716;
    wire [63:0] _7720;
    wire [63:0] _7722;
    wire [63:0] _744;
    reg [63:0] _7719;
    wire _7724;
    wire _7725;
    wire [63:0] _7729;
    wire [63:0] _7731;
    wire [63:0] _745;
    reg [63:0] _7728;
    wire _7733;
    wire _7734;
    wire [63:0] _7738;
    wire [63:0] _7740;
    wire [63:0] _746;
    reg [63:0] _7737;
    wire _7742;
    wire _7743;
    wire [63:0] _7747;
    wire [63:0] _7749;
    wire [63:0] _747;
    reg [63:0] _7746;
    wire _7751;
    wire _7752;
    wire [63:0] _7756;
    wire [63:0] _7758;
    wire [63:0] _748;
    reg [63:0] _7755;
    wire _7760;
    wire _7761;
    wire [63:0] _7765;
    wire [63:0] _7767;
    wire [63:0] _749;
    reg [63:0] _7764;
    wire _7769;
    wire _7770;
    wire [63:0] _7774;
    wire [63:0] _7776;
    wire [63:0] _750;
    reg [63:0] _7773;
    wire _7778;
    wire _7779;
    wire [63:0] _7783;
    wire [63:0] _7785;
    wire [63:0] _751;
    reg [63:0] _7782;
    wire _7787;
    wire _7788;
    wire [63:0] _7792;
    wire [63:0] _7794;
    wire [63:0] _752;
    reg [63:0] _7791;
    wire _7796;
    wire _7797;
    wire [63:0] _7801;
    wire [63:0] _7803;
    wire [63:0] _753;
    reg [63:0] _7800;
    wire _7805;
    wire _7806;
    wire [63:0] _7810;
    wire [63:0] _7812;
    wire [63:0] _754;
    reg [63:0] _7809;
    wire _7814;
    wire _7815;
    wire [63:0] _7819;
    wire [63:0] _7821;
    wire [63:0] _755;
    reg [63:0] _7818;
    wire _7823;
    wire _7824;
    wire [63:0] _7828;
    wire [63:0] _7830;
    wire [63:0] _756;
    reg [63:0] _7827;
    wire _7832;
    wire _7833;
    wire [63:0] _7837;
    wire [63:0] _7839;
    wire [63:0] _757;
    reg [63:0] _7836;
    wire _7841;
    wire _7842;
    wire [63:0] _7846;
    wire [63:0] _7848;
    wire [63:0] _758;
    reg [63:0] _7845;
    wire _7850;
    wire _7851;
    wire [63:0] _7855;
    wire [63:0] _7857;
    wire [63:0] _759;
    reg [63:0] _7854;
    wire _7859;
    wire _7860;
    wire [63:0] _7864;
    wire [63:0] _7866;
    wire [63:0] _760;
    reg [63:0] _7863;
    wire _7868;
    wire _7869;
    wire [63:0] _7873;
    wire [63:0] _7875;
    wire [63:0] _761;
    reg [63:0] _7872;
    wire _7877;
    wire _7878;
    wire [63:0] _7882;
    wire [63:0] _7884;
    wire [63:0] _762;
    reg [63:0] _7881;
    wire _7886;
    wire _7887;
    wire [63:0] _7891;
    wire [63:0] _7893;
    wire [63:0] _763;
    reg [63:0] _7890;
    wire _7895;
    wire _7896;
    wire [63:0] _7900;
    wire [63:0] _7902;
    wire [63:0] _764;
    reg [63:0] _7899;
    wire _7904;
    wire _7905;
    wire [63:0] _7909;
    wire [63:0] _7911;
    wire [63:0] _765;
    reg [63:0] _7908;
    wire _7913;
    wire _7914;
    wire [63:0] _7918;
    wire [63:0] _7920;
    wire [63:0] _766;
    reg [63:0] _7917;
    wire _7922;
    wire _7923;
    wire [63:0] _7927;
    wire [63:0] _7929;
    wire [63:0] _767;
    reg [63:0] _7926;
    wire _7931;
    wire _7932;
    wire [63:0] _7936;
    wire [63:0] _7938;
    wire [63:0] _768;
    reg [63:0] _7935;
    wire _7940;
    wire _7941;
    wire [63:0] _7945;
    wire [63:0] _7947;
    wire [63:0] _769;
    reg [63:0] _7944;
    wire _7949;
    wire _7950;
    wire [63:0] _7954;
    wire [63:0] _7956;
    wire [63:0] _770;
    reg [63:0] _7953;
    wire _7958;
    wire _7959;
    wire [63:0] _7963;
    wire [63:0] _7965;
    wire [63:0] _771;
    reg [63:0] _7962;
    wire _7967;
    wire _7968;
    wire [63:0] _7972;
    wire [63:0] _7974;
    wire [63:0] _772;
    reg [63:0] _7971;
    wire _7976;
    wire _7977;
    wire [63:0] _7981;
    wire [63:0] _7983;
    wire [63:0] _773;
    reg [63:0] _7980;
    wire _7985;
    wire _7986;
    wire [63:0] _7990;
    wire [63:0] _7992;
    wire [63:0] _774;
    reg [63:0] _7989;
    wire _7994;
    wire _7995;
    wire [63:0] _7999;
    wire [63:0] _8001;
    wire [63:0] _775;
    reg [63:0] _7998;
    wire _8003;
    wire _8004;
    wire [63:0] _8008;
    wire [63:0] _8010;
    wire [63:0] _776;
    reg [63:0] _8007;
    wire _8012;
    wire _8013;
    wire [63:0] _8017;
    wire [63:0] _8019;
    wire [63:0] _777;
    reg [63:0] _8016;
    wire _8021;
    wire _8022;
    wire [63:0] _8026;
    wire [63:0] _8028;
    wire [63:0] _778;
    reg [63:0] _8025;
    wire _8030;
    wire _8031;
    wire [63:0] _8035;
    wire [63:0] _8037;
    wire [63:0] _779;
    reg [63:0] _8034;
    wire _8039;
    wire _8040;
    wire [63:0] _8044;
    wire [63:0] _8046;
    wire [63:0] _780;
    reg [63:0] _8043;
    wire _8048;
    wire _8049;
    wire [63:0] _8053;
    wire [63:0] _8055;
    wire [63:0] _781;
    reg [63:0] _8052;
    wire _8057;
    wire _8058;
    wire [63:0] _8062;
    wire [63:0] _8064;
    wire [63:0] _782;
    reg [63:0] _8061;
    wire _8066;
    wire _8067;
    wire [63:0] _8071;
    wire [63:0] _8073;
    wire [63:0] _783;
    reg [63:0] _8070;
    wire _8075;
    wire _8076;
    wire [63:0] _8080;
    wire [63:0] _8082;
    wire [63:0] _784;
    reg [63:0] _8079;
    wire _8084;
    wire _8085;
    wire [63:0] _8089;
    wire [63:0] _8091;
    wire [63:0] _785;
    reg [63:0] _8088;
    wire _8093;
    wire _8094;
    wire [63:0] _8098;
    wire [63:0] _8100;
    wire [63:0] _786;
    reg [63:0] _8097;
    wire _8102;
    wire _8103;
    wire [63:0] _8107;
    wire [63:0] _8109;
    wire [63:0] _787;
    reg [63:0] _8106;
    wire _8111;
    wire _8112;
    wire [63:0] _8116;
    wire [63:0] _8118;
    wire [63:0] _788;
    reg [63:0] _8115;
    wire _8120;
    wire _8121;
    wire [63:0] _8125;
    wire [63:0] _8127;
    wire [63:0] _789;
    reg [63:0] _8124;
    wire _8129;
    wire _8130;
    wire [63:0] _8134;
    wire [63:0] _8136;
    wire [63:0] _790;
    reg [63:0] _8133;
    wire _8138;
    wire _8139;
    wire [63:0] _8143;
    wire [63:0] _8145;
    wire [63:0] _791;
    reg [63:0] _8142;
    wire _8147;
    wire _8148;
    wire [63:0] _8152;
    wire [63:0] _8154;
    wire [63:0] _792;
    reg [63:0] _8151;
    wire _8156;
    wire _8157;
    wire [63:0] _8161;
    wire [63:0] _8163;
    wire [63:0] _793;
    reg [63:0] _8160;
    wire _8165;
    wire _8166;
    wire [63:0] _8170;
    wire [63:0] _8172;
    wire [63:0] _794;
    reg [63:0] _8169;
    wire _8174;
    wire _8175;
    wire [63:0] _8179;
    wire [63:0] _8181;
    wire [63:0] _795;
    reg [63:0] _8178;
    wire _8183;
    wire _8184;
    wire [63:0] _8188;
    wire [63:0] _8190;
    wire [63:0] _796;
    reg [63:0] _8187;
    wire _8192;
    wire _8193;
    wire [63:0] _8197;
    wire [63:0] _8199;
    wire [63:0] _797;
    reg [63:0] _8196;
    wire _8201;
    wire _8202;
    wire [63:0] _8206;
    wire [63:0] _8208;
    wire [63:0] _798;
    reg [63:0] _8205;
    wire _8210;
    wire _8211;
    wire [63:0] _8215;
    wire [63:0] _8217;
    wire [63:0] _799;
    reg [63:0] _8214;
    wire _8219;
    wire _8220;
    wire [63:0] _8224;
    wire [63:0] _8226;
    wire [63:0] _800;
    reg [63:0] _8223;
    wire _8228;
    wire _8229;
    wire [63:0] _8233;
    wire [63:0] _8235;
    wire [63:0] _801;
    reg [63:0] _8232;
    wire _8237;
    wire _8238;
    wire [63:0] _8242;
    wire [63:0] _8244;
    wire [63:0] _802;
    reg [63:0] _8241;
    wire _8246;
    wire _8247;
    wire [63:0] _8251;
    wire [63:0] _8253;
    wire [63:0] _803;
    reg [63:0] _8250;
    wire _8255;
    wire _8256;
    wire [63:0] _8260;
    wire [63:0] _8262;
    wire [63:0] _804;
    reg [63:0] _8259;
    wire _8264;
    wire _8265;
    wire [63:0] _8269;
    wire [63:0] _8271;
    wire [63:0] _805;
    reg [63:0] _8268;
    wire _8273;
    wire _8274;
    wire [63:0] _8278;
    wire [63:0] _8280;
    wire [63:0] _806;
    reg [63:0] _8277;
    wire _8282;
    wire _8283;
    wire [63:0] _8287;
    wire [63:0] _8289;
    wire [63:0] _807;
    reg [63:0] _8286;
    wire _8291;
    wire _8292;
    wire [63:0] _8296;
    wire [63:0] _8298;
    wire [63:0] _808;
    reg [63:0] _8295;
    wire _8300;
    wire _8301;
    wire [63:0] _8305;
    wire [63:0] _8307;
    wire [63:0] _809;
    reg [63:0] _8304;
    wire _8309;
    wire _8310;
    wire [63:0] _8314;
    wire [63:0] _8316;
    wire [63:0] _810;
    reg [63:0] _8313;
    wire _8318;
    wire _8319;
    wire [63:0] _8323;
    wire [63:0] _8325;
    wire [63:0] _811;
    reg [63:0] _8322;
    wire _8327;
    wire _8328;
    wire [63:0] _8332;
    wire [63:0] _8334;
    wire [63:0] _812;
    reg [63:0] _8331;
    wire _8336;
    wire _8337;
    wire [63:0] _8341;
    wire [63:0] _8343;
    wire [63:0] _813;
    reg [63:0] _8340;
    wire _8345;
    wire _8346;
    wire [63:0] _8350;
    wire [63:0] _8352;
    wire [63:0] _814;
    reg [63:0] _8349;
    wire _8354;
    wire _8355;
    wire [63:0] _8359;
    wire [63:0] _8361;
    wire [63:0] _815;
    reg [63:0] _8358;
    wire _8363;
    wire _8364;
    wire [63:0] _8368;
    wire [63:0] _8370;
    wire [63:0] _816;
    reg [63:0] _8367;
    wire _8372;
    wire _8373;
    wire [63:0] _8377;
    wire [63:0] _8379;
    wire [63:0] _817;
    reg [63:0] _8376;
    wire _8381;
    wire _8382;
    wire [63:0] _8386;
    wire [63:0] _8388;
    wire [63:0] _818;
    reg [63:0] _8385;
    wire _8390;
    wire _8391;
    wire [63:0] _8395;
    wire [63:0] _8397;
    wire [63:0] _819;
    reg [63:0] _8394;
    wire _8399;
    wire _8400;
    wire [63:0] _8404;
    wire [63:0] _8406;
    wire [63:0] _820;
    reg [63:0] _8403;
    wire _8408;
    wire _8409;
    wire [63:0] _8413;
    wire [63:0] _8415;
    wire [63:0] _821;
    reg [63:0] _8412;
    wire _8417;
    wire _8418;
    wire [63:0] _8422;
    wire [63:0] _8424;
    wire [63:0] _822;
    reg [63:0] _8421;
    wire _8426;
    wire _8427;
    wire [63:0] _8431;
    wire [63:0] _8433;
    wire [63:0] _823;
    reg [63:0] _8430;
    wire _8435;
    wire _8436;
    wire [63:0] _8440;
    wire [63:0] _8442;
    wire [63:0] _824;
    reg [63:0] _8439;
    wire _8444;
    wire _8445;
    wire [63:0] _8449;
    wire [63:0] _8451;
    wire [63:0] _825;
    reg [63:0] _8448;
    wire _8453;
    wire _8454;
    wire [63:0] _8458;
    wire [63:0] _8460;
    wire [63:0] _826;
    reg [63:0] _8457;
    wire _8462;
    wire _8463;
    wire [63:0] _8467;
    wire [63:0] _8469;
    wire [63:0] _827;
    reg [63:0] _8466;
    wire _8471;
    wire _8472;
    wire [63:0] _8476;
    wire [63:0] _8478;
    wire [63:0] _828;
    reg [63:0] _8475;
    wire _8480;
    wire _8481;
    wire [63:0] _8485;
    wire [63:0] _8487;
    wire [63:0] _829;
    reg [63:0] _8484;
    wire _8489;
    wire _8490;
    wire [63:0] _8494;
    wire [63:0] _8496;
    wire [63:0] _830;
    reg [63:0] _8493;
    wire _8498;
    wire _8499;
    wire [63:0] _8503;
    wire [63:0] _8505;
    wire [63:0] _831;
    reg [63:0] _8502;
    wire _8507;
    wire _8508;
    wire [63:0] _8512;
    wire [63:0] _8514;
    wire [63:0] _832;
    reg [63:0] _8511;
    wire _8516;
    wire _8517;
    wire [63:0] _8521;
    wire [63:0] _8523;
    wire [63:0] _833;
    reg [63:0] _8520;
    wire _8525;
    wire _8526;
    wire [63:0] _8530;
    wire [63:0] _8532;
    wire [63:0] _834;
    reg [63:0] _8529;
    wire _8534;
    wire _8535;
    wire [63:0] _8539;
    wire [63:0] _8541;
    wire [63:0] _835;
    reg [63:0] _8538;
    wire _8543;
    wire _8544;
    wire [63:0] _8548;
    wire [63:0] _8550;
    wire [63:0] _836;
    reg [63:0] _8547;
    wire _8552;
    wire _8553;
    wire [63:0] _8557;
    wire [63:0] _8559;
    wire [63:0] _837;
    reg [63:0] _8556;
    wire _8561;
    wire _8562;
    wire [63:0] _8566;
    wire [63:0] _8568;
    wire [63:0] _838;
    reg [63:0] _8565;
    wire _8570;
    wire _8571;
    wire [63:0] _8575;
    wire [63:0] _8577;
    wire [63:0] _839;
    reg [63:0] _8574;
    wire _8579;
    wire _8580;
    wire [63:0] _8584;
    wire [63:0] _8586;
    wire [63:0] _840;
    reg [63:0] _8583;
    wire _8588;
    wire _8589;
    wire [63:0] _8593;
    wire [63:0] _8595;
    wire [63:0] _841;
    reg [63:0] _8592;
    wire _8597;
    wire _8598;
    wire [63:0] _8602;
    wire [63:0] _8604;
    wire [63:0] _842;
    reg [63:0] _8601;
    wire _8606;
    wire _8607;
    wire [63:0] _8611;
    wire [63:0] _8613;
    wire [63:0] _843;
    reg [63:0] _8610;
    wire _8615;
    wire _8616;
    wire [63:0] _8620;
    wire [63:0] _8622;
    wire [63:0] _844;
    reg [63:0] _8619;
    wire _8624;
    wire _8625;
    wire [63:0] _8629;
    wire [63:0] _8631;
    wire [63:0] _845;
    reg [63:0] _8628;
    wire _8633;
    wire _8634;
    wire [63:0] _8638;
    wire [63:0] _8640;
    wire [63:0] _846;
    reg [63:0] _8637;
    wire _8642;
    wire _8643;
    wire [63:0] _8647;
    wire [63:0] _8649;
    wire [63:0] _847;
    reg [63:0] _8646;
    wire _8651;
    wire _8652;
    wire [63:0] _8656;
    wire [63:0] _8658;
    wire [63:0] _848;
    reg [63:0] _8655;
    wire _8660;
    wire _8661;
    wire [63:0] _8665;
    wire [63:0] _8667;
    wire [63:0] _849;
    reg [63:0] _8664;
    wire _8669;
    wire _8670;
    wire [63:0] _8674;
    wire [63:0] _8676;
    wire [63:0] _850;
    reg [63:0] _8673;
    wire _8678;
    wire _8679;
    wire [63:0] _8683;
    wire [63:0] _8685;
    wire [63:0] _851;
    reg [63:0] _8682;
    wire _8687;
    wire _8688;
    wire [63:0] _8692;
    wire [63:0] _8694;
    wire [63:0] _852;
    reg [63:0] _8691;
    wire _8696;
    wire _8697;
    wire [63:0] _8701;
    wire [63:0] _8703;
    wire [63:0] _853;
    reg [63:0] _8700;
    wire _8705;
    wire _8706;
    wire [63:0] _8710;
    wire [63:0] _8712;
    wire [63:0] _854;
    reg [63:0] _8709;
    wire _8714;
    wire _8715;
    wire [63:0] _8719;
    wire [63:0] _8721;
    wire [63:0] _855;
    reg [63:0] _8718;
    wire _8723;
    wire _8724;
    wire [63:0] _8728;
    wire [63:0] _8730;
    wire [63:0] _856;
    reg [63:0] _8727;
    wire _8732;
    wire _8733;
    wire [63:0] _8737;
    wire [63:0] _8739;
    wire [63:0] _857;
    reg [63:0] _8736;
    wire _8741;
    wire _8742;
    wire [63:0] _8746;
    wire [63:0] _8748;
    wire [63:0] _858;
    reg [63:0] _8745;
    wire _8750;
    wire _8751;
    wire [63:0] _8755;
    wire [63:0] _8757;
    wire [63:0] _859;
    reg [63:0] _8754;
    wire _8759;
    wire _8760;
    wire [63:0] _8764;
    wire [63:0] _8766;
    wire [63:0] _860;
    reg [63:0] _8763;
    wire _8768;
    wire _8769;
    wire [63:0] _8773;
    wire [63:0] _8775;
    wire [63:0] _861;
    reg [63:0] _8772;
    wire _8777;
    wire _8778;
    wire [63:0] _8782;
    wire [63:0] _8784;
    wire [63:0] _862;
    reg [63:0] _8781;
    wire _8786;
    wire _8787;
    wire [63:0] _8791;
    wire [63:0] _8793;
    wire [63:0] _863;
    reg [63:0] _8790;
    wire _8795;
    wire _8796;
    wire [63:0] _8800;
    wire [63:0] _8802;
    wire [63:0] _864;
    reg [63:0] _8799;
    wire _8804;
    wire _8805;
    wire [63:0] _8809;
    wire [63:0] _8811;
    wire [63:0] _865;
    reg [63:0] _8808;
    wire _8813;
    wire _8814;
    wire [63:0] _8818;
    wire [63:0] _8820;
    wire [63:0] _866;
    reg [63:0] _8817;
    wire _8822;
    wire _8823;
    wire [63:0] _8827;
    wire [63:0] _8829;
    wire [63:0] _867;
    reg [63:0] _8826;
    wire _8831;
    wire _8832;
    wire [63:0] _8836;
    wire [63:0] _8838;
    wire [63:0] _868;
    reg [63:0] _8835;
    wire _8840;
    wire _8841;
    wire [63:0] _8845;
    wire [63:0] _8847;
    wire [63:0] _869;
    reg [63:0] _8844;
    wire _8849;
    wire _8850;
    wire [63:0] _8854;
    wire [63:0] _8856;
    wire [63:0] _870;
    reg [63:0] _8853;
    wire _8858;
    wire _8859;
    wire [63:0] _8863;
    wire [63:0] _8865;
    wire [63:0] _871;
    reg [63:0] _8862;
    wire _8867;
    wire _8868;
    wire [63:0] _8872;
    wire [63:0] _8874;
    wire [63:0] _872;
    reg [63:0] _8871;
    wire _8876;
    wire _8877;
    wire [63:0] _8881;
    wire [63:0] _8883;
    wire [63:0] _873;
    reg [63:0] _8880;
    wire _8885;
    wire _8886;
    wire [63:0] _8890;
    wire [63:0] _8892;
    wire [63:0] _874;
    reg [63:0] _8889;
    wire _8894;
    wire _8895;
    wire [63:0] _8899;
    wire [63:0] _8901;
    wire [63:0] _875;
    reg [63:0] _8898;
    wire _8903;
    wire _8904;
    wire [63:0] _8908;
    wire [63:0] _8910;
    wire [63:0] _876;
    reg [63:0] _8907;
    wire _8912;
    wire _8913;
    wire [63:0] _8917;
    wire [63:0] _8919;
    wire [63:0] _877;
    reg [63:0] _8916;
    wire _8921;
    wire _8922;
    wire [63:0] _8926;
    wire [63:0] _8928;
    wire [63:0] _878;
    reg [63:0] _8925;
    wire _8930;
    wire _8931;
    wire [63:0] _8935;
    wire [63:0] _8937;
    wire [63:0] _879;
    reg [63:0] _8934;
    wire _8939;
    wire _8940;
    wire [63:0] _8944;
    wire [63:0] _8946;
    wire [63:0] _880;
    reg [63:0] _8943;
    wire _8948;
    wire _8949;
    wire [63:0] _8953;
    wire [63:0] _8955;
    wire [63:0] _881;
    reg [63:0] _8952;
    wire _8957;
    wire _8958;
    wire [63:0] _8962;
    wire [63:0] _8964;
    wire [63:0] _882;
    reg [63:0] _8961;
    wire _8966;
    wire _8967;
    wire [63:0] _8971;
    wire [63:0] _8973;
    wire [63:0] _883;
    reg [63:0] _8970;
    wire _8975;
    wire _8976;
    wire [63:0] _8980;
    wire [63:0] _8982;
    wire [63:0] _884;
    reg [63:0] _8979;
    wire _8984;
    wire _8985;
    wire [63:0] _8989;
    wire [63:0] _8991;
    wire [63:0] _885;
    reg [63:0] _8988;
    wire _8993;
    wire _8994;
    wire [63:0] _8998;
    wire [63:0] _9000;
    wire [63:0] _886;
    reg [63:0] _8997;
    wire _9002;
    wire _9003;
    wire [63:0] _9007;
    wire [63:0] _9009;
    wire [63:0] _887;
    reg [63:0] _9006;
    wire _9011;
    wire _9012;
    wire [63:0] _9016;
    wire [63:0] _9018;
    wire [63:0] _888;
    reg [63:0] _9015;
    wire _9020;
    wire _9021;
    wire [63:0] _9025;
    wire [63:0] _9027;
    wire [63:0] _889;
    reg [63:0] _9024;
    wire _9029;
    wire _9030;
    wire [63:0] _9034;
    wire [63:0] _9036;
    wire [63:0] _890;
    reg [63:0] _9033;
    wire _9038;
    wire _9039;
    wire [63:0] _9043;
    wire [63:0] _9045;
    wire [63:0] _891;
    reg [63:0] _9042;
    wire _9047;
    wire _9048;
    wire [63:0] _9052;
    wire [63:0] _9054;
    wire [63:0] _892;
    reg [63:0] _9051;
    wire _9056;
    wire _9057;
    wire [63:0] _9061;
    wire [63:0] _9063;
    wire [63:0] _893;
    reg [63:0] _9060;
    wire _9065;
    wire _9066;
    wire [63:0] _9070;
    wire [63:0] _9072;
    wire [63:0] _894;
    reg [63:0] _9069;
    wire _9074;
    wire _9075;
    wire [63:0] _9079;
    wire [63:0] _9081;
    wire [63:0] _895;
    reg [63:0] _9078;
    wire _9083;
    wire _9084;
    wire [63:0] _9088;
    wire [63:0] _9090;
    wire [63:0] _896;
    reg [63:0] _9087;
    wire _9092;
    wire _9093;
    wire [63:0] _9097;
    wire [63:0] _9099;
    wire [63:0] _897;
    reg [63:0] _9096;
    wire _9101;
    wire _9102;
    wire [63:0] _9106;
    wire [63:0] _9108;
    wire [63:0] _898;
    reg [63:0] _9105;
    wire _9110;
    wire _9111;
    wire [63:0] _9115;
    wire [63:0] _9117;
    wire [63:0] _899;
    reg [63:0] _9114;
    wire _9119;
    wire _9120;
    wire [63:0] _9124;
    wire [63:0] _9126;
    wire [63:0] _900;
    reg [63:0] _9123;
    wire _9128;
    wire _9129;
    wire [63:0] _9133;
    wire [63:0] _9135;
    wire [63:0] _901;
    reg [63:0] _9132;
    wire _9137;
    wire _9138;
    wire [63:0] _9142;
    wire [63:0] _9144;
    wire [63:0] _902;
    reg [63:0] _9141;
    wire _9146;
    wire _9147;
    wire [63:0] _9151;
    wire [63:0] _9153;
    wire [63:0] _903;
    reg [63:0] _9150;
    wire _9155;
    wire _9156;
    wire [63:0] _9160;
    wire [63:0] _9162;
    wire [63:0] _904;
    reg [63:0] _9159;
    wire _9164;
    wire _9165;
    wire [63:0] _9169;
    wire [63:0] _9171;
    wire [63:0] _905;
    reg [63:0] _9168;
    wire _9173;
    wire _9174;
    wire [63:0] _9178;
    wire [63:0] _9180;
    wire [63:0] _906;
    reg [63:0] _9177;
    wire _9182;
    wire _9183;
    wire [63:0] _9187;
    wire [63:0] _9189;
    wire [63:0] _907;
    reg [63:0] _9186;
    wire _9191;
    wire _9192;
    wire [63:0] _9196;
    wire [63:0] _9198;
    wire [63:0] _908;
    reg [63:0] _9195;
    wire _9200;
    wire _9201;
    wire [63:0] _9205;
    wire [63:0] _9207;
    wire [63:0] _909;
    reg [63:0] _9204;
    wire _9209;
    wire _9210;
    wire [63:0] _9214;
    wire [63:0] _9216;
    wire [63:0] _910;
    reg [63:0] _9213;
    wire _9218;
    wire _9219;
    wire [63:0] _9223;
    wire [63:0] _9225;
    wire [63:0] _911;
    reg [63:0] _9222;
    wire _9227;
    wire _9228;
    wire [63:0] _9232;
    wire [63:0] _9234;
    wire [63:0] _912;
    reg [63:0] _9231;
    wire _9236;
    wire _9237;
    wire [63:0] _9241;
    wire [63:0] _9243;
    wire [63:0] _913;
    reg [63:0] _9240;
    wire _9245;
    wire _9246;
    wire [63:0] _9250;
    wire [63:0] _9252;
    wire [63:0] _914;
    reg [63:0] _9249;
    wire _9254;
    wire _9255;
    wire [63:0] _9259;
    wire [63:0] _9261;
    wire [63:0] _915;
    reg [63:0] _9258;
    wire _9263;
    wire _9264;
    wire [63:0] _9268;
    wire [63:0] _9270;
    wire [63:0] _916;
    reg [63:0] _9267;
    wire _9272;
    wire _9273;
    wire [63:0] _9277;
    wire [63:0] _9279;
    wire [63:0] _917;
    reg [63:0] _9276;
    wire _9281;
    wire _9282;
    wire [63:0] _9286;
    wire [63:0] _9288;
    wire [63:0] _918;
    reg [63:0] _9285;
    wire _9290;
    wire _9291;
    wire [63:0] _9295;
    wire [63:0] _9297;
    wire [63:0] _919;
    reg [63:0] _9294;
    wire _9299;
    wire _9300;
    wire [63:0] _9304;
    wire [63:0] _9306;
    wire [63:0] _920;
    reg [63:0] _9303;
    wire _9308;
    wire _9309;
    wire [63:0] _9313;
    wire [63:0] _9315;
    wire [63:0] _921;
    reg [63:0] _9312;
    wire _9317;
    wire _9318;
    wire [63:0] _9322;
    wire [63:0] _9324;
    wire [63:0] _922;
    reg [63:0] _9321;
    wire _9326;
    wire _9327;
    wire [63:0] _9331;
    wire [63:0] _9333;
    wire [63:0] _923;
    reg [63:0] _9330;
    wire _9335;
    wire _9336;
    wire [63:0] _9340;
    wire [63:0] _9342;
    wire [63:0] _924;
    reg [63:0] _9339;
    wire _9344;
    wire _9345;
    wire [63:0] _9349;
    wire [63:0] _9351;
    wire [63:0] _925;
    reg [63:0] _9348;
    wire _9353;
    wire _9354;
    wire [63:0] _9358;
    wire [63:0] _9360;
    wire [63:0] _926;
    reg [63:0] _9357;
    wire _9362;
    wire _9363;
    wire [63:0] _9367;
    wire [63:0] _9369;
    wire [63:0] _927;
    reg [63:0] _9366;
    wire _9371;
    wire _9372;
    wire [63:0] _9376;
    wire [63:0] _9378;
    wire [63:0] _928;
    reg [63:0] _9375;
    wire _9380;
    wire _9381;
    wire [63:0] _9385;
    wire [63:0] _9387;
    wire [63:0] _929;
    reg [63:0] _9384;
    wire _9389;
    wire _9390;
    wire [63:0] _9394;
    wire [63:0] _9396;
    wire [63:0] _930;
    reg [63:0] _9393;
    wire _9398;
    wire _9399;
    wire [63:0] _9403;
    wire [63:0] _9405;
    wire [63:0] _931;
    reg [63:0] _9402;
    wire _9407;
    wire _9408;
    wire [63:0] _9412;
    wire [63:0] _9414;
    wire [63:0] _932;
    reg [63:0] _9411;
    wire _9416;
    wire _9417;
    wire [63:0] _9421;
    wire [63:0] _9423;
    wire [63:0] _933;
    reg [63:0] _9420;
    wire _9425;
    wire _9426;
    wire [63:0] _9430;
    wire [63:0] _9432;
    wire [63:0] _934;
    reg [63:0] _9429;
    wire _9434;
    wire _9435;
    wire [63:0] _9439;
    wire [63:0] _9441;
    wire [63:0] _935;
    reg [63:0] _9438;
    wire _9443;
    wire _9444;
    wire [63:0] _9448;
    wire [63:0] _9450;
    wire [63:0] _936;
    reg [63:0] _9447;
    wire _9452;
    wire _9453;
    wire [63:0] _9457;
    wire [63:0] _9459;
    wire [63:0] _937;
    reg [63:0] _9456;
    wire _9461;
    wire _9462;
    wire [63:0] _9466;
    wire [63:0] _9468;
    wire [63:0] _938;
    reg [63:0] _9465;
    wire _9470;
    wire _9471;
    wire [63:0] _9475;
    wire [63:0] _9477;
    wire [63:0] _939;
    reg [63:0] _9474;
    wire _9479;
    wire _9480;
    wire [63:0] _9484;
    wire [63:0] _9486;
    wire [63:0] _940;
    reg [63:0] _9483;
    wire _9488;
    wire _9489;
    wire [63:0] _9493;
    wire [63:0] _9495;
    wire [63:0] _941;
    reg [63:0] _9492;
    wire _9497;
    wire _9498;
    wire [63:0] _9502;
    wire [63:0] _9504;
    wire [63:0] _942;
    reg [63:0] _9501;
    wire _9506;
    wire _9507;
    wire [63:0] _9511;
    wire [63:0] _9513;
    wire [63:0] _943;
    reg [63:0] _9510;
    wire _9515;
    wire _9516;
    wire [63:0] _9520;
    wire [63:0] _9522;
    wire [63:0] _944;
    reg [63:0] _9519;
    wire _9524;
    wire _9525;
    wire [63:0] _9529;
    wire [63:0] _9531;
    wire [63:0] _945;
    reg [63:0] _9528;
    wire _9533;
    wire _9534;
    wire [63:0] _9538;
    wire [63:0] _9540;
    wire [63:0] _946;
    reg [63:0] _9537;
    wire _9542;
    wire _9543;
    wire [63:0] _9547;
    wire [63:0] _9549;
    wire [63:0] _947;
    reg [63:0] _9546;
    wire _9551;
    wire _9552;
    wire [63:0] _9556;
    wire [63:0] _9558;
    wire [63:0] _948;
    reg [63:0] _9555;
    wire _9560;
    wire _9561;
    wire [63:0] _9565;
    wire [63:0] _9567;
    wire [63:0] _949;
    reg [63:0] _9564;
    wire _9569;
    wire _9570;
    wire [63:0] _9574;
    wire [63:0] _9576;
    wire [63:0] _950;
    reg [63:0] _9573;
    wire _9578;
    wire _9579;
    wire [63:0] _9583;
    wire [63:0] _9585;
    wire [63:0] _951;
    reg [63:0] _9582;
    wire _9587;
    wire _9588;
    wire [63:0] _9592;
    wire [63:0] _9594;
    wire [63:0] _952;
    reg [63:0] _9591;
    wire _9596;
    wire _9597;
    wire [63:0] _9601;
    wire [63:0] _9603;
    wire [63:0] _953;
    reg [63:0] _9600;
    wire _9605;
    wire _9606;
    wire [63:0] _9610;
    wire [63:0] _9612;
    wire [63:0] _954;
    reg [63:0] _9609;
    wire _9614;
    wire _9615;
    wire [63:0] _9619;
    wire [63:0] _9621;
    wire [63:0] _955;
    reg [63:0] _9618;
    wire _9623;
    wire _9624;
    wire [63:0] _9628;
    wire [63:0] _9630;
    wire [63:0] _956;
    reg [63:0] _9627;
    wire _9632;
    wire _9633;
    wire [63:0] _9637;
    wire [63:0] _9639;
    wire [63:0] _957;
    reg [63:0] _9636;
    wire _9641;
    wire _9642;
    wire [63:0] _9646;
    wire [63:0] _9648;
    wire [63:0] _958;
    reg [63:0] _9645;
    wire _9650;
    wire _9651;
    wire [63:0] _9655;
    wire [63:0] _9657;
    wire [63:0] _959;
    reg [63:0] _9654;
    wire _9659;
    wire _9660;
    wire [63:0] _9664;
    wire [63:0] _9666;
    wire [63:0] _960;
    reg [63:0] _9663;
    wire _9668;
    wire _9669;
    wire [63:0] _9673;
    wire [63:0] _9675;
    wire [63:0] _961;
    reg [63:0] _9672;
    wire _9677;
    wire _9678;
    wire [63:0] _9682;
    wire [63:0] _9684;
    wire [63:0] _962;
    reg [63:0] _9681;
    wire _9686;
    wire _9687;
    wire [63:0] _9691;
    wire [63:0] _9693;
    wire [63:0] _963;
    reg [63:0] _9690;
    wire _9695;
    wire _9696;
    wire [63:0] _9700;
    wire [63:0] _9702;
    wire [63:0] _964;
    reg [63:0] _9699;
    wire _9704;
    wire _9705;
    wire [63:0] _9709;
    wire [63:0] _9711;
    wire [63:0] _965;
    reg [63:0] _9708;
    wire _9713;
    wire _9714;
    wire [63:0] _9718;
    wire [63:0] _9720;
    wire [63:0] _966;
    reg [63:0] _9717;
    wire _9722;
    wire _9723;
    wire [63:0] _9727;
    wire [63:0] _9729;
    wire [63:0] _967;
    reg [63:0] _9726;
    wire _9731;
    wire _9732;
    wire [63:0] _9736;
    wire [63:0] _9738;
    wire [63:0] _968;
    reg [63:0] _9735;
    wire _9740;
    wire _9741;
    wire [63:0] _9745;
    wire [63:0] _9747;
    wire [63:0] _969;
    reg [63:0] _9744;
    wire _9749;
    wire _9750;
    wire [63:0] _9754;
    wire [63:0] _9756;
    wire [63:0] _970;
    reg [63:0] _9753;
    wire _9758;
    wire _9759;
    wire [63:0] _9763;
    wire [63:0] _9765;
    wire [63:0] _971;
    reg [63:0] _9762;
    wire _9767;
    wire _9768;
    wire [63:0] _9772;
    wire [63:0] _9774;
    wire [63:0] _972;
    reg [63:0] _9771;
    wire _9776;
    wire _9777;
    wire [63:0] _9781;
    wire [63:0] _9783;
    wire [63:0] _973;
    reg [63:0] _9780;
    wire _9785;
    wire _9786;
    wire [63:0] _9790;
    wire [63:0] _9792;
    wire [63:0] _974;
    reg [63:0] _9789;
    wire _9794;
    wire _9795;
    wire [63:0] _9799;
    wire [63:0] _9801;
    wire [63:0] _975;
    reg [63:0] _9798;
    wire _9803;
    wire _9804;
    wire [63:0] _9808;
    wire [63:0] _9810;
    wire [63:0] _976;
    reg [63:0] _9807;
    wire _9812;
    wire _9813;
    wire [63:0] _9817;
    wire [63:0] _9819;
    wire [63:0] _977;
    reg [63:0] _9816;
    wire _9821;
    wire _9822;
    wire [63:0] _9826;
    wire [63:0] _9828;
    wire [63:0] _978;
    reg [63:0] _9825;
    wire _9830;
    wire _9831;
    wire [63:0] _9835;
    wire [63:0] _9837;
    wire [63:0] _979;
    reg [63:0] _9834;
    wire _9839;
    wire _9840;
    wire [63:0] _9844;
    wire [63:0] _9846;
    wire [63:0] _980;
    reg [63:0] _9843;
    wire _9848;
    wire _9849;
    wire [63:0] _9853;
    wire [63:0] _9855;
    wire [63:0] _981;
    reg [63:0] _9852;
    wire _9857;
    wire _9858;
    wire [63:0] _9862;
    wire [63:0] _9864;
    wire [63:0] _982;
    reg [63:0] _9861;
    wire _9866;
    wire _9867;
    wire [63:0] _9871;
    wire [63:0] _9873;
    wire [63:0] _983;
    reg [63:0] _9870;
    wire _9875;
    wire _9876;
    wire [63:0] _9880;
    wire [63:0] _9882;
    wire [63:0] _984;
    reg [63:0] _9879;
    wire _9884;
    wire _9885;
    wire [63:0] _9889;
    wire [63:0] _9891;
    wire [63:0] _985;
    reg [63:0] _9888;
    wire _9893;
    wire _9894;
    wire [63:0] _9898;
    wire [63:0] _9900;
    wire [63:0] _986;
    reg [63:0] _9897;
    wire _9902;
    wire _9903;
    wire [63:0] _9907;
    wire [63:0] _9909;
    wire [63:0] _987;
    reg [63:0] _9906;
    wire _9911;
    wire _9912;
    wire [63:0] _9916;
    wire [63:0] _9918;
    wire [63:0] _988;
    reg [63:0] _9915;
    wire _9920;
    wire _9921;
    wire [63:0] _9925;
    wire [63:0] _9927;
    wire [63:0] _989;
    reg [63:0] _9924;
    wire _9929;
    wire _9930;
    wire [63:0] _9934;
    wire [63:0] _9936;
    wire [63:0] _990;
    reg [63:0] _9933;
    wire _9938;
    wire _9939;
    wire [63:0] _9943;
    wire [63:0] _9945;
    wire [63:0] _991;
    reg [63:0] _9942;
    wire _9947;
    wire _9948;
    wire [63:0] _9952;
    wire [63:0] _9954;
    wire [63:0] _992;
    reg [63:0] _9951;
    wire _9956;
    wire _9957;
    wire [63:0] _9961;
    wire [63:0] _9963;
    wire [63:0] _993;
    reg [63:0] _9960;
    wire _9965;
    wire _9966;
    wire [63:0] _9970;
    wire [63:0] _9972;
    wire [63:0] _994;
    reg [63:0] _9969;
    wire _9974;
    wire _9975;
    wire [63:0] _9979;
    wire [63:0] _9981;
    wire [63:0] _995;
    reg [63:0] _9978;
    wire _9983;
    wire _9984;
    wire [63:0] _9988;
    wire [63:0] _9990;
    wire [63:0] _996;
    reg [63:0] _9987;
    wire _9992;
    wire _9993;
    wire [63:0] _9997;
    wire [63:0] _9999;
    wire [63:0] _997;
    reg [63:0] _9996;
    wire _10001;
    wire _10002;
    wire [63:0] _10006;
    wire [63:0] _10008;
    wire [63:0] _998;
    reg [63:0] _10005;
    wire _10010;
    wire _10011;
    wire [63:0] _10015;
    wire [63:0] _10017;
    wire [63:0] _999;
    reg [63:0] _10014;
    wire _10019;
    wire _10020;
    wire [63:0] _10024;
    wire [63:0] _10026;
    wire [63:0] _1000;
    reg [63:0] _10023;
    wire _10028;
    wire _10029;
    wire [63:0] _10033;
    wire [63:0] _10035;
    wire [63:0] _1001;
    reg [63:0] _10032;
    wire _10037;
    wire _10038;
    wire [63:0] _10042;
    wire [63:0] _10044;
    wire [63:0] _1002;
    reg [63:0] _10041;
    wire _10046;
    wire _10047;
    wire [63:0] _10051;
    wire [63:0] _10053;
    wire [63:0] _1003;
    reg [63:0] _10050;
    wire _10055;
    wire _10056;
    wire [63:0] _10060;
    wire [63:0] _10062;
    wire [63:0] _1004;
    reg [63:0] _10059;
    wire _10064;
    wire _10065;
    wire [63:0] _10069;
    wire [63:0] _10071;
    wire [63:0] _1005;
    reg [63:0] _10068;
    wire _10073;
    wire _10074;
    wire [63:0] _10078;
    wire [63:0] _10080;
    wire [63:0] _1006;
    reg [63:0] _10077;
    wire _10082;
    wire _10083;
    wire [63:0] _10087;
    wire [63:0] _10089;
    wire [63:0] _1007;
    reg [63:0] _10086;
    wire _10091;
    wire _10092;
    wire [63:0] _10096;
    wire [63:0] _10098;
    wire [63:0] _1008;
    reg [63:0] _10095;
    wire _10100;
    wire _10101;
    wire [63:0] _10105;
    wire [63:0] _10107;
    wire [63:0] _1009;
    reg [63:0] _10104;
    wire _10109;
    wire _10110;
    wire [63:0] _10114;
    wire [63:0] _10116;
    wire [63:0] _1010;
    reg [63:0] _10113;
    wire _10118;
    wire _10119;
    wire [63:0] _10123;
    wire [63:0] _10125;
    wire [63:0] _1011;
    reg [63:0] _10122;
    wire _10127;
    wire _10128;
    wire [63:0] _10132;
    wire [63:0] _10134;
    wire [63:0] _1012;
    reg [63:0] _10131;
    wire _10136;
    wire _10137;
    wire [63:0] _10141;
    wire [63:0] _10143;
    wire [63:0] _1013;
    reg [63:0] _10140;
    wire _10145;
    wire _10146;
    wire [63:0] _10150;
    wire [63:0] _10152;
    wire [63:0] _1014;
    reg [63:0] _10149;
    wire _10154;
    wire _10155;
    wire [63:0] _10159;
    wire [63:0] _10161;
    wire [63:0] _1015;
    reg [63:0] _10158;
    wire _10163;
    wire _10164;
    wire [63:0] _10168;
    wire [63:0] _10170;
    wire [63:0] _1016;
    reg [63:0] _10167;
    wire _10172;
    wire _10173;
    wire [63:0] _10177;
    wire [63:0] _10179;
    wire [63:0] _1017;
    reg [63:0] _10176;
    wire _10181;
    wire _10182;
    wire [63:0] _10186;
    wire [63:0] _10188;
    wire [63:0] _1018;
    reg [63:0] _10185;
    wire _10190;
    wire _10191;
    wire [63:0] _10195;
    wire [63:0] _10197;
    wire [63:0] _1019;
    reg [63:0] _10194;
    wire _10199;
    wire _10200;
    wire [63:0] _10204;
    wire [63:0] _10206;
    wire [63:0] _1020;
    reg [63:0] _10203;
    wire _10208;
    wire _10209;
    wire [63:0] _10213;
    wire [63:0] _10215;
    wire [63:0] _1021;
    reg [63:0] _10212;
    wire _10217;
    wire _10218;
    wire [63:0] _10222;
    wire [63:0] _10224;
    wire [63:0] _1022;
    reg [63:0] _10221;
    wire _10226;
    wire _10227;
    wire [63:0] _10231;
    wire [63:0] _10233;
    wire [63:0] _1023;
    reg [63:0] _10230;
    wire _10235;
    wire _10236;
    wire [63:0] _10240;
    wire [63:0] _10242;
    wire [63:0] _1024;
    reg [63:0] _10239;
    wire _10244;
    wire _10245;
    wire [63:0] _10249;
    wire [63:0] _10251;
    wire [63:0] _1025;
    reg [63:0] _10248;
    wire _10253;
    wire _10254;
    wire [63:0] _10258;
    wire [63:0] _10260;
    wire [63:0] _1026;
    reg [63:0] _10257;
    wire _10262;
    wire _10263;
    wire [63:0] _10267;
    wire [63:0] _10269;
    wire [63:0] _1027;
    reg [63:0] _10266;
    wire [63:0] _1029;
    wire _10271;
    wire _10272;
    wire [63:0] _10276;
    wire [63:0] _10278;
    wire [63:0] _1030;
    reg [63:0] _10275;
    reg [63:0] _10295;
    wire _10297;
    wire _10298;
    wire [63:0] _10301;
    wire [63:0] _10303;
    wire [127:0] _10313;
    wire [63:0] _10314;
    wire _10315;
    wire _10294;
    wire _10316;
    wire [63:0] _10322;
    wire [63:0] _1031;
    reg [63:0] _1056;
    wire _10324;
    wire [1:0] _1051;
    wire [1:0] _10323;
    wire [8:0] _10363;
    wire [8:0] _10359;
    wire [8:0] _10355;
    wire _10353;
    wire [8:0] _10357;
    wire [8:0] _10337;
    wire [8:0] _10335;
    wire [8:0] _10332;
    wire _10333;
    wire [8:0] _10338;
    wire [8:0] _10328;
    wire _10326;
    wire [8:0] _10330;
    wire _10325;
    wire [8:0] _10339;
    wire [8:0] _1034;
    reg [8:0] _10291;
    wire _10292;
    wire vdd;
    wire _1036;
    wire _1038;
    wire [8:0] _10343;
    wire [8:0] _10341;
    wire [8:0] _10344;
    wire [8:0] _1039;
    reg [8:0] _1062;
    wire [8:0] _10349;
    wire [8:0] _10347;
    wire _10345;
    wire [8:0] _10350;
    wire [8:0] _1040;
    reg [8:0] _10286;
    wire _10287;
    wire _10288;
    wire _10293;
    wire _10351;
    wire _10352;
    wire [8:0] _10360;
    wire [8:0] _1041;
    reg [8:0] _10283;
    wire _10364;
    wire [1:0] _10279;
    wire _10280;
    wire _10365;
    wire _10366;
    wire [1:0] _10367;
    wire _1043;
    wire _1045;
    wire _1059;
    wire _10361;
    wire [1:0] _10368;
    wire _1047;
    wire [1:0] _10369;
    wire [1:0] _1048;
    reg [1:0] _1053;
    wire _1058;
    assign _1055 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign _10319 = _1047 ? _1055 : _1056;
    assign _10317 = _1059 & _1043;
    assign _10321 = _10317 ? _1055 : _10319;
    assign _10311 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    assign _10309 = _10304 - _10305;
    assign _10308 = _10305 - _10304;
    always @* begin
        case (_10291)
        0:
            _10305 <= _5667;
        1:
            _10305 <= _5658;
        2:
            _10305 <= _5649;
        3:
            _10305 <= _5640;
        4:
            _10305 <= _5631;
        5:
            _10305 <= _5622;
        6:
            _10305 <= _5613;
        7:
            _10305 <= _5604;
        8:
            _10305 <= _5595;
        9:
            _10305 <= _5586;
        10:
            _10305 <= _5577;
        11:
            _10305 <= _5568;
        12:
            _10305 <= _5559;
        13:
            _10305 <= _5550;
        14:
            _10305 <= _5541;
        15:
            _10305 <= _5532;
        16:
            _10305 <= _5523;
        17:
            _10305 <= _5514;
        18:
            _10305 <= _5505;
        19:
            _10305 <= _5496;
        20:
            _10305 <= _5487;
        21:
            _10305 <= _5478;
        22:
            _10305 <= _5469;
        23:
            _10305 <= _5460;
        24:
            _10305 <= _5451;
        25:
            _10305 <= _5442;
        26:
            _10305 <= _5433;
        27:
            _10305 <= _5424;
        28:
            _10305 <= _5415;
        29:
            _10305 <= _5406;
        30:
            _10305 <= _5397;
        31:
            _10305 <= _5388;
        32:
            _10305 <= _5379;
        33:
            _10305 <= _5370;
        34:
            _10305 <= _5361;
        35:
            _10305 <= _5352;
        36:
            _10305 <= _5343;
        37:
            _10305 <= _5334;
        38:
            _10305 <= _5325;
        39:
            _10305 <= _5316;
        40:
            _10305 <= _5307;
        41:
            _10305 <= _5298;
        42:
            _10305 <= _5289;
        43:
            _10305 <= _5280;
        44:
            _10305 <= _5271;
        45:
            _10305 <= _5262;
        46:
            _10305 <= _5253;
        47:
            _10305 <= _5244;
        48:
            _10305 <= _5235;
        49:
            _10305 <= _5226;
        50:
            _10305 <= _5217;
        51:
            _10305 <= _5208;
        52:
            _10305 <= _5199;
        53:
            _10305 <= _5190;
        54:
            _10305 <= _5181;
        55:
            _10305 <= _5172;
        56:
            _10305 <= _5163;
        57:
            _10305 <= _5154;
        58:
            _10305 <= _5145;
        59:
            _10305 <= _5136;
        60:
            _10305 <= _5127;
        61:
            _10305 <= _5118;
        62:
            _10305 <= _5109;
        63:
            _10305 <= _5100;
        64:
            _10305 <= _5091;
        65:
            _10305 <= _5082;
        66:
            _10305 <= _5073;
        67:
            _10305 <= _5064;
        68:
            _10305 <= _5055;
        69:
            _10305 <= _5046;
        70:
            _10305 <= _5037;
        71:
            _10305 <= _5028;
        72:
            _10305 <= _5019;
        73:
            _10305 <= _5010;
        74:
            _10305 <= _5001;
        75:
            _10305 <= _4992;
        76:
            _10305 <= _4983;
        77:
            _10305 <= _4974;
        78:
            _10305 <= _4965;
        79:
            _10305 <= _4956;
        80:
            _10305 <= _4947;
        81:
            _10305 <= _4938;
        82:
            _10305 <= _4929;
        83:
            _10305 <= _4920;
        84:
            _10305 <= _4911;
        85:
            _10305 <= _4902;
        86:
            _10305 <= _4893;
        87:
            _10305 <= _4884;
        88:
            _10305 <= _4875;
        89:
            _10305 <= _4866;
        90:
            _10305 <= _4857;
        91:
            _10305 <= _4848;
        92:
            _10305 <= _4839;
        93:
            _10305 <= _4830;
        94:
            _10305 <= _4821;
        95:
            _10305 <= _4812;
        96:
            _10305 <= _4803;
        97:
            _10305 <= _4794;
        98:
            _10305 <= _4785;
        99:
            _10305 <= _4776;
        100:
            _10305 <= _4767;
        101:
            _10305 <= _4758;
        102:
            _10305 <= _4749;
        103:
            _10305 <= _4740;
        104:
            _10305 <= _4731;
        105:
            _10305 <= _4722;
        106:
            _10305 <= _4713;
        107:
            _10305 <= _4704;
        108:
            _10305 <= _4695;
        109:
            _10305 <= _4686;
        110:
            _10305 <= _4677;
        111:
            _10305 <= _4668;
        112:
            _10305 <= _4659;
        113:
            _10305 <= _4650;
        114:
            _10305 <= _4641;
        115:
            _10305 <= _4632;
        116:
            _10305 <= _4623;
        117:
            _10305 <= _4614;
        118:
            _10305 <= _4605;
        119:
            _10305 <= _4596;
        120:
            _10305 <= _4587;
        121:
            _10305 <= _4578;
        122:
            _10305 <= _4569;
        123:
            _10305 <= _4560;
        124:
            _10305 <= _4551;
        125:
            _10305 <= _4542;
        126:
            _10305 <= _4533;
        127:
            _10305 <= _4524;
        128:
            _10305 <= _4515;
        129:
            _10305 <= _4506;
        130:
            _10305 <= _4497;
        131:
            _10305 <= _4488;
        132:
            _10305 <= _4479;
        133:
            _10305 <= _4470;
        134:
            _10305 <= _4461;
        135:
            _10305 <= _4452;
        136:
            _10305 <= _4443;
        137:
            _10305 <= _4434;
        138:
            _10305 <= _4425;
        139:
            _10305 <= _4416;
        140:
            _10305 <= _4407;
        141:
            _10305 <= _4398;
        142:
            _10305 <= _4389;
        143:
            _10305 <= _4380;
        144:
            _10305 <= _4371;
        145:
            _10305 <= _4362;
        146:
            _10305 <= _4353;
        147:
            _10305 <= _4344;
        148:
            _10305 <= _4335;
        149:
            _10305 <= _4326;
        150:
            _10305 <= _4317;
        151:
            _10305 <= _4308;
        152:
            _10305 <= _4299;
        153:
            _10305 <= _4290;
        154:
            _10305 <= _4281;
        155:
            _10305 <= _4272;
        156:
            _10305 <= _4263;
        157:
            _10305 <= _4254;
        158:
            _10305 <= _4245;
        159:
            _10305 <= _4236;
        160:
            _10305 <= _4227;
        161:
            _10305 <= _4218;
        162:
            _10305 <= _4209;
        163:
            _10305 <= _4200;
        164:
            _10305 <= _4191;
        165:
            _10305 <= _4182;
        166:
            _10305 <= _4173;
        167:
            _10305 <= _4164;
        168:
            _10305 <= _4155;
        169:
            _10305 <= _4146;
        170:
            _10305 <= _4137;
        171:
            _10305 <= _4128;
        172:
            _10305 <= _4119;
        173:
            _10305 <= _4110;
        174:
            _10305 <= _4101;
        175:
            _10305 <= _4092;
        176:
            _10305 <= _4083;
        177:
            _10305 <= _4074;
        178:
            _10305 <= _4065;
        179:
            _10305 <= _4056;
        180:
            _10305 <= _4047;
        181:
            _10305 <= _4038;
        182:
            _10305 <= _4029;
        183:
            _10305 <= _4020;
        184:
            _10305 <= _4011;
        185:
            _10305 <= _4002;
        186:
            _10305 <= _3993;
        187:
            _10305 <= _3984;
        188:
            _10305 <= _3975;
        189:
            _10305 <= _3966;
        190:
            _10305 <= _3957;
        191:
            _10305 <= _3948;
        192:
            _10305 <= _3939;
        193:
            _10305 <= _3930;
        194:
            _10305 <= _3921;
        195:
            _10305 <= _3912;
        196:
            _10305 <= _3903;
        197:
            _10305 <= _3894;
        198:
            _10305 <= _3885;
        199:
            _10305 <= _3876;
        200:
            _10305 <= _3867;
        201:
            _10305 <= _3858;
        202:
            _10305 <= _3849;
        203:
            _10305 <= _3840;
        204:
            _10305 <= _3831;
        205:
            _10305 <= _3822;
        206:
            _10305 <= _3813;
        207:
            _10305 <= _3804;
        208:
            _10305 <= _3795;
        209:
            _10305 <= _3786;
        210:
            _10305 <= _3777;
        211:
            _10305 <= _3768;
        212:
            _10305 <= _3759;
        213:
            _10305 <= _3750;
        214:
            _10305 <= _3741;
        215:
            _10305 <= _3732;
        216:
            _10305 <= _3723;
        217:
            _10305 <= _3714;
        218:
            _10305 <= _3705;
        219:
            _10305 <= _3696;
        220:
            _10305 <= _3687;
        221:
            _10305 <= _3678;
        222:
            _10305 <= _3669;
        223:
            _10305 <= _3660;
        224:
            _10305 <= _3651;
        225:
            _10305 <= _3642;
        226:
            _10305 <= _3633;
        227:
            _10305 <= _3624;
        228:
            _10305 <= _3615;
        229:
            _10305 <= _3606;
        230:
            _10305 <= _3597;
        231:
            _10305 <= _3588;
        232:
            _10305 <= _3579;
        233:
            _10305 <= _3570;
        234:
            _10305 <= _3561;
        235:
            _10305 <= _3552;
        236:
            _10305 <= _3543;
        237:
            _10305 <= _3534;
        238:
            _10305 <= _3525;
        239:
            _10305 <= _3516;
        240:
            _10305 <= _3507;
        241:
            _10305 <= _3498;
        242:
            _10305 <= _3489;
        243:
            _10305 <= _3480;
        244:
            _10305 <= _3471;
        245:
            _10305 <= _3462;
        246:
            _10305 <= _3453;
        247:
            _10305 <= _3444;
        248:
            _10305 <= _3435;
        249:
            _10305 <= _3426;
        250:
            _10305 <= _3417;
        251:
            _10305 <= _3408;
        252:
            _10305 <= _3399;
        253:
            _10305 <= _3390;
        254:
            _10305 <= _3381;
        255:
            _10305 <= _3372;
        256:
            _10305 <= _3363;
        257:
            _10305 <= _3354;
        258:
            _10305 <= _3345;
        259:
            _10305 <= _3336;
        260:
            _10305 <= _3327;
        261:
            _10305 <= _3318;
        262:
            _10305 <= _3309;
        263:
            _10305 <= _3300;
        264:
            _10305 <= _3291;
        265:
            _10305 <= _3282;
        266:
            _10305 <= _3273;
        267:
            _10305 <= _3264;
        268:
            _10305 <= _3255;
        269:
            _10305 <= _3246;
        270:
            _10305 <= _3237;
        271:
            _10305 <= _3228;
        272:
            _10305 <= _3219;
        273:
            _10305 <= _3210;
        274:
            _10305 <= _3201;
        275:
            _10305 <= _3192;
        276:
            _10305 <= _3183;
        277:
            _10305 <= _3174;
        278:
            _10305 <= _3165;
        279:
            _10305 <= _3156;
        280:
            _10305 <= _3147;
        281:
            _10305 <= _3138;
        282:
            _10305 <= _3129;
        283:
            _10305 <= _3120;
        284:
            _10305 <= _3111;
        285:
            _10305 <= _3102;
        286:
            _10305 <= _3093;
        287:
            _10305 <= _3084;
        288:
            _10305 <= _3075;
        289:
            _10305 <= _3066;
        290:
            _10305 <= _3057;
        291:
            _10305 <= _3048;
        292:
            _10305 <= _3039;
        293:
            _10305 <= _3030;
        294:
            _10305 <= _3021;
        295:
            _10305 <= _3012;
        296:
            _10305 <= _3003;
        297:
            _10305 <= _2994;
        298:
            _10305 <= _2985;
        299:
            _10305 <= _2976;
        300:
            _10305 <= _2967;
        301:
            _10305 <= _2958;
        302:
            _10305 <= _2949;
        303:
            _10305 <= _2940;
        304:
            _10305 <= _2931;
        305:
            _10305 <= _2922;
        306:
            _10305 <= _2913;
        307:
            _10305 <= _2904;
        308:
            _10305 <= _2895;
        309:
            _10305 <= _2886;
        310:
            _10305 <= _2877;
        311:
            _10305 <= _2868;
        312:
            _10305 <= _2859;
        313:
            _10305 <= _2850;
        314:
            _10305 <= _2841;
        315:
            _10305 <= _2832;
        316:
            _10305 <= _2823;
        317:
            _10305 <= _2814;
        318:
            _10305 <= _2805;
        319:
            _10305 <= _2796;
        320:
            _10305 <= _2787;
        321:
            _10305 <= _2778;
        322:
            _10305 <= _2769;
        323:
            _10305 <= _2760;
        324:
            _10305 <= _2751;
        325:
            _10305 <= _2742;
        326:
            _10305 <= _2733;
        327:
            _10305 <= _2724;
        328:
            _10305 <= _2715;
        329:
            _10305 <= _2706;
        330:
            _10305 <= _2697;
        331:
            _10305 <= _2688;
        332:
            _10305 <= _2679;
        333:
            _10305 <= _2670;
        334:
            _10305 <= _2661;
        335:
            _10305 <= _2652;
        336:
            _10305 <= _2643;
        337:
            _10305 <= _2634;
        338:
            _10305 <= _2625;
        339:
            _10305 <= _2616;
        340:
            _10305 <= _2607;
        341:
            _10305 <= _2598;
        342:
            _10305 <= _2589;
        343:
            _10305 <= _2580;
        344:
            _10305 <= _2571;
        345:
            _10305 <= _2562;
        346:
            _10305 <= _2553;
        347:
            _10305 <= _2544;
        348:
            _10305 <= _2535;
        349:
            _10305 <= _2526;
        350:
            _10305 <= _2517;
        351:
            _10305 <= _2508;
        352:
            _10305 <= _2499;
        353:
            _10305 <= _2490;
        354:
            _10305 <= _2481;
        355:
            _10305 <= _2472;
        356:
            _10305 <= _2463;
        357:
            _10305 <= _2454;
        358:
            _10305 <= _2445;
        359:
            _10305 <= _2436;
        360:
            _10305 <= _2427;
        361:
            _10305 <= _2418;
        362:
            _10305 <= _2409;
        363:
            _10305 <= _2400;
        364:
            _10305 <= _2391;
        365:
            _10305 <= _2382;
        366:
            _10305 <= _2373;
        367:
            _10305 <= _2364;
        368:
            _10305 <= _2355;
        369:
            _10305 <= _2346;
        370:
            _10305 <= _2337;
        371:
            _10305 <= _2328;
        372:
            _10305 <= _2319;
        373:
            _10305 <= _2310;
        374:
            _10305 <= _2301;
        375:
            _10305 <= _2292;
        376:
            _10305 <= _2283;
        377:
            _10305 <= _2274;
        378:
            _10305 <= _2265;
        379:
            _10305 <= _2256;
        380:
            _10305 <= _2247;
        381:
            _10305 <= _2238;
        382:
            _10305 <= _2229;
        383:
            _10305 <= _2220;
        384:
            _10305 <= _2211;
        385:
            _10305 <= _2202;
        386:
            _10305 <= _2193;
        387:
            _10305 <= _2184;
        388:
            _10305 <= _2175;
        389:
            _10305 <= _2166;
        390:
            _10305 <= _2157;
        391:
            _10305 <= _2148;
        392:
            _10305 <= _2139;
        393:
            _10305 <= _2130;
        394:
            _10305 <= _2121;
        395:
            _10305 <= _2112;
        396:
            _10305 <= _2103;
        397:
            _10305 <= _2094;
        398:
            _10305 <= _2085;
        399:
            _10305 <= _2076;
        400:
            _10305 <= _2067;
        401:
            _10305 <= _2058;
        402:
            _10305 <= _2049;
        403:
            _10305 <= _2040;
        404:
            _10305 <= _2031;
        405:
            _10305 <= _2022;
        406:
            _10305 <= _2013;
        407:
            _10305 <= _2004;
        408:
            _10305 <= _1995;
        409:
            _10305 <= _1986;
        410:
            _10305 <= _1977;
        411:
            _10305 <= _1968;
        412:
            _10305 <= _1959;
        413:
            _10305 <= _1950;
        414:
            _10305 <= _1941;
        415:
            _10305 <= _1932;
        416:
            _10305 <= _1923;
        417:
            _10305 <= _1914;
        418:
            _10305 <= _1905;
        419:
            _10305 <= _1896;
        420:
            _10305 <= _1887;
        421:
            _10305 <= _1878;
        422:
            _10305 <= _1869;
        423:
            _10305 <= _1860;
        424:
            _10305 <= _1851;
        425:
            _10305 <= _1842;
        426:
            _10305 <= _1833;
        427:
            _10305 <= _1824;
        428:
            _10305 <= _1815;
        429:
            _10305 <= _1806;
        430:
            _10305 <= _1797;
        431:
            _10305 <= _1788;
        432:
            _10305 <= _1779;
        433:
            _10305 <= _1770;
        434:
            _10305 <= _1761;
        435:
            _10305 <= _1752;
        436:
            _10305 <= _1743;
        437:
            _10305 <= _1734;
        438:
            _10305 <= _1725;
        439:
            _10305 <= _1716;
        440:
            _10305 <= _1707;
        441:
            _10305 <= _1698;
        442:
            _10305 <= _1689;
        443:
            _10305 <= _1680;
        444:
            _10305 <= _1671;
        445:
            _10305 <= _1662;
        446:
            _10305 <= _1653;
        447:
            _10305 <= _1644;
        448:
            _10305 <= _1635;
        449:
            _10305 <= _1626;
        450:
            _10305 <= _1617;
        451:
            _10305 <= _1608;
        452:
            _10305 <= _1599;
        453:
            _10305 <= _1590;
        454:
            _10305 <= _1581;
        455:
            _10305 <= _1572;
        456:
            _10305 <= _1563;
        457:
            _10305 <= _1554;
        458:
            _10305 <= _1545;
        459:
            _10305 <= _1536;
        460:
            _10305 <= _1527;
        461:
            _10305 <= _1518;
        462:
            _10305 <= _1509;
        463:
            _10305 <= _1500;
        464:
            _10305 <= _1491;
        465:
            _10305 <= _1482;
        466:
            _10305 <= _1473;
        467:
            _10305 <= _1464;
        468:
            _10305 <= _1455;
        469:
            _10305 <= _1446;
        470:
            _10305 <= _1437;
        471:
            _10305 <= _1428;
        472:
            _10305 <= _1419;
        473:
            _10305 <= _1410;
        474:
            _10305 <= _1401;
        475:
            _10305 <= _1392;
        476:
            _10305 <= _1383;
        477:
            _10305 <= _1374;
        478:
            _10305 <= _1365;
        479:
            _10305 <= _1356;
        480:
            _10305 <= _1347;
        481:
            _10305 <= _1338;
        482:
            _10305 <= _1329;
        483:
            _10305 <= _1320;
        484:
            _10305 <= _1311;
        485:
            _10305 <= _1302;
        486:
            _10305 <= _1293;
        487:
            _10305 <= _1284;
        488:
            _10305 <= _1275;
        489:
            _10305 <= _1266;
        490:
            _10305 <= _1257;
        491:
            _10305 <= _1248;
        492:
            _10305 <= _1239;
        493:
            _10305 <= _1230;
        494:
            _10305 <= _1221;
        495:
            _10305 <= _1212;
        496:
            _10305 <= _1203;
        497:
            _10305 <= _1194;
        498:
            _10305 <= _1185;
        499:
            _10305 <= _1176;
        500:
            _10305 <= _1167;
        501:
            _10305 <= _1158;
        502:
            _10305 <= _1149;
        503:
            _10305 <= _1140;
        504:
            _10305 <= _1131;
        505:
            _10305 <= _1122;
        506:
            _10305 <= _1113;
        507:
            _10305 <= _1104;
        508:
            _10305 <= _1095;
        509:
            _10305 <= _1086;
        510:
            _10305 <= _1077;
        default:
            _10305 <= _1068;
        endcase
    end
    assign _1063 = 9'b111111111;
    assign _1064 = _1062 == _1063;
    assign _1065 = _1059 & _1064;
    assign _1069 = _1065 ? _515 : _1068;
    assign _1071 = _1047 ? _1055 : _1069;
    assign _3 = _1071;
    always @(posedge _1038) begin
        if (_1036)
            _1068 <= _1055;
        else
            _1068 <= _3;
    end
    assign _1072 = 9'b111111110;
    assign _1073 = _1062 == _1072;
    assign _1074 = _1059 & _1073;
    assign _1078 = _1074 ? _515 : _1077;
    assign _1080 = _1047 ? _1055 : _1078;
    assign _4 = _1080;
    always @(posedge _1038) begin
        if (_1036)
            _1077 <= _1055;
        else
            _1077 <= _4;
    end
    assign _1081 = 9'b111111101;
    assign _1082 = _1062 == _1081;
    assign _1083 = _1059 & _1082;
    assign _1087 = _1083 ? _515 : _1086;
    assign _1089 = _1047 ? _1055 : _1087;
    assign _5 = _1089;
    always @(posedge _1038) begin
        if (_1036)
            _1086 <= _1055;
        else
            _1086 <= _5;
    end
    assign _1090 = 9'b111111100;
    assign _1091 = _1062 == _1090;
    assign _1092 = _1059 & _1091;
    assign _1096 = _1092 ? _515 : _1095;
    assign _1098 = _1047 ? _1055 : _1096;
    assign _6 = _1098;
    always @(posedge _1038) begin
        if (_1036)
            _1095 <= _1055;
        else
            _1095 <= _6;
    end
    assign _1099 = 9'b111111011;
    assign _1100 = _1062 == _1099;
    assign _1101 = _1059 & _1100;
    assign _1105 = _1101 ? _515 : _1104;
    assign _1107 = _1047 ? _1055 : _1105;
    assign _7 = _1107;
    always @(posedge _1038) begin
        if (_1036)
            _1104 <= _1055;
        else
            _1104 <= _7;
    end
    assign _1108 = 9'b111111010;
    assign _1109 = _1062 == _1108;
    assign _1110 = _1059 & _1109;
    assign _1114 = _1110 ? _515 : _1113;
    assign _1116 = _1047 ? _1055 : _1114;
    assign _8 = _1116;
    always @(posedge _1038) begin
        if (_1036)
            _1113 <= _1055;
        else
            _1113 <= _8;
    end
    assign _1117 = 9'b111111001;
    assign _1118 = _1062 == _1117;
    assign _1119 = _1059 & _1118;
    assign _1123 = _1119 ? _515 : _1122;
    assign _1125 = _1047 ? _1055 : _1123;
    assign _9 = _1125;
    always @(posedge _1038) begin
        if (_1036)
            _1122 <= _1055;
        else
            _1122 <= _9;
    end
    assign _1126 = 9'b111111000;
    assign _1127 = _1062 == _1126;
    assign _1128 = _1059 & _1127;
    assign _1132 = _1128 ? _515 : _1131;
    assign _1134 = _1047 ? _1055 : _1132;
    assign _10 = _1134;
    always @(posedge _1038) begin
        if (_1036)
            _1131 <= _1055;
        else
            _1131 <= _10;
    end
    assign _1135 = 9'b111110111;
    assign _1136 = _1062 == _1135;
    assign _1137 = _1059 & _1136;
    assign _1141 = _1137 ? _515 : _1140;
    assign _1143 = _1047 ? _1055 : _1141;
    assign _11 = _1143;
    always @(posedge _1038) begin
        if (_1036)
            _1140 <= _1055;
        else
            _1140 <= _11;
    end
    assign _1144 = 9'b111110110;
    assign _1145 = _1062 == _1144;
    assign _1146 = _1059 & _1145;
    assign _1150 = _1146 ? _515 : _1149;
    assign _1152 = _1047 ? _1055 : _1150;
    assign _12 = _1152;
    always @(posedge _1038) begin
        if (_1036)
            _1149 <= _1055;
        else
            _1149 <= _12;
    end
    assign _1153 = 9'b111110101;
    assign _1154 = _1062 == _1153;
    assign _1155 = _1059 & _1154;
    assign _1159 = _1155 ? _515 : _1158;
    assign _1161 = _1047 ? _1055 : _1159;
    assign _13 = _1161;
    always @(posedge _1038) begin
        if (_1036)
            _1158 <= _1055;
        else
            _1158 <= _13;
    end
    assign _1162 = 9'b111110100;
    assign _1163 = _1062 == _1162;
    assign _1164 = _1059 & _1163;
    assign _1168 = _1164 ? _515 : _1167;
    assign _1170 = _1047 ? _1055 : _1168;
    assign _14 = _1170;
    always @(posedge _1038) begin
        if (_1036)
            _1167 <= _1055;
        else
            _1167 <= _14;
    end
    assign _1171 = 9'b111110011;
    assign _1172 = _1062 == _1171;
    assign _1173 = _1059 & _1172;
    assign _1177 = _1173 ? _515 : _1176;
    assign _1179 = _1047 ? _1055 : _1177;
    assign _15 = _1179;
    always @(posedge _1038) begin
        if (_1036)
            _1176 <= _1055;
        else
            _1176 <= _15;
    end
    assign _1180 = 9'b111110010;
    assign _1181 = _1062 == _1180;
    assign _1182 = _1059 & _1181;
    assign _1186 = _1182 ? _515 : _1185;
    assign _1188 = _1047 ? _1055 : _1186;
    assign _16 = _1188;
    always @(posedge _1038) begin
        if (_1036)
            _1185 <= _1055;
        else
            _1185 <= _16;
    end
    assign _1189 = 9'b111110001;
    assign _1190 = _1062 == _1189;
    assign _1191 = _1059 & _1190;
    assign _1195 = _1191 ? _515 : _1194;
    assign _1197 = _1047 ? _1055 : _1195;
    assign _17 = _1197;
    always @(posedge _1038) begin
        if (_1036)
            _1194 <= _1055;
        else
            _1194 <= _17;
    end
    assign _1198 = 9'b111110000;
    assign _1199 = _1062 == _1198;
    assign _1200 = _1059 & _1199;
    assign _1204 = _1200 ? _515 : _1203;
    assign _1206 = _1047 ? _1055 : _1204;
    assign _18 = _1206;
    always @(posedge _1038) begin
        if (_1036)
            _1203 <= _1055;
        else
            _1203 <= _18;
    end
    assign _1207 = 9'b111101111;
    assign _1208 = _1062 == _1207;
    assign _1209 = _1059 & _1208;
    assign _1213 = _1209 ? _515 : _1212;
    assign _1215 = _1047 ? _1055 : _1213;
    assign _19 = _1215;
    always @(posedge _1038) begin
        if (_1036)
            _1212 <= _1055;
        else
            _1212 <= _19;
    end
    assign _1216 = 9'b111101110;
    assign _1217 = _1062 == _1216;
    assign _1218 = _1059 & _1217;
    assign _1222 = _1218 ? _515 : _1221;
    assign _1224 = _1047 ? _1055 : _1222;
    assign _20 = _1224;
    always @(posedge _1038) begin
        if (_1036)
            _1221 <= _1055;
        else
            _1221 <= _20;
    end
    assign _1225 = 9'b111101101;
    assign _1226 = _1062 == _1225;
    assign _1227 = _1059 & _1226;
    assign _1231 = _1227 ? _515 : _1230;
    assign _1233 = _1047 ? _1055 : _1231;
    assign _21 = _1233;
    always @(posedge _1038) begin
        if (_1036)
            _1230 <= _1055;
        else
            _1230 <= _21;
    end
    assign _1234 = 9'b111101100;
    assign _1235 = _1062 == _1234;
    assign _1236 = _1059 & _1235;
    assign _1240 = _1236 ? _515 : _1239;
    assign _1242 = _1047 ? _1055 : _1240;
    assign _22 = _1242;
    always @(posedge _1038) begin
        if (_1036)
            _1239 <= _1055;
        else
            _1239 <= _22;
    end
    assign _1243 = 9'b111101011;
    assign _1244 = _1062 == _1243;
    assign _1245 = _1059 & _1244;
    assign _1249 = _1245 ? _515 : _1248;
    assign _1251 = _1047 ? _1055 : _1249;
    assign _23 = _1251;
    always @(posedge _1038) begin
        if (_1036)
            _1248 <= _1055;
        else
            _1248 <= _23;
    end
    assign _1252 = 9'b111101010;
    assign _1253 = _1062 == _1252;
    assign _1254 = _1059 & _1253;
    assign _1258 = _1254 ? _515 : _1257;
    assign _1260 = _1047 ? _1055 : _1258;
    assign _24 = _1260;
    always @(posedge _1038) begin
        if (_1036)
            _1257 <= _1055;
        else
            _1257 <= _24;
    end
    assign _1261 = 9'b111101001;
    assign _1262 = _1062 == _1261;
    assign _1263 = _1059 & _1262;
    assign _1267 = _1263 ? _515 : _1266;
    assign _1269 = _1047 ? _1055 : _1267;
    assign _25 = _1269;
    always @(posedge _1038) begin
        if (_1036)
            _1266 <= _1055;
        else
            _1266 <= _25;
    end
    assign _1270 = 9'b111101000;
    assign _1271 = _1062 == _1270;
    assign _1272 = _1059 & _1271;
    assign _1276 = _1272 ? _515 : _1275;
    assign _1278 = _1047 ? _1055 : _1276;
    assign _26 = _1278;
    always @(posedge _1038) begin
        if (_1036)
            _1275 <= _1055;
        else
            _1275 <= _26;
    end
    assign _1279 = 9'b111100111;
    assign _1280 = _1062 == _1279;
    assign _1281 = _1059 & _1280;
    assign _1285 = _1281 ? _515 : _1284;
    assign _1287 = _1047 ? _1055 : _1285;
    assign _27 = _1287;
    always @(posedge _1038) begin
        if (_1036)
            _1284 <= _1055;
        else
            _1284 <= _27;
    end
    assign _1288 = 9'b111100110;
    assign _1289 = _1062 == _1288;
    assign _1290 = _1059 & _1289;
    assign _1294 = _1290 ? _515 : _1293;
    assign _1296 = _1047 ? _1055 : _1294;
    assign _28 = _1296;
    always @(posedge _1038) begin
        if (_1036)
            _1293 <= _1055;
        else
            _1293 <= _28;
    end
    assign _1297 = 9'b111100101;
    assign _1298 = _1062 == _1297;
    assign _1299 = _1059 & _1298;
    assign _1303 = _1299 ? _515 : _1302;
    assign _1305 = _1047 ? _1055 : _1303;
    assign _29 = _1305;
    always @(posedge _1038) begin
        if (_1036)
            _1302 <= _1055;
        else
            _1302 <= _29;
    end
    assign _1306 = 9'b111100100;
    assign _1307 = _1062 == _1306;
    assign _1308 = _1059 & _1307;
    assign _1312 = _1308 ? _515 : _1311;
    assign _1314 = _1047 ? _1055 : _1312;
    assign _30 = _1314;
    always @(posedge _1038) begin
        if (_1036)
            _1311 <= _1055;
        else
            _1311 <= _30;
    end
    assign _1315 = 9'b111100011;
    assign _1316 = _1062 == _1315;
    assign _1317 = _1059 & _1316;
    assign _1321 = _1317 ? _515 : _1320;
    assign _1323 = _1047 ? _1055 : _1321;
    assign _31 = _1323;
    always @(posedge _1038) begin
        if (_1036)
            _1320 <= _1055;
        else
            _1320 <= _31;
    end
    assign _1324 = 9'b111100010;
    assign _1325 = _1062 == _1324;
    assign _1326 = _1059 & _1325;
    assign _1330 = _1326 ? _515 : _1329;
    assign _1332 = _1047 ? _1055 : _1330;
    assign _32 = _1332;
    always @(posedge _1038) begin
        if (_1036)
            _1329 <= _1055;
        else
            _1329 <= _32;
    end
    assign _1333 = 9'b111100001;
    assign _1334 = _1062 == _1333;
    assign _1335 = _1059 & _1334;
    assign _1339 = _1335 ? _515 : _1338;
    assign _1341 = _1047 ? _1055 : _1339;
    assign _33 = _1341;
    always @(posedge _1038) begin
        if (_1036)
            _1338 <= _1055;
        else
            _1338 <= _33;
    end
    assign _1342 = 9'b111100000;
    assign _1343 = _1062 == _1342;
    assign _1344 = _1059 & _1343;
    assign _1348 = _1344 ? _515 : _1347;
    assign _1350 = _1047 ? _1055 : _1348;
    assign _34 = _1350;
    always @(posedge _1038) begin
        if (_1036)
            _1347 <= _1055;
        else
            _1347 <= _34;
    end
    assign _1351 = 9'b111011111;
    assign _1352 = _1062 == _1351;
    assign _1353 = _1059 & _1352;
    assign _1357 = _1353 ? _515 : _1356;
    assign _1359 = _1047 ? _1055 : _1357;
    assign _35 = _1359;
    always @(posedge _1038) begin
        if (_1036)
            _1356 <= _1055;
        else
            _1356 <= _35;
    end
    assign _1360 = 9'b111011110;
    assign _1361 = _1062 == _1360;
    assign _1362 = _1059 & _1361;
    assign _1366 = _1362 ? _515 : _1365;
    assign _1368 = _1047 ? _1055 : _1366;
    assign _36 = _1368;
    always @(posedge _1038) begin
        if (_1036)
            _1365 <= _1055;
        else
            _1365 <= _36;
    end
    assign _1369 = 9'b111011101;
    assign _1370 = _1062 == _1369;
    assign _1371 = _1059 & _1370;
    assign _1375 = _1371 ? _515 : _1374;
    assign _1377 = _1047 ? _1055 : _1375;
    assign _37 = _1377;
    always @(posedge _1038) begin
        if (_1036)
            _1374 <= _1055;
        else
            _1374 <= _37;
    end
    assign _1378 = 9'b111011100;
    assign _1379 = _1062 == _1378;
    assign _1380 = _1059 & _1379;
    assign _1384 = _1380 ? _515 : _1383;
    assign _1386 = _1047 ? _1055 : _1384;
    assign _38 = _1386;
    always @(posedge _1038) begin
        if (_1036)
            _1383 <= _1055;
        else
            _1383 <= _38;
    end
    assign _1387 = 9'b111011011;
    assign _1388 = _1062 == _1387;
    assign _1389 = _1059 & _1388;
    assign _1393 = _1389 ? _515 : _1392;
    assign _1395 = _1047 ? _1055 : _1393;
    assign _39 = _1395;
    always @(posedge _1038) begin
        if (_1036)
            _1392 <= _1055;
        else
            _1392 <= _39;
    end
    assign _1396 = 9'b111011010;
    assign _1397 = _1062 == _1396;
    assign _1398 = _1059 & _1397;
    assign _1402 = _1398 ? _515 : _1401;
    assign _1404 = _1047 ? _1055 : _1402;
    assign _40 = _1404;
    always @(posedge _1038) begin
        if (_1036)
            _1401 <= _1055;
        else
            _1401 <= _40;
    end
    assign _1405 = 9'b111011001;
    assign _1406 = _1062 == _1405;
    assign _1407 = _1059 & _1406;
    assign _1411 = _1407 ? _515 : _1410;
    assign _1413 = _1047 ? _1055 : _1411;
    assign _41 = _1413;
    always @(posedge _1038) begin
        if (_1036)
            _1410 <= _1055;
        else
            _1410 <= _41;
    end
    assign _1414 = 9'b111011000;
    assign _1415 = _1062 == _1414;
    assign _1416 = _1059 & _1415;
    assign _1420 = _1416 ? _515 : _1419;
    assign _1422 = _1047 ? _1055 : _1420;
    assign _42 = _1422;
    always @(posedge _1038) begin
        if (_1036)
            _1419 <= _1055;
        else
            _1419 <= _42;
    end
    assign _1423 = 9'b111010111;
    assign _1424 = _1062 == _1423;
    assign _1425 = _1059 & _1424;
    assign _1429 = _1425 ? _515 : _1428;
    assign _1431 = _1047 ? _1055 : _1429;
    assign _43 = _1431;
    always @(posedge _1038) begin
        if (_1036)
            _1428 <= _1055;
        else
            _1428 <= _43;
    end
    assign _1432 = 9'b111010110;
    assign _1433 = _1062 == _1432;
    assign _1434 = _1059 & _1433;
    assign _1438 = _1434 ? _515 : _1437;
    assign _1440 = _1047 ? _1055 : _1438;
    assign _44 = _1440;
    always @(posedge _1038) begin
        if (_1036)
            _1437 <= _1055;
        else
            _1437 <= _44;
    end
    assign _1441 = 9'b111010101;
    assign _1442 = _1062 == _1441;
    assign _1443 = _1059 & _1442;
    assign _1447 = _1443 ? _515 : _1446;
    assign _1449 = _1047 ? _1055 : _1447;
    assign _45 = _1449;
    always @(posedge _1038) begin
        if (_1036)
            _1446 <= _1055;
        else
            _1446 <= _45;
    end
    assign _1450 = 9'b111010100;
    assign _1451 = _1062 == _1450;
    assign _1452 = _1059 & _1451;
    assign _1456 = _1452 ? _515 : _1455;
    assign _1458 = _1047 ? _1055 : _1456;
    assign _46 = _1458;
    always @(posedge _1038) begin
        if (_1036)
            _1455 <= _1055;
        else
            _1455 <= _46;
    end
    assign _1459 = 9'b111010011;
    assign _1460 = _1062 == _1459;
    assign _1461 = _1059 & _1460;
    assign _1465 = _1461 ? _515 : _1464;
    assign _1467 = _1047 ? _1055 : _1465;
    assign _47 = _1467;
    always @(posedge _1038) begin
        if (_1036)
            _1464 <= _1055;
        else
            _1464 <= _47;
    end
    assign _1468 = 9'b111010010;
    assign _1469 = _1062 == _1468;
    assign _1470 = _1059 & _1469;
    assign _1474 = _1470 ? _515 : _1473;
    assign _1476 = _1047 ? _1055 : _1474;
    assign _48 = _1476;
    always @(posedge _1038) begin
        if (_1036)
            _1473 <= _1055;
        else
            _1473 <= _48;
    end
    assign _1477 = 9'b111010001;
    assign _1478 = _1062 == _1477;
    assign _1479 = _1059 & _1478;
    assign _1483 = _1479 ? _515 : _1482;
    assign _1485 = _1047 ? _1055 : _1483;
    assign _49 = _1485;
    always @(posedge _1038) begin
        if (_1036)
            _1482 <= _1055;
        else
            _1482 <= _49;
    end
    assign _1486 = 9'b111010000;
    assign _1487 = _1062 == _1486;
    assign _1488 = _1059 & _1487;
    assign _1492 = _1488 ? _515 : _1491;
    assign _1494 = _1047 ? _1055 : _1492;
    assign _50 = _1494;
    always @(posedge _1038) begin
        if (_1036)
            _1491 <= _1055;
        else
            _1491 <= _50;
    end
    assign _1495 = 9'b111001111;
    assign _1496 = _1062 == _1495;
    assign _1497 = _1059 & _1496;
    assign _1501 = _1497 ? _515 : _1500;
    assign _1503 = _1047 ? _1055 : _1501;
    assign _51 = _1503;
    always @(posedge _1038) begin
        if (_1036)
            _1500 <= _1055;
        else
            _1500 <= _51;
    end
    assign _1504 = 9'b111001110;
    assign _1505 = _1062 == _1504;
    assign _1506 = _1059 & _1505;
    assign _1510 = _1506 ? _515 : _1509;
    assign _1512 = _1047 ? _1055 : _1510;
    assign _52 = _1512;
    always @(posedge _1038) begin
        if (_1036)
            _1509 <= _1055;
        else
            _1509 <= _52;
    end
    assign _1513 = 9'b111001101;
    assign _1514 = _1062 == _1513;
    assign _1515 = _1059 & _1514;
    assign _1519 = _1515 ? _515 : _1518;
    assign _1521 = _1047 ? _1055 : _1519;
    assign _53 = _1521;
    always @(posedge _1038) begin
        if (_1036)
            _1518 <= _1055;
        else
            _1518 <= _53;
    end
    assign _1522 = 9'b111001100;
    assign _1523 = _1062 == _1522;
    assign _1524 = _1059 & _1523;
    assign _1528 = _1524 ? _515 : _1527;
    assign _1530 = _1047 ? _1055 : _1528;
    assign _54 = _1530;
    always @(posedge _1038) begin
        if (_1036)
            _1527 <= _1055;
        else
            _1527 <= _54;
    end
    assign _1531 = 9'b111001011;
    assign _1532 = _1062 == _1531;
    assign _1533 = _1059 & _1532;
    assign _1537 = _1533 ? _515 : _1536;
    assign _1539 = _1047 ? _1055 : _1537;
    assign _55 = _1539;
    always @(posedge _1038) begin
        if (_1036)
            _1536 <= _1055;
        else
            _1536 <= _55;
    end
    assign _1540 = 9'b111001010;
    assign _1541 = _1062 == _1540;
    assign _1542 = _1059 & _1541;
    assign _1546 = _1542 ? _515 : _1545;
    assign _1548 = _1047 ? _1055 : _1546;
    assign _56 = _1548;
    always @(posedge _1038) begin
        if (_1036)
            _1545 <= _1055;
        else
            _1545 <= _56;
    end
    assign _1549 = 9'b111001001;
    assign _1550 = _1062 == _1549;
    assign _1551 = _1059 & _1550;
    assign _1555 = _1551 ? _515 : _1554;
    assign _1557 = _1047 ? _1055 : _1555;
    assign _57 = _1557;
    always @(posedge _1038) begin
        if (_1036)
            _1554 <= _1055;
        else
            _1554 <= _57;
    end
    assign _1558 = 9'b111001000;
    assign _1559 = _1062 == _1558;
    assign _1560 = _1059 & _1559;
    assign _1564 = _1560 ? _515 : _1563;
    assign _1566 = _1047 ? _1055 : _1564;
    assign _58 = _1566;
    always @(posedge _1038) begin
        if (_1036)
            _1563 <= _1055;
        else
            _1563 <= _58;
    end
    assign _1567 = 9'b111000111;
    assign _1568 = _1062 == _1567;
    assign _1569 = _1059 & _1568;
    assign _1573 = _1569 ? _515 : _1572;
    assign _1575 = _1047 ? _1055 : _1573;
    assign _59 = _1575;
    always @(posedge _1038) begin
        if (_1036)
            _1572 <= _1055;
        else
            _1572 <= _59;
    end
    assign _1576 = 9'b111000110;
    assign _1577 = _1062 == _1576;
    assign _1578 = _1059 & _1577;
    assign _1582 = _1578 ? _515 : _1581;
    assign _1584 = _1047 ? _1055 : _1582;
    assign _60 = _1584;
    always @(posedge _1038) begin
        if (_1036)
            _1581 <= _1055;
        else
            _1581 <= _60;
    end
    assign _1585 = 9'b111000101;
    assign _1586 = _1062 == _1585;
    assign _1587 = _1059 & _1586;
    assign _1591 = _1587 ? _515 : _1590;
    assign _1593 = _1047 ? _1055 : _1591;
    assign _61 = _1593;
    always @(posedge _1038) begin
        if (_1036)
            _1590 <= _1055;
        else
            _1590 <= _61;
    end
    assign _1594 = 9'b111000100;
    assign _1595 = _1062 == _1594;
    assign _1596 = _1059 & _1595;
    assign _1600 = _1596 ? _515 : _1599;
    assign _1602 = _1047 ? _1055 : _1600;
    assign _62 = _1602;
    always @(posedge _1038) begin
        if (_1036)
            _1599 <= _1055;
        else
            _1599 <= _62;
    end
    assign _1603 = 9'b111000011;
    assign _1604 = _1062 == _1603;
    assign _1605 = _1059 & _1604;
    assign _1609 = _1605 ? _515 : _1608;
    assign _1611 = _1047 ? _1055 : _1609;
    assign _63 = _1611;
    always @(posedge _1038) begin
        if (_1036)
            _1608 <= _1055;
        else
            _1608 <= _63;
    end
    assign _1612 = 9'b111000010;
    assign _1613 = _1062 == _1612;
    assign _1614 = _1059 & _1613;
    assign _1618 = _1614 ? _515 : _1617;
    assign _1620 = _1047 ? _1055 : _1618;
    assign _64 = _1620;
    always @(posedge _1038) begin
        if (_1036)
            _1617 <= _1055;
        else
            _1617 <= _64;
    end
    assign _1621 = 9'b111000001;
    assign _1622 = _1062 == _1621;
    assign _1623 = _1059 & _1622;
    assign _1627 = _1623 ? _515 : _1626;
    assign _1629 = _1047 ? _1055 : _1627;
    assign _65 = _1629;
    always @(posedge _1038) begin
        if (_1036)
            _1626 <= _1055;
        else
            _1626 <= _65;
    end
    assign _1630 = 9'b111000000;
    assign _1631 = _1062 == _1630;
    assign _1632 = _1059 & _1631;
    assign _1636 = _1632 ? _515 : _1635;
    assign _1638 = _1047 ? _1055 : _1636;
    assign _66 = _1638;
    always @(posedge _1038) begin
        if (_1036)
            _1635 <= _1055;
        else
            _1635 <= _66;
    end
    assign _1639 = 9'b110111111;
    assign _1640 = _1062 == _1639;
    assign _1641 = _1059 & _1640;
    assign _1645 = _1641 ? _515 : _1644;
    assign _1647 = _1047 ? _1055 : _1645;
    assign _67 = _1647;
    always @(posedge _1038) begin
        if (_1036)
            _1644 <= _1055;
        else
            _1644 <= _67;
    end
    assign _1648 = 9'b110111110;
    assign _1649 = _1062 == _1648;
    assign _1650 = _1059 & _1649;
    assign _1654 = _1650 ? _515 : _1653;
    assign _1656 = _1047 ? _1055 : _1654;
    assign _68 = _1656;
    always @(posedge _1038) begin
        if (_1036)
            _1653 <= _1055;
        else
            _1653 <= _68;
    end
    assign _1657 = 9'b110111101;
    assign _1658 = _1062 == _1657;
    assign _1659 = _1059 & _1658;
    assign _1663 = _1659 ? _515 : _1662;
    assign _1665 = _1047 ? _1055 : _1663;
    assign _69 = _1665;
    always @(posedge _1038) begin
        if (_1036)
            _1662 <= _1055;
        else
            _1662 <= _69;
    end
    assign _1666 = 9'b110111100;
    assign _1667 = _1062 == _1666;
    assign _1668 = _1059 & _1667;
    assign _1672 = _1668 ? _515 : _1671;
    assign _1674 = _1047 ? _1055 : _1672;
    assign _70 = _1674;
    always @(posedge _1038) begin
        if (_1036)
            _1671 <= _1055;
        else
            _1671 <= _70;
    end
    assign _1675 = 9'b110111011;
    assign _1676 = _1062 == _1675;
    assign _1677 = _1059 & _1676;
    assign _1681 = _1677 ? _515 : _1680;
    assign _1683 = _1047 ? _1055 : _1681;
    assign _71 = _1683;
    always @(posedge _1038) begin
        if (_1036)
            _1680 <= _1055;
        else
            _1680 <= _71;
    end
    assign _1684 = 9'b110111010;
    assign _1685 = _1062 == _1684;
    assign _1686 = _1059 & _1685;
    assign _1690 = _1686 ? _515 : _1689;
    assign _1692 = _1047 ? _1055 : _1690;
    assign _72 = _1692;
    always @(posedge _1038) begin
        if (_1036)
            _1689 <= _1055;
        else
            _1689 <= _72;
    end
    assign _1693 = 9'b110111001;
    assign _1694 = _1062 == _1693;
    assign _1695 = _1059 & _1694;
    assign _1699 = _1695 ? _515 : _1698;
    assign _1701 = _1047 ? _1055 : _1699;
    assign _73 = _1701;
    always @(posedge _1038) begin
        if (_1036)
            _1698 <= _1055;
        else
            _1698 <= _73;
    end
    assign _1702 = 9'b110111000;
    assign _1703 = _1062 == _1702;
    assign _1704 = _1059 & _1703;
    assign _1708 = _1704 ? _515 : _1707;
    assign _1710 = _1047 ? _1055 : _1708;
    assign _74 = _1710;
    always @(posedge _1038) begin
        if (_1036)
            _1707 <= _1055;
        else
            _1707 <= _74;
    end
    assign _1711 = 9'b110110111;
    assign _1712 = _1062 == _1711;
    assign _1713 = _1059 & _1712;
    assign _1717 = _1713 ? _515 : _1716;
    assign _1719 = _1047 ? _1055 : _1717;
    assign _75 = _1719;
    always @(posedge _1038) begin
        if (_1036)
            _1716 <= _1055;
        else
            _1716 <= _75;
    end
    assign _1720 = 9'b110110110;
    assign _1721 = _1062 == _1720;
    assign _1722 = _1059 & _1721;
    assign _1726 = _1722 ? _515 : _1725;
    assign _1728 = _1047 ? _1055 : _1726;
    assign _76 = _1728;
    always @(posedge _1038) begin
        if (_1036)
            _1725 <= _1055;
        else
            _1725 <= _76;
    end
    assign _1729 = 9'b110110101;
    assign _1730 = _1062 == _1729;
    assign _1731 = _1059 & _1730;
    assign _1735 = _1731 ? _515 : _1734;
    assign _1737 = _1047 ? _1055 : _1735;
    assign _77 = _1737;
    always @(posedge _1038) begin
        if (_1036)
            _1734 <= _1055;
        else
            _1734 <= _77;
    end
    assign _1738 = 9'b110110100;
    assign _1739 = _1062 == _1738;
    assign _1740 = _1059 & _1739;
    assign _1744 = _1740 ? _515 : _1743;
    assign _1746 = _1047 ? _1055 : _1744;
    assign _78 = _1746;
    always @(posedge _1038) begin
        if (_1036)
            _1743 <= _1055;
        else
            _1743 <= _78;
    end
    assign _1747 = 9'b110110011;
    assign _1748 = _1062 == _1747;
    assign _1749 = _1059 & _1748;
    assign _1753 = _1749 ? _515 : _1752;
    assign _1755 = _1047 ? _1055 : _1753;
    assign _79 = _1755;
    always @(posedge _1038) begin
        if (_1036)
            _1752 <= _1055;
        else
            _1752 <= _79;
    end
    assign _1756 = 9'b110110010;
    assign _1757 = _1062 == _1756;
    assign _1758 = _1059 & _1757;
    assign _1762 = _1758 ? _515 : _1761;
    assign _1764 = _1047 ? _1055 : _1762;
    assign _80 = _1764;
    always @(posedge _1038) begin
        if (_1036)
            _1761 <= _1055;
        else
            _1761 <= _80;
    end
    assign _1765 = 9'b110110001;
    assign _1766 = _1062 == _1765;
    assign _1767 = _1059 & _1766;
    assign _1771 = _1767 ? _515 : _1770;
    assign _1773 = _1047 ? _1055 : _1771;
    assign _81 = _1773;
    always @(posedge _1038) begin
        if (_1036)
            _1770 <= _1055;
        else
            _1770 <= _81;
    end
    assign _1774 = 9'b110110000;
    assign _1775 = _1062 == _1774;
    assign _1776 = _1059 & _1775;
    assign _1780 = _1776 ? _515 : _1779;
    assign _1782 = _1047 ? _1055 : _1780;
    assign _82 = _1782;
    always @(posedge _1038) begin
        if (_1036)
            _1779 <= _1055;
        else
            _1779 <= _82;
    end
    assign _1783 = 9'b110101111;
    assign _1784 = _1062 == _1783;
    assign _1785 = _1059 & _1784;
    assign _1789 = _1785 ? _515 : _1788;
    assign _1791 = _1047 ? _1055 : _1789;
    assign _83 = _1791;
    always @(posedge _1038) begin
        if (_1036)
            _1788 <= _1055;
        else
            _1788 <= _83;
    end
    assign _1792 = 9'b110101110;
    assign _1793 = _1062 == _1792;
    assign _1794 = _1059 & _1793;
    assign _1798 = _1794 ? _515 : _1797;
    assign _1800 = _1047 ? _1055 : _1798;
    assign _84 = _1800;
    always @(posedge _1038) begin
        if (_1036)
            _1797 <= _1055;
        else
            _1797 <= _84;
    end
    assign _1801 = 9'b110101101;
    assign _1802 = _1062 == _1801;
    assign _1803 = _1059 & _1802;
    assign _1807 = _1803 ? _515 : _1806;
    assign _1809 = _1047 ? _1055 : _1807;
    assign _85 = _1809;
    always @(posedge _1038) begin
        if (_1036)
            _1806 <= _1055;
        else
            _1806 <= _85;
    end
    assign _1810 = 9'b110101100;
    assign _1811 = _1062 == _1810;
    assign _1812 = _1059 & _1811;
    assign _1816 = _1812 ? _515 : _1815;
    assign _1818 = _1047 ? _1055 : _1816;
    assign _86 = _1818;
    always @(posedge _1038) begin
        if (_1036)
            _1815 <= _1055;
        else
            _1815 <= _86;
    end
    assign _1819 = 9'b110101011;
    assign _1820 = _1062 == _1819;
    assign _1821 = _1059 & _1820;
    assign _1825 = _1821 ? _515 : _1824;
    assign _1827 = _1047 ? _1055 : _1825;
    assign _87 = _1827;
    always @(posedge _1038) begin
        if (_1036)
            _1824 <= _1055;
        else
            _1824 <= _87;
    end
    assign _1828 = 9'b110101010;
    assign _1829 = _1062 == _1828;
    assign _1830 = _1059 & _1829;
    assign _1834 = _1830 ? _515 : _1833;
    assign _1836 = _1047 ? _1055 : _1834;
    assign _88 = _1836;
    always @(posedge _1038) begin
        if (_1036)
            _1833 <= _1055;
        else
            _1833 <= _88;
    end
    assign _1837 = 9'b110101001;
    assign _1838 = _1062 == _1837;
    assign _1839 = _1059 & _1838;
    assign _1843 = _1839 ? _515 : _1842;
    assign _1845 = _1047 ? _1055 : _1843;
    assign _89 = _1845;
    always @(posedge _1038) begin
        if (_1036)
            _1842 <= _1055;
        else
            _1842 <= _89;
    end
    assign _1846 = 9'b110101000;
    assign _1847 = _1062 == _1846;
    assign _1848 = _1059 & _1847;
    assign _1852 = _1848 ? _515 : _1851;
    assign _1854 = _1047 ? _1055 : _1852;
    assign _90 = _1854;
    always @(posedge _1038) begin
        if (_1036)
            _1851 <= _1055;
        else
            _1851 <= _90;
    end
    assign _1855 = 9'b110100111;
    assign _1856 = _1062 == _1855;
    assign _1857 = _1059 & _1856;
    assign _1861 = _1857 ? _515 : _1860;
    assign _1863 = _1047 ? _1055 : _1861;
    assign _91 = _1863;
    always @(posedge _1038) begin
        if (_1036)
            _1860 <= _1055;
        else
            _1860 <= _91;
    end
    assign _1864 = 9'b110100110;
    assign _1865 = _1062 == _1864;
    assign _1866 = _1059 & _1865;
    assign _1870 = _1866 ? _515 : _1869;
    assign _1872 = _1047 ? _1055 : _1870;
    assign _92 = _1872;
    always @(posedge _1038) begin
        if (_1036)
            _1869 <= _1055;
        else
            _1869 <= _92;
    end
    assign _1873 = 9'b110100101;
    assign _1874 = _1062 == _1873;
    assign _1875 = _1059 & _1874;
    assign _1879 = _1875 ? _515 : _1878;
    assign _1881 = _1047 ? _1055 : _1879;
    assign _93 = _1881;
    always @(posedge _1038) begin
        if (_1036)
            _1878 <= _1055;
        else
            _1878 <= _93;
    end
    assign _1882 = 9'b110100100;
    assign _1883 = _1062 == _1882;
    assign _1884 = _1059 & _1883;
    assign _1888 = _1884 ? _515 : _1887;
    assign _1890 = _1047 ? _1055 : _1888;
    assign _94 = _1890;
    always @(posedge _1038) begin
        if (_1036)
            _1887 <= _1055;
        else
            _1887 <= _94;
    end
    assign _1891 = 9'b110100011;
    assign _1892 = _1062 == _1891;
    assign _1893 = _1059 & _1892;
    assign _1897 = _1893 ? _515 : _1896;
    assign _1899 = _1047 ? _1055 : _1897;
    assign _95 = _1899;
    always @(posedge _1038) begin
        if (_1036)
            _1896 <= _1055;
        else
            _1896 <= _95;
    end
    assign _1900 = 9'b110100010;
    assign _1901 = _1062 == _1900;
    assign _1902 = _1059 & _1901;
    assign _1906 = _1902 ? _515 : _1905;
    assign _1908 = _1047 ? _1055 : _1906;
    assign _96 = _1908;
    always @(posedge _1038) begin
        if (_1036)
            _1905 <= _1055;
        else
            _1905 <= _96;
    end
    assign _1909 = 9'b110100001;
    assign _1910 = _1062 == _1909;
    assign _1911 = _1059 & _1910;
    assign _1915 = _1911 ? _515 : _1914;
    assign _1917 = _1047 ? _1055 : _1915;
    assign _97 = _1917;
    always @(posedge _1038) begin
        if (_1036)
            _1914 <= _1055;
        else
            _1914 <= _97;
    end
    assign _1918 = 9'b110100000;
    assign _1919 = _1062 == _1918;
    assign _1920 = _1059 & _1919;
    assign _1924 = _1920 ? _515 : _1923;
    assign _1926 = _1047 ? _1055 : _1924;
    assign _98 = _1926;
    always @(posedge _1038) begin
        if (_1036)
            _1923 <= _1055;
        else
            _1923 <= _98;
    end
    assign _1927 = 9'b110011111;
    assign _1928 = _1062 == _1927;
    assign _1929 = _1059 & _1928;
    assign _1933 = _1929 ? _515 : _1932;
    assign _1935 = _1047 ? _1055 : _1933;
    assign _99 = _1935;
    always @(posedge _1038) begin
        if (_1036)
            _1932 <= _1055;
        else
            _1932 <= _99;
    end
    assign _1936 = 9'b110011110;
    assign _1937 = _1062 == _1936;
    assign _1938 = _1059 & _1937;
    assign _1942 = _1938 ? _515 : _1941;
    assign _1944 = _1047 ? _1055 : _1942;
    assign _100 = _1944;
    always @(posedge _1038) begin
        if (_1036)
            _1941 <= _1055;
        else
            _1941 <= _100;
    end
    assign _1945 = 9'b110011101;
    assign _1946 = _1062 == _1945;
    assign _1947 = _1059 & _1946;
    assign _1951 = _1947 ? _515 : _1950;
    assign _1953 = _1047 ? _1055 : _1951;
    assign _101 = _1953;
    always @(posedge _1038) begin
        if (_1036)
            _1950 <= _1055;
        else
            _1950 <= _101;
    end
    assign _1954 = 9'b110011100;
    assign _1955 = _1062 == _1954;
    assign _1956 = _1059 & _1955;
    assign _1960 = _1956 ? _515 : _1959;
    assign _1962 = _1047 ? _1055 : _1960;
    assign _102 = _1962;
    always @(posedge _1038) begin
        if (_1036)
            _1959 <= _1055;
        else
            _1959 <= _102;
    end
    assign _1963 = 9'b110011011;
    assign _1964 = _1062 == _1963;
    assign _1965 = _1059 & _1964;
    assign _1969 = _1965 ? _515 : _1968;
    assign _1971 = _1047 ? _1055 : _1969;
    assign _103 = _1971;
    always @(posedge _1038) begin
        if (_1036)
            _1968 <= _1055;
        else
            _1968 <= _103;
    end
    assign _1972 = 9'b110011010;
    assign _1973 = _1062 == _1972;
    assign _1974 = _1059 & _1973;
    assign _1978 = _1974 ? _515 : _1977;
    assign _1980 = _1047 ? _1055 : _1978;
    assign _104 = _1980;
    always @(posedge _1038) begin
        if (_1036)
            _1977 <= _1055;
        else
            _1977 <= _104;
    end
    assign _1981 = 9'b110011001;
    assign _1982 = _1062 == _1981;
    assign _1983 = _1059 & _1982;
    assign _1987 = _1983 ? _515 : _1986;
    assign _1989 = _1047 ? _1055 : _1987;
    assign _105 = _1989;
    always @(posedge _1038) begin
        if (_1036)
            _1986 <= _1055;
        else
            _1986 <= _105;
    end
    assign _1990 = 9'b110011000;
    assign _1991 = _1062 == _1990;
    assign _1992 = _1059 & _1991;
    assign _1996 = _1992 ? _515 : _1995;
    assign _1998 = _1047 ? _1055 : _1996;
    assign _106 = _1998;
    always @(posedge _1038) begin
        if (_1036)
            _1995 <= _1055;
        else
            _1995 <= _106;
    end
    assign _1999 = 9'b110010111;
    assign _2000 = _1062 == _1999;
    assign _2001 = _1059 & _2000;
    assign _2005 = _2001 ? _515 : _2004;
    assign _2007 = _1047 ? _1055 : _2005;
    assign _107 = _2007;
    always @(posedge _1038) begin
        if (_1036)
            _2004 <= _1055;
        else
            _2004 <= _107;
    end
    assign _2008 = 9'b110010110;
    assign _2009 = _1062 == _2008;
    assign _2010 = _1059 & _2009;
    assign _2014 = _2010 ? _515 : _2013;
    assign _2016 = _1047 ? _1055 : _2014;
    assign _108 = _2016;
    always @(posedge _1038) begin
        if (_1036)
            _2013 <= _1055;
        else
            _2013 <= _108;
    end
    assign _2017 = 9'b110010101;
    assign _2018 = _1062 == _2017;
    assign _2019 = _1059 & _2018;
    assign _2023 = _2019 ? _515 : _2022;
    assign _2025 = _1047 ? _1055 : _2023;
    assign _109 = _2025;
    always @(posedge _1038) begin
        if (_1036)
            _2022 <= _1055;
        else
            _2022 <= _109;
    end
    assign _2026 = 9'b110010100;
    assign _2027 = _1062 == _2026;
    assign _2028 = _1059 & _2027;
    assign _2032 = _2028 ? _515 : _2031;
    assign _2034 = _1047 ? _1055 : _2032;
    assign _110 = _2034;
    always @(posedge _1038) begin
        if (_1036)
            _2031 <= _1055;
        else
            _2031 <= _110;
    end
    assign _2035 = 9'b110010011;
    assign _2036 = _1062 == _2035;
    assign _2037 = _1059 & _2036;
    assign _2041 = _2037 ? _515 : _2040;
    assign _2043 = _1047 ? _1055 : _2041;
    assign _111 = _2043;
    always @(posedge _1038) begin
        if (_1036)
            _2040 <= _1055;
        else
            _2040 <= _111;
    end
    assign _2044 = 9'b110010010;
    assign _2045 = _1062 == _2044;
    assign _2046 = _1059 & _2045;
    assign _2050 = _2046 ? _515 : _2049;
    assign _2052 = _1047 ? _1055 : _2050;
    assign _112 = _2052;
    always @(posedge _1038) begin
        if (_1036)
            _2049 <= _1055;
        else
            _2049 <= _112;
    end
    assign _2053 = 9'b110010001;
    assign _2054 = _1062 == _2053;
    assign _2055 = _1059 & _2054;
    assign _2059 = _2055 ? _515 : _2058;
    assign _2061 = _1047 ? _1055 : _2059;
    assign _113 = _2061;
    always @(posedge _1038) begin
        if (_1036)
            _2058 <= _1055;
        else
            _2058 <= _113;
    end
    assign _2062 = 9'b110010000;
    assign _2063 = _1062 == _2062;
    assign _2064 = _1059 & _2063;
    assign _2068 = _2064 ? _515 : _2067;
    assign _2070 = _1047 ? _1055 : _2068;
    assign _114 = _2070;
    always @(posedge _1038) begin
        if (_1036)
            _2067 <= _1055;
        else
            _2067 <= _114;
    end
    assign _2071 = 9'b110001111;
    assign _2072 = _1062 == _2071;
    assign _2073 = _1059 & _2072;
    assign _2077 = _2073 ? _515 : _2076;
    assign _2079 = _1047 ? _1055 : _2077;
    assign _115 = _2079;
    always @(posedge _1038) begin
        if (_1036)
            _2076 <= _1055;
        else
            _2076 <= _115;
    end
    assign _2080 = 9'b110001110;
    assign _2081 = _1062 == _2080;
    assign _2082 = _1059 & _2081;
    assign _2086 = _2082 ? _515 : _2085;
    assign _2088 = _1047 ? _1055 : _2086;
    assign _116 = _2088;
    always @(posedge _1038) begin
        if (_1036)
            _2085 <= _1055;
        else
            _2085 <= _116;
    end
    assign _2089 = 9'b110001101;
    assign _2090 = _1062 == _2089;
    assign _2091 = _1059 & _2090;
    assign _2095 = _2091 ? _515 : _2094;
    assign _2097 = _1047 ? _1055 : _2095;
    assign _117 = _2097;
    always @(posedge _1038) begin
        if (_1036)
            _2094 <= _1055;
        else
            _2094 <= _117;
    end
    assign _2098 = 9'b110001100;
    assign _2099 = _1062 == _2098;
    assign _2100 = _1059 & _2099;
    assign _2104 = _2100 ? _515 : _2103;
    assign _2106 = _1047 ? _1055 : _2104;
    assign _118 = _2106;
    always @(posedge _1038) begin
        if (_1036)
            _2103 <= _1055;
        else
            _2103 <= _118;
    end
    assign _2107 = 9'b110001011;
    assign _2108 = _1062 == _2107;
    assign _2109 = _1059 & _2108;
    assign _2113 = _2109 ? _515 : _2112;
    assign _2115 = _1047 ? _1055 : _2113;
    assign _119 = _2115;
    always @(posedge _1038) begin
        if (_1036)
            _2112 <= _1055;
        else
            _2112 <= _119;
    end
    assign _2116 = 9'b110001010;
    assign _2117 = _1062 == _2116;
    assign _2118 = _1059 & _2117;
    assign _2122 = _2118 ? _515 : _2121;
    assign _2124 = _1047 ? _1055 : _2122;
    assign _120 = _2124;
    always @(posedge _1038) begin
        if (_1036)
            _2121 <= _1055;
        else
            _2121 <= _120;
    end
    assign _2125 = 9'b110001001;
    assign _2126 = _1062 == _2125;
    assign _2127 = _1059 & _2126;
    assign _2131 = _2127 ? _515 : _2130;
    assign _2133 = _1047 ? _1055 : _2131;
    assign _121 = _2133;
    always @(posedge _1038) begin
        if (_1036)
            _2130 <= _1055;
        else
            _2130 <= _121;
    end
    assign _2134 = 9'b110001000;
    assign _2135 = _1062 == _2134;
    assign _2136 = _1059 & _2135;
    assign _2140 = _2136 ? _515 : _2139;
    assign _2142 = _1047 ? _1055 : _2140;
    assign _122 = _2142;
    always @(posedge _1038) begin
        if (_1036)
            _2139 <= _1055;
        else
            _2139 <= _122;
    end
    assign _2143 = 9'b110000111;
    assign _2144 = _1062 == _2143;
    assign _2145 = _1059 & _2144;
    assign _2149 = _2145 ? _515 : _2148;
    assign _2151 = _1047 ? _1055 : _2149;
    assign _123 = _2151;
    always @(posedge _1038) begin
        if (_1036)
            _2148 <= _1055;
        else
            _2148 <= _123;
    end
    assign _2152 = 9'b110000110;
    assign _2153 = _1062 == _2152;
    assign _2154 = _1059 & _2153;
    assign _2158 = _2154 ? _515 : _2157;
    assign _2160 = _1047 ? _1055 : _2158;
    assign _124 = _2160;
    always @(posedge _1038) begin
        if (_1036)
            _2157 <= _1055;
        else
            _2157 <= _124;
    end
    assign _2161 = 9'b110000101;
    assign _2162 = _1062 == _2161;
    assign _2163 = _1059 & _2162;
    assign _2167 = _2163 ? _515 : _2166;
    assign _2169 = _1047 ? _1055 : _2167;
    assign _125 = _2169;
    always @(posedge _1038) begin
        if (_1036)
            _2166 <= _1055;
        else
            _2166 <= _125;
    end
    assign _2170 = 9'b110000100;
    assign _2171 = _1062 == _2170;
    assign _2172 = _1059 & _2171;
    assign _2176 = _2172 ? _515 : _2175;
    assign _2178 = _1047 ? _1055 : _2176;
    assign _126 = _2178;
    always @(posedge _1038) begin
        if (_1036)
            _2175 <= _1055;
        else
            _2175 <= _126;
    end
    assign _2179 = 9'b110000011;
    assign _2180 = _1062 == _2179;
    assign _2181 = _1059 & _2180;
    assign _2185 = _2181 ? _515 : _2184;
    assign _2187 = _1047 ? _1055 : _2185;
    assign _127 = _2187;
    always @(posedge _1038) begin
        if (_1036)
            _2184 <= _1055;
        else
            _2184 <= _127;
    end
    assign _2188 = 9'b110000010;
    assign _2189 = _1062 == _2188;
    assign _2190 = _1059 & _2189;
    assign _2194 = _2190 ? _515 : _2193;
    assign _2196 = _1047 ? _1055 : _2194;
    assign _128 = _2196;
    always @(posedge _1038) begin
        if (_1036)
            _2193 <= _1055;
        else
            _2193 <= _128;
    end
    assign _2197 = 9'b110000001;
    assign _2198 = _1062 == _2197;
    assign _2199 = _1059 & _2198;
    assign _2203 = _2199 ? _515 : _2202;
    assign _2205 = _1047 ? _1055 : _2203;
    assign _129 = _2205;
    always @(posedge _1038) begin
        if (_1036)
            _2202 <= _1055;
        else
            _2202 <= _129;
    end
    assign _2206 = 9'b110000000;
    assign _2207 = _1062 == _2206;
    assign _2208 = _1059 & _2207;
    assign _2212 = _2208 ? _515 : _2211;
    assign _2214 = _1047 ? _1055 : _2212;
    assign _130 = _2214;
    always @(posedge _1038) begin
        if (_1036)
            _2211 <= _1055;
        else
            _2211 <= _130;
    end
    assign _2215 = 9'b101111111;
    assign _2216 = _1062 == _2215;
    assign _2217 = _1059 & _2216;
    assign _2221 = _2217 ? _515 : _2220;
    assign _2223 = _1047 ? _1055 : _2221;
    assign _131 = _2223;
    always @(posedge _1038) begin
        if (_1036)
            _2220 <= _1055;
        else
            _2220 <= _131;
    end
    assign _2224 = 9'b101111110;
    assign _2225 = _1062 == _2224;
    assign _2226 = _1059 & _2225;
    assign _2230 = _2226 ? _515 : _2229;
    assign _2232 = _1047 ? _1055 : _2230;
    assign _132 = _2232;
    always @(posedge _1038) begin
        if (_1036)
            _2229 <= _1055;
        else
            _2229 <= _132;
    end
    assign _2233 = 9'b101111101;
    assign _2234 = _1062 == _2233;
    assign _2235 = _1059 & _2234;
    assign _2239 = _2235 ? _515 : _2238;
    assign _2241 = _1047 ? _1055 : _2239;
    assign _133 = _2241;
    always @(posedge _1038) begin
        if (_1036)
            _2238 <= _1055;
        else
            _2238 <= _133;
    end
    assign _2242 = 9'b101111100;
    assign _2243 = _1062 == _2242;
    assign _2244 = _1059 & _2243;
    assign _2248 = _2244 ? _515 : _2247;
    assign _2250 = _1047 ? _1055 : _2248;
    assign _134 = _2250;
    always @(posedge _1038) begin
        if (_1036)
            _2247 <= _1055;
        else
            _2247 <= _134;
    end
    assign _2251 = 9'b101111011;
    assign _2252 = _1062 == _2251;
    assign _2253 = _1059 & _2252;
    assign _2257 = _2253 ? _515 : _2256;
    assign _2259 = _1047 ? _1055 : _2257;
    assign _135 = _2259;
    always @(posedge _1038) begin
        if (_1036)
            _2256 <= _1055;
        else
            _2256 <= _135;
    end
    assign _2260 = 9'b101111010;
    assign _2261 = _1062 == _2260;
    assign _2262 = _1059 & _2261;
    assign _2266 = _2262 ? _515 : _2265;
    assign _2268 = _1047 ? _1055 : _2266;
    assign _136 = _2268;
    always @(posedge _1038) begin
        if (_1036)
            _2265 <= _1055;
        else
            _2265 <= _136;
    end
    assign _2269 = 9'b101111001;
    assign _2270 = _1062 == _2269;
    assign _2271 = _1059 & _2270;
    assign _2275 = _2271 ? _515 : _2274;
    assign _2277 = _1047 ? _1055 : _2275;
    assign _137 = _2277;
    always @(posedge _1038) begin
        if (_1036)
            _2274 <= _1055;
        else
            _2274 <= _137;
    end
    assign _2278 = 9'b101111000;
    assign _2279 = _1062 == _2278;
    assign _2280 = _1059 & _2279;
    assign _2284 = _2280 ? _515 : _2283;
    assign _2286 = _1047 ? _1055 : _2284;
    assign _138 = _2286;
    always @(posedge _1038) begin
        if (_1036)
            _2283 <= _1055;
        else
            _2283 <= _138;
    end
    assign _2287 = 9'b101110111;
    assign _2288 = _1062 == _2287;
    assign _2289 = _1059 & _2288;
    assign _2293 = _2289 ? _515 : _2292;
    assign _2295 = _1047 ? _1055 : _2293;
    assign _139 = _2295;
    always @(posedge _1038) begin
        if (_1036)
            _2292 <= _1055;
        else
            _2292 <= _139;
    end
    assign _2296 = 9'b101110110;
    assign _2297 = _1062 == _2296;
    assign _2298 = _1059 & _2297;
    assign _2302 = _2298 ? _515 : _2301;
    assign _2304 = _1047 ? _1055 : _2302;
    assign _140 = _2304;
    always @(posedge _1038) begin
        if (_1036)
            _2301 <= _1055;
        else
            _2301 <= _140;
    end
    assign _2305 = 9'b101110101;
    assign _2306 = _1062 == _2305;
    assign _2307 = _1059 & _2306;
    assign _2311 = _2307 ? _515 : _2310;
    assign _2313 = _1047 ? _1055 : _2311;
    assign _141 = _2313;
    always @(posedge _1038) begin
        if (_1036)
            _2310 <= _1055;
        else
            _2310 <= _141;
    end
    assign _2314 = 9'b101110100;
    assign _2315 = _1062 == _2314;
    assign _2316 = _1059 & _2315;
    assign _2320 = _2316 ? _515 : _2319;
    assign _2322 = _1047 ? _1055 : _2320;
    assign _142 = _2322;
    always @(posedge _1038) begin
        if (_1036)
            _2319 <= _1055;
        else
            _2319 <= _142;
    end
    assign _2323 = 9'b101110011;
    assign _2324 = _1062 == _2323;
    assign _2325 = _1059 & _2324;
    assign _2329 = _2325 ? _515 : _2328;
    assign _2331 = _1047 ? _1055 : _2329;
    assign _143 = _2331;
    always @(posedge _1038) begin
        if (_1036)
            _2328 <= _1055;
        else
            _2328 <= _143;
    end
    assign _2332 = 9'b101110010;
    assign _2333 = _1062 == _2332;
    assign _2334 = _1059 & _2333;
    assign _2338 = _2334 ? _515 : _2337;
    assign _2340 = _1047 ? _1055 : _2338;
    assign _144 = _2340;
    always @(posedge _1038) begin
        if (_1036)
            _2337 <= _1055;
        else
            _2337 <= _144;
    end
    assign _2341 = 9'b101110001;
    assign _2342 = _1062 == _2341;
    assign _2343 = _1059 & _2342;
    assign _2347 = _2343 ? _515 : _2346;
    assign _2349 = _1047 ? _1055 : _2347;
    assign _145 = _2349;
    always @(posedge _1038) begin
        if (_1036)
            _2346 <= _1055;
        else
            _2346 <= _145;
    end
    assign _2350 = 9'b101110000;
    assign _2351 = _1062 == _2350;
    assign _2352 = _1059 & _2351;
    assign _2356 = _2352 ? _515 : _2355;
    assign _2358 = _1047 ? _1055 : _2356;
    assign _146 = _2358;
    always @(posedge _1038) begin
        if (_1036)
            _2355 <= _1055;
        else
            _2355 <= _146;
    end
    assign _2359 = 9'b101101111;
    assign _2360 = _1062 == _2359;
    assign _2361 = _1059 & _2360;
    assign _2365 = _2361 ? _515 : _2364;
    assign _2367 = _1047 ? _1055 : _2365;
    assign _147 = _2367;
    always @(posedge _1038) begin
        if (_1036)
            _2364 <= _1055;
        else
            _2364 <= _147;
    end
    assign _2368 = 9'b101101110;
    assign _2369 = _1062 == _2368;
    assign _2370 = _1059 & _2369;
    assign _2374 = _2370 ? _515 : _2373;
    assign _2376 = _1047 ? _1055 : _2374;
    assign _148 = _2376;
    always @(posedge _1038) begin
        if (_1036)
            _2373 <= _1055;
        else
            _2373 <= _148;
    end
    assign _2377 = 9'b101101101;
    assign _2378 = _1062 == _2377;
    assign _2379 = _1059 & _2378;
    assign _2383 = _2379 ? _515 : _2382;
    assign _2385 = _1047 ? _1055 : _2383;
    assign _149 = _2385;
    always @(posedge _1038) begin
        if (_1036)
            _2382 <= _1055;
        else
            _2382 <= _149;
    end
    assign _2386 = 9'b101101100;
    assign _2387 = _1062 == _2386;
    assign _2388 = _1059 & _2387;
    assign _2392 = _2388 ? _515 : _2391;
    assign _2394 = _1047 ? _1055 : _2392;
    assign _150 = _2394;
    always @(posedge _1038) begin
        if (_1036)
            _2391 <= _1055;
        else
            _2391 <= _150;
    end
    assign _2395 = 9'b101101011;
    assign _2396 = _1062 == _2395;
    assign _2397 = _1059 & _2396;
    assign _2401 = _2397 ? _515 : _2400;
    assign _2403 = _1047 ? _1055 : _2401;
    assign _151 = _2403;
    always @(posedge _1038) begin
        if (_1036)
            _2400 <= _1055;
        else
            _2400 <= _151;
    end
    assign _2404 = 9'b101101010;
    assign _2405 = _1062 == _2404;
    assign _2406 = _1059 & _2405;
    assign _2410 = _2406 ? _515 : _2409;
    assign _2412 = _1047 ? _1055 : _2410;
    assign _152 = _2412;
    always @(posedge _1038) begin
        if (_1036)
            _2409 <= _1055;
        else
            _2409 <= _152;
    end
    assign _2413 = 9'b101101001;
    assign _2414 = _1062 == _2413;
    assign _2415 = _1059 & _2414;
    assign _2419 = _2415 ? _515 : _2418;
    assign _2421 = _1047 ? _1055 : _2419;
    assign _153 = _2421;
    always @(posedge _1038) begin
        if (_1036)
            _2418 <= _1055;
        else
            _2418 <= _153;
    end
    assign _2422 = 9'b101101000;
    assign _2423 = _1062 == _2422;
    assign _2424 = _1059 & _2423;
    assign _2428 = _2424 ? _515 : _2427;
    assign _2430 = _1047 ? _1055 : _2428;
    assign _154 = _2430;
    always @(posedge _1038) begin
        if (_1036)
            _2427 <= _1055;
        else
            _2427 <= _154;
    end
    assign _2431 = 9'b101100111;
    assign _2432 = _1062 == _2431;
    assign _2433 = _1059 & _2432;
    assign _2437 = _2433 ? _515 : _2436;
    assign _2439 = _1047 ? _1055 : _2437;
    assign _155 = _2439;
    always @(posedge _1038) begin
        if (_1036)
            _2436 <= _1055;
        else
            _2436 <= _155;
    end
    assign _2440 = 9'b101100110;
    assign _2441 = _1062 == _2440;
    assign _2442 = _1059 & _2441;
    assign _2446 = _2442 ? _515 : _2445;
    assign _2448 = _1047 ? _1055 : _2446;
    assign _156 = _2448;
    always @(posedge _1038) begin
        if (_1036)
            _2445 <= _1055;
        else
            _2445 <= _156;
    end
    assign _2449 = 9'b101100101;
    assign _2450 = _1062 == _2449;
    assign _2451 = _1059 & _2450;
    assign _2455 = _2451 ? _515 : _2454;
    assign _2457 = _1047 ? _1055 : _2455;
    assign _157 = _2457;
    always @(posedge _1038) begin
        if (_1036)
            _2454 <= _1055;
        else
            _2454 <= _157;
    end
    assign _2458 = 9'b101100100;
    assign _2459 = _1062 == _2458;
    assign _2460 = _1059 & _2459;
    assign _2464 = _2460 ? _515 : _2463;
    assign _2466 = _1047 ? _1055 : _2464;
    assign _158 = _2466;
    always @(posedge _1038) begin
        if (_1036)
            _2463 <= _1055;
        else
            _2463 <= _158;
    end
    assign _2467 = 9'b101100011;
    assign _2468 = _1062 == _2467;
    assign _2469 = _1059 & _2468;
    assign _2473 = _2469 ? _515 : _2472;
    assign _2475 = _1047 ? _1055 : _2473;
    assign _159 = _2475;
    always @(posedge _1038) begin
        if (_1036)
            _2472 <= _1055;
        else
            _2472 <= _159;
    end
    assign _2476 = 9'b101100010;
    assign _2477 = _1062 == _2476;
    assign _2478 = _1059 & _2477;
    assign _2482 = _2478 ? _515 : _2481;
    assign _2484 = _1047 ? _1055 : _2482;
    assign _160 = _2484;
    always @(posedge _1038) begin
        if (_1036)
            _2481 <= _1055;
        else
            _2481 <= _160;
    end
    assign _2485 = 9'b101100001;
    assign _2486 = _1062 == _2485;
    assign _2487 = _1059 & _2486;
    assign _2491 = _2487 ? _515 : _2490;
    assign _2493 = _1047 ? _1055 : _2491;
    assign _161 = _2493;
    always @(posedge _1038) begin
        if (_1036)
            _2490 <= _1055;
        else
            _2490 <= _161;
    end
    assign _2494 = 9'b101100000;
    assign _2495 = _1062 == _2494;
    assign _2496 = _1059 & _2495;
    assign _2500 = _2496 ? _515 : _2499;
    assign _2502 = _1047 ? _1055 : _2500;
    assign _162 = _2502;
    always @(posedge _1038) begin
        if (_1036)
            _2499 <= _1055;
        else
            _2499 <= _162;
    end
    assign _2503 = 9'b101011111;
    assign _2504 = _1062 == _2503;
    assign _2505 = _1059 & _2504;
    assign _2509 = _2505 ? _515 : _2508;
    assign _2511 = _1047 ? _1055 : _2509;
    assign _163 = _2511;
    always @(posedge _1038) begin
        if (_1036)
            _2508 <= _1055;
        else
            _2508 <= _163;
    end
    assign _2512 = 9'b101011110;
    assign _2513 = _1062 == _2512;
    assign _2514 = _1059 & _2513;
    assign _2518 = _2514 ? _515 : _2517;
    assign _2520 = _1047 ? _1055 : _2518;
    assign _164 = _2520;
    always @(posedge _1038) begin
        if (_1036)
            _2517 <= _1055;
        else
            _2517 <= _164;
    end
    assign _2521 = 9'b101011101;
    assign _2522 = _1062 == _2521;
    assign _2523 = _1059 & _2522;
    assign _2527 = _2523 ? _515 : _2526;
    assign _2529 = _1047 ? _1055 : _2527;
    assign _165 = _2529;
    always @(posedge _1038) begin
        if (_1036)
            _2526 <= _1055;
        else
            _2526 <= _165;
    end
    assign _2530 = 9'b101011100;
    assign _2531 = _1062 == _2530;
    assign _2532 = _1059 & _2531;
    assign _2536 = _2532 ? _515 : _2535;
    assign _2538 = _1047 ? _1055 : _2536;
    assign _166 = _2538;
    always @(posedge _1038) begin
        if (_1036)
            _2535 <= _1055;
        else
            _2535 <= _166;
    end
    assign _2539 = 9'b101011011;
    assign _2540 = _1062 == _2539;
    assign _2541 = _1059 & _2540;
    assign _2545 = _2541 ? _515 : _2544;
    assign _2547 = _1047 ? _1055 : _2545;
    assign _167 = _2547;
    always @(posedge _1038) begin
        if (_1036)
            _2544 <= _1055;
        else
            _2544 <= _167;
    end
    assign _2548 = 9'b101011010;
    assign _2549 = _1062 == _2548;
    assign _2550 = _1059 & _2549;
    assign _2554 = _2550 ? _515 : _2553;
    assign _2556 = _1047 ? _1055 : _2554;
    assign _168 = _2556;
    always @(posedge _1038) begin
        if (_1036)
            _2553 <= _1055;
        else
            _2553 <= _168;
    end
    assign _2557 = 9'b101011001;
    assign _2558 = _1062 == _2557;
    assign _2559 = _1059 & _2558;
    assign _2563 = _2559 ? _515 : _2562;
    assign _2565 = _1047 ? _1055 : _2563;
    assign _169 = _2565;
    always @(posedge _1038) begin
        if (_1036)
            _2562 <= _1055;
        else
            _2562 <= _169;
    end
    assign _2566 = 9'b101011000;
    assign _2567 = _1062 == _2566;
    assign _2568 = _1059 & _2567;
    assign _2572 = _2568 ? _515 : _2571;
    assign _2574 = _1047 ? _1055 : _2572;
    assign _170 = _2574;
    always @(posedge _1038) begin
        if (_1036)
            _2571 <= _1055;
        else
            _2571 <= _170;
    end
    assign _2575 = 9'b101010111;
    assign _2576 = _1062 == _2575;
    assign _2577 = _1059 & _2576;
    assign _2581 = _2577 ? _515 : _2580;
    assign _2583 = _1047 ? _1055 : _2581;
    assign _171 = _2583;
    always @(posedge _1038) begin
        if (_1036)
            _2580 <= _1055;
        else
            _2580 <= _171;
    end
    assign _2584 = 9'b101010110;
    assign _2585 = _1062 == _2584;
    assign _2586 = _1059 & _2585;
    assign _2590 = _2586 ? _515 : _2589;
    assign _2592 = _1047 ? _1055 : _2590;
    assign _172 = _2592;
    always @(posedge _1038) begin
        if (_1036)
            _2589 <= _1055;
        else
            _2589 <= _172;
    end
    assign _2593 = 9'b101010101;
    assign _2594 = _1062 == _2593;
    assign _2595 = _1059 & _2594;
    assign _2599 = _2595 ? _515 : _2598;
    assign _2601 = _1047 ? _1055 : _2599;
    assign _173 = _2601;
    always @(posedge _1038) begin
        if (_1036)
            _2598 <= _1055;
        else
            _2598 <= _173;
    end
    assign _2602 = 9'b101010100;
    assign _2603 = _1062 == _2602;
    assign _2604 = _1059 & _2603;
    assign _2608 = _2604 ? _515 : _2607;
    assign _2610 = _1047 ? _1055 : _2608;
    assign _174 = _2610;
    always @(posedge _1038) begin
        if (_1036)
            _2607 <= _1055;
        else
            _2607 <= _174;
    end
    assign _2611 = 9'b101010011;
    assign _2612 = _1062 == _2611;
    assign _2613 = _1059 & _2612;
    assign _2617 = _2613 ? _515 : _2616;
    assign _2619 = _1047 ? _1055 : _2617;
    assign _175 = _2619;
    always @(posedge _1038) begin
        if (_1036)
            _2616 <= _1055;
        else
            _2616 <= _175;
    end
    assign _2620 = 9'b101010010;
    assign _2621 = _1062 == _2620;
    assign _2622 = _1059 & _2621;
    assign _2626 = _2622 ? _515 : _2625;
    assign _2628 = _1047 ? _1055 : _2626;
    assign _176 = _2628;
    always @(posedge _1038) begin
        if (_1036)
            _2625 <= _1055;
        else
            _2625 <= _176;
    end
    assign _2629 = 9'b101010001;
    assign _2630 = _1062 == _2629;
    assign _2631 = _1059 & _2630;
    assign _2635 = _2631 ? _515 : _2634;
    assign _2637 = _1047 ? _1055 : _2635;
    assign _177 = _2637;
    always @(posedge _1038) begin
        if (_1036)
            _2634 <= _1055;
        else
            _2634 <= _177;
    end
    assign _2638 = 9'b101010000;
    assign _2639 = _1062 == _2638;
    assign _2640 = _1059 & _2639;
    assign _2644 = _2640 ? _515 : _2643;
    assign _2646 = _1047 ? _1055 : _2644;
    assign _178 = _2646;
    always @(posedge _1038) begin
        if (_1036)
            _2643 <= _1055;
        else
            _2643 <= _178;
    end
    assign _2647 = 9'b101001111;
    assign _2648 = _1062 == _2647;
    assign _2649 = _1059 & _2648;
    assign _2653 = _2649 ? _515 : _2652;
    assign _2655 = _1047 ? _1055 : _2653;
    assign _179 = _2655;
    always @(posedge _1038) begin
        if (_1036)
            _2652 <= _1055;
        else
            _2652 <= _179;
    end
    assign _2656 = 9'b101001110;
    assign _2657 = _1062 == _2656;
    assign _2658 = _1059 & _2657;
    assign _2662 = _2658 ? _515 : _2661;
    assign _2664 = _1047 ? _1055 : _2662;
    assign _180 = _2664;
    always @(posedge _1038) begin
        if (_1036)
            _2661 <= _1055;
        else
            _2661 <= _180;
    end
    assign _2665 = 9'b101001101;
    assign _2666 = _1062 == _2665;
    assign _2667 = _1059 & _2666;
    assign _2671 = _2667 ? _515 : _2670;
    assign _2673 = _1047 ? _1055 : _2671;
    assign _181 = _2673;
    always @(posedge _1038) begin
        if (_1036)
            _2670 <= _1055;
        else
            _2670 <= _181;
    end
    assign _2674 = 9'b101001100;
    assign _2675 = _1062 == _2674;
    assign _2676 = _1059 & _2675;
    assign _2680 = _2676 ? _515 : _2679;
    assign _2682 = _1047 ? _1055 : _2680;
    assign _182 = _2682;
    always @(posedge _1038) begin
        if (_1036)
            _2679 <= _1055;
        else
            _2679 <= _182;
    end
    assign _2683 = 9'b101001011;
    assign _2684 = _1062 == _2683;
    assign _2685 = _1059 & _2684;
    assign _2689 = _2685 ? _515 : _2688;
    assign _2691 = _1047 ? _1055 : _2689;
    assign _183 = _2691;
    always @(posedge _1038) begin
        if (_1036)
            _2688 <= _1055;
        else
            _2688 <= _183;
    end
    assign _2692 = 9'b101001010;
    assign _2693 = _1062 == _2692;
    assign _2694 = _1059 & _2693;
    assign _2698 = _2694 ? _515 : _2697;
    assign _2700 = _1047 ? _1055 : _2698;
    assign _184 = _2700;
    always @(posedge _1038) begin
        if (_1036)
            _2697 <= _1055;
        else
            _2697 <= _184;
    end
    assign _2701 = 9'b101001001;
    assign _2702 = _1062 == _2701;
    assign _2703 = _1059 & _2702;
    assign _2707 = _2703 ? _515 : _2706;
    assign _2709 = _1047 ? _1055 : _2707;
    assign _185 = _2709;
    always @(posedge _1038) begin
        if (_1036)
            _2706 <= _1055;
        else
            _2706 <= _185;
    end
    assign _2710 = 9'b101001000;
    assign _2711 = _1062 == _2710;
    assign _2712 = _1059 & _2711;
    assign _2716 = _2712 ? _515 : _2715;
    assign _2718 = _1047 ? _1055 : _2716;
    assign _186 = _2718;
    always @(posedge _1038) begin
        if (_1036)
            _2715 <= _1055;
        else
            _2715 <= _186;
    end
    assign _2719 = 9'b101000111;
    assign _2720 = _1062 == _2719;
    assign _2721 = _1059 & _2720;
    assign _2725 = _2721 ? _515 : _2724;
    assign _2727 = _1047 ? _1055 : _2725;
    assign _187 = _2727;
    always @(posedge _1038) begin
        if (_1036)
            _2724 <= _1055;
        else
            _2724 <= _187;
    end
    assign _2728 = 9'b101000110;
    assign _2729 = _1062 == _2728;
    assign _2730 = _1059 & _2729;
    assign _2734 = _2730 ? _515 : _2733;
    assign _2736 = _1047 ? _1055 : _2734;
    assign _188 = _2736;
    always @(posedge _1038) begin
        if (_1036)
            _2733 <= _1055;
        else
            _2733 <= _188;
    end
    assign _2737 = 9'b101000101;
    assign _2738 = _1062 == _2737;
    assign _2739 = _1059 & _2738;
    assign _2743 = _2739 ? _515 : _2742;
    assign _2745 = _1047 ? _1055 : _2743;
    assign _189 = _2745;
    always @(posedge _1038) begin
        if (_1036)
            _2742 <= _1055;
        else
            _2742 <= _189;
    end
    assign _2746 = 9'b101000100;
    assign _2747 = _1062 == _2746;
    assign _2748 = _1059 & _2747;
    assign _2752 = _2748 ? _515 : _2751;
    assign _2754 = _1047 ? _1055 : _2752;
    assign _190 = _2754;
    always @(posedge _1038) begin
        if (_1036)
            _2751 <= _1055;
        else
            _2751 <= _190;
    end
    assign _2755 = 9'b101000011;
    assign _2756 = _1062 == _2755;
    assign _2757 = _1059 & _2756;
    assign _2761 = _2757 ? _515 : _2760;
    assign _2763 = _1047 ? _1055 : _2761;
    assign _191 = _2763;
    always @(posedge _1038) begin
        if (_1036)
            _2760 <= _1055;
        else
            _2760 <= _191;
    end
    assign _2764 = 9'b101000010;
    assign _2765 = _1062 == _2764;
    assign _2766 = _1059 & _2765;
    assign _2770 = _2766 ? _515 : _2769;
    assign _2772 = _1047 ? _1055 : _2770;
    assign _192 = _2772;
    always @(posedge _1038) begin
        if (_1036)
            _2769 <= _1055;
        else
            _2769 <= _192;
    end
    assign _2773 = 9'b101000001;
    assign _2774 = _1062 == _2773;
    assign _2775 = _1059 & _2774;
    assign _2779 = _2775 ? _515 : _2778;
    assign _2781 = _1047 ? _1055 : _2779;
    assign _193 = _2781;
    always @(posedge _1038) begin
        if (_1036)
            _2778 <= _1055;
        else
            _2778 <= _193;
    end
    assign _2782 = 9'b101000000;
    assign _2783 = _1062 == _2782;
    assign _2784 = _1059 & _2783;
    assign _2788 = _2784 ? _515 : _2787;
    assign _2790 = _1047 ? _1055 : _2788;
    assign _194 = _2790;
    always @(posedge _1038) begin
        if (_1036)
            _2787 <= _1055;
        else
            _2787 <= _194;
    end
    assign _2791 = 9'b100111111;
    assign _2792 = _1062 == _2791;
    assign _2793 = _1059 & _2792;
    assign _2797 = _2793 ? _515 : _2796;
    assign _2799 = _1047 ? _1055 : _2797;
    assign _195 = _2799;
    always @(posedge _1038) begin
        if (_1036)
            _2796 <= _1055;
        else
            _2796 <= _195;
    end
    assign _2800 = 9'b100111110;
    assign _2801 = _1062 == _2800;
    assign _2802 = _1059 & _2801;
    assign _2806 = _2802 ? _515 : _2805;
    assign _2808 = _1047 ? _1055 : _2806;
    assign _196 = _2808;
    always @(posedge _1038) begin
        if (_1036)
            _2805 <= _1055;
        else
            _2805 <= _196;
    end
    assign _2809 = 9'b100111101;
    assign _2810 = _1062 == _2809;
    assign _2811 = _1059 & _2810;
    assign _2815 = _2811 ? _515 : _2814;
    assign _2817 = _1047 ? _1055 : _2815;
    assign _197 = _2817;
    always @(posedge _1038) begin
        if (_1036)
            _2814 <= _1055;
        else
            _2814 <= _197;
    end
    assign _2818 = 9'b100111100;
    assign _2819 = _1062 == _2818;
    assign _2820 = _1059 & _2819;
    assign _2824 = _2820 ? _515 : _2823;
    assign _2826 = _1047 ? _1055 : _2824;
    assign _198 = _2826;
    always @(posedge _1038) begin
        if (_1036)
            _2823 <= _1055;
        else
            _2823 <= _198;
    end
    assign _2827 = 9'b100111011;
    assign _2828 = _1062 == _2827;
    assign _2829 = _1059 & _2828;
    assign _2833 = _2829 ? _515 : _2832;
    assign _2835 = _1047 ? _1055 : _2833;
    assign _199 = _2835;
    always @(posedge _1038) begin
        if (_1036)
            _2832 <= _1055;
        else
            _2832 <= _199;
    end
    assign _2836 = 9'b100111010;
    assign _2837 = _1062 == _2836;
    assign _2838 = _1059 & _2837;
    assign _2842 = _2838 ? _515 : _2841;
    assign _2844 = _1047 ? _1055 : _2842;
    assign _200 = _2844;
    always @(posedge _1038) begin
        if (_1036)
            _2841 <= _1055;
        else
            _2841 <= _200;
    end
    assign _2845 = 9'b100111001;
    assign _2846 = _1062 == _2845;
    assign _2847 = _1059 & _2846;
    assign _2851 = _2847 ? _515 : _2850;
    assign _2853 = _1047 ? _1055 : _2851;
    assign _201 = _2853;
    always @(posedge _1038) begin
        if (_1036)
            _2850 <= _1055;
        else
            _2850 <= _201;
    end
    assign _2854 = 9'b100111000;
    assign _2855 = _1062 == _2854;
    assign _2856 = _1059 & _2855;
    assign _2860 = _2856 ? _515 : _2859;
    assign _2862 = _1047 ? _1055 : _2860;
    assign _202 = _2862;
    always @(posedge _1038) begin
        if (_1036)
            _2859 <= _1055;
        else
            _2859 <= _202;
    end
    assign _2863 = 9'b100110111;
    assign _2864 = _1062 == _2863;
    assign _2865 = _1059 & _2864;
    assign _2869 = _2865 ? _515 : _2868;
    assign _2871 = _1047 ? _1055 : _2869;
    assign _203 = _2871;
    always @(posedge _1038) begin
        if (_1036)
            _2868 <= _1055;
        else
            _2868 <= _203;
    end
    assign _2872 = 9'b100110110;
    assign _2873 = _1062 == _2872;
    assign _2874 = _1059 & _2873;
    assign _2878 = _2874 ? _515 : _2877;
    assign _2880 = _1047 ? _1055 : _2878;
    assign _204 = _2880;
    always @(posedge _1038) begin
        if (_1036)
            _2877 <= _1055;
        else
            _2877 <= _204;
    end
    assign _2881 = 9'b100110101;
    assign _2882 = _1062 == _2881;
    assign _2883 = _1059 & _2882;
    assign _2887 = _2883 ? _515 : _2886;
    assign _2889 = _1047 ? _1055 : _2887;
    assign _205 = _2889;
    always @(posedge _1038) begin
        if (_1036)
            _2886 <= _1055;
        else
            _2886 <= _205;
    end
    assign _2890 = 9'b100110100;
    assign _2891 = _1062 == _2890;
    assign _2892 = _1059 & _2891;
    assign _2896 = _2892 ? _515 : _2895;
    assign _2898 = _1047 ? _1055 : _2896;
    assign _206 = _2898;
    always @(posedge _1038) begin
        if (_1036)
            _2895 <= _1055;
        else
            _2895 <= _206;
    end
    assign _2899 = 9'b100110011;
    assign _2900 = _1062 == _2899;
    assign _2901 = _1059 & _2900;
    assign _2905 = _2901 ? _515 : _2904;
    assign _2907 = _1047 ? _1055 : _2905;
    assign _207 = _2907;
    always @(posedge _1038) begin
        if (_1036)
            _2904 <= _1055;
        else
            _2904 <= _207;
    end
    assign _2908 = 9'b100110010;
    assign _2909 = _1062 == _2908;
    assign _2910 = _1059 & _2909;
    assign _2914 = _2910 ? _515 : _2913;
    assign _2916 = _1047 ? _1055 : _2914;
    assign _208 = _2916;
    always @(posedge _1038) begin
        if (_1036)
            _2913 <= _1055;
        else
            _2913 <= _208;
    end
    assign _2917 = 9'b100110001;
    assign _2918 = _1062 == _2917;
    assign _2919 = _1059 & _2918;
    assign _2923 = _2919 ? _515 : _2922;
    assign _2925 = _1047 ? _1055 : _2923;
    assign _209 = _2925;
    always @(posedge _1038) begin
        if (_1036)
            _2922 <= _1055;
        else
            _2922 <= _209;
    end
    assign _2926 = 9'b100110000;
    assign _2927 = _1062 == _2926;
    assign _2928 = _1059 & _2927;
    assign _2932 = _2928 ? _515 : _2931;
    assign _2934 = _1047 ? _1055 : _2932;
    assign _210 = _2934;
    always @(posedge _1038) begin
        if (_1036)
            _2931 <= _1055;
        else
            _2931 <= _210;
    end
    assign _2935 = 9'b100101111;
    assign _2936 = _1062 == _2935;
    assign _2937 = _1059 & _2936;
    assign _2941 = _2937 ? _515 : _2940;
    assign _2943 = _1047 ? _1055 : _2941;
    assign _211 = _2943;
    always @(posedge _1038) begin
        if (_1036)
            _2940 <= _1055;
        else
            _2940 <= _211;
    end
    assign _2944 = 9'b100101110;
    assign _2945 = _1062 == _2944;
    assign _2946 = _1059 & _2945;
    assign _2950 = _2946 ? _515 : _2949;
    assign _2952 = _1047 ? _1055 : _2950;
    assign _212 = _2952;
    always @(posedge _1038) begin
        if (_1036)
            _2949 <= _1055;
        else
            _2949 <= _212;
    end
    assign _2953 = 9'b100101101;
    assign _2954 = _1062 == _2953;
    assign _2955 = _1059 & _2954;
    assign _2959 = _2955 ? _515 : _2958;
    assign _2961 = _1047 ? _1055 : _2959;
    assign _213 = _2961;
    always @(posedge _1038) begin
        if (_1036)
            _2958 <= _1055;
        else
            _2958 <= _213;
    end
    assign _2962 = 9'b100101100;
    assign _2963 = _1062 == _2962;
    assign _2964 = _1059 & _2963;
    assign _2968 = _2964 ? _515 : _2967;
    assign _2970 = _1047 ? _1055 : _2968;
    assign _214 = _2970;
    always @(posedge _1038) begin
        if (_1036)
            _2967 <= _1055;
        else
            _2967 <= _214;
    end
    assign _2971 = 9'b100101011;
    assign _2972 = _1062 == _2971;
    assign _2973 = _1059 & _2972;
    assign _2977 = _2973 ? _515 : _2976;
    assign _2979 = _1047 ? _1055 : _2977;
    assign _215 = _2979;
    always @(posedge _1038) begin
        if (_1036)
            _2976 <= _1055;
        else
            _2976 <= _215;
    end
    assign _2980 = 9'b100101010;
    assign _2981 = _1062 == _2980;
    assign _2982 = _1059 & _2981;
    assign _2986 = _2982 ? _515 : _2985;
    assign _2988 = _1047 ? _1055 : _2986;
    assign _216 = _2988;
    always @(posedge _1038) begin
        if (_1036)
            _2985 <= _1055;
        else
            _2985 <= _216;
    end
    assign _2989 = 9'b100101001;
    assign _2990 = _1062 == _2989;
    assign _2991 = _1059 & _2990;
    assign _2995 = _2991 ? _515 : _2994;
    assign _2997 = _1047 ? _1055 : _2995;
    assign _217 = _2997;
    always @(posedge _1038) begin
        if (_1036)
            _2994 <= _1055;
        else
            _2994 <= _217;
    end
    assign _2998 = 9'b100101000;
    assign _2999 = _1062 == _2998;
    assign _3000 = _1059 & _2999;
    assign _3004 = _3000 ? _515 : _3003;
    assign _3006 = _1047 ? _1055 : _3004;
    assign _218 = _3006;
    always @(posedge _1038) begin
        if (_1036)
            _3003 <= _1055;
        else
            _3003 <= _218;
    end
    assign _3007 = 9'b100100111;
    assign _3008 = _1062 == _3007;
    assign _3009 = _1059 & _3008;
    assign _3013 = _3009 ? _515 : _3012;
    assign _3015 = _1047 ? _1055 : _3013;
    assign _219 = _3015;
    always @(posedge _1038) begin
        if (_1036)
            _3012 <= _1055;
        else
            _3012 <= _219;
    end
    assign _3016 = 9'b100100110;
    assign _3017 = _1062 == _3016;
    assign _3018 = _1059 & _3017;
    assign _3022 = _3018 ? _515 : _3021;
    assign _3024 = _1047 ? _1055 : _3022;
    assign _220 = _3024;
    always @(posedge _1038) begin
        if (_1036)
            _3021 <= _1055;
        else
            _3021 <= _220;
    end
    assign _3025 = 9'b100100101;
    assign _3026 = _1062 == _3025;
    assign _3027 = _1059 & _3026;
    assign _3031 = _3027 ? _515 : _3030;
    assign _3033 = _1047 ? _1055 : _3031;
    assign _221 = _3033;
    always @(posedge _1038) begin
        if (_1036)
            _3030 <= _1055;
        else
            _3030 <= _221;
    end
    assign _3034 = 9'b100100100;
    assign _3035 = _1062 == _3034;
    assign _3036 = _1059 & _3035;
    assign _3040 = _3036 ? _515 : _3039;
    assign _3042 = _1047 ? _1055 : _3040;
    assign _222 = _3042;
    always @(posedge _1038) begin
        if (_1036)
            _3039 <= _1055;
        else
            _3039 <= _222;
    end
    assign _3043 = 9'b100100011;
    assign _3044 = _1062 == _3043;
    assign _3045 = _1059 & _3044;
    assign _3049 = _3045 ? _515 : _3048;
    assign _3051 = _1047 ? _1055 : _3049;
    assign _223 = _3051;
    always @(posedge _1038) begin
        if (_1036)
            _3048 <= _1055;
        else
            _3048 <= _223;
    end
    assign _3052 = 9'b100100010;
    assign _3053 = _1062 == _3052;
    assign _3054 = _1059 & _3053;
    assign _3058 = _3054 ? _515 : _3057;
    assign _3060 = _1047 ? _1055 : _3058;
    assign _224 = _3060;
    always @(posedge _1038) begin
        if (_1036)
            _3057 <= _1055;
        else
            _3057 <= _224;
    end
    assign _3061 = 9'b100100001;
    assign _3062 = _1062 == _3061;
    assign _3063 = _1059 & _3062;
    assign _3067 = _3063 ? _515 : _3066;
    assign _3069 = _1047 ? _1055 : _3067;
    assign _225 = _3069;
    always @(posedge _1038) begin
        if (_1036)
            _3066 <= _1055;
        else
            _3066 <= _225;
    end
    assign _3070 = 9'b100100000;
    assign _3071 = _1062 == _3070;
    assign _3072 = _1059 & _3071;
    assign _3076 = _3072 ? _515 : _3075;
    assign _3078 = _1047 ? _1055 : _3076;
    assign _226 = _3078;
    always @(posedge _1038) begin
        if (_1036)
            _3075 <= _1055;
        else
            _3075 <= _226;
    end
    assign _3079 = 9'b100011111;
    assign _3080 = _1062 == _3079;
    assign _3081 = _1059 & _3080;
    assign _3085 = _3081 ? _515 : _3084;
    assign _3087 = _1047 ? _1055 : _3085;
    assign _227 = _3087;
    always @(posedge _1038) begin
        if (_1036)
            _3084 <= _1055;
        else
            _3084 <= _227;
    end
    assign _3088 = 9'b100011110;
    assign _3089 = _1062 == _3088;
    assign _3090 = _1059 & _3089;
    assign _3094 = _3090 ? _515 : _3093;
    assign _3096 = _1047 ? _1055 : _3094;
    assign _228 = _3096;
    always @(posedge _1038) begin
        if (_1036)
            _3093 <= _1055;
        else
            _3093 <= _228;
    end
    assign _3097 = 9'b100011101;
    assign _3098 = _1062 == _3097;
    assign _3099 = _1059 & _3098;
    assign _3103 = _3099 ? _515 : _3102;
    assign _3105 = _1047 ? _1055 : _3103;
    assign _229 = _3105;
    always @(posedge _1038) begin
        if (_1036)
            _3102 <= _1055;
        else
            _3102 <= _229;
    end
    assign _3106 = 9'b100011100;
    assign _3107 = _1062 == _3106;
    assign _3108 = _1059 & _3107;
    assign _3112 = _3108 ? _515 : _3111;
    assign _3114 = _1047 ? _1055 : _3112;
    assign _230 = _3114;
    always @(posedge _1038) begin
        if (_1036)
            _3111 <= _1055;
        else
            _3111 <= _230;
    end
    assign _3115 = 9'b100011011;
    assign _3116 = _1062 == _3115;
    assign _3117 = _1059 & _3116;
    assign _3121 = _3117 ? _515 : _3120;
    assign _3123 = _1047 ? _1055 : _3121;
    assign _231 = _3123;
    always @(posedge _1038) begin
        if (_1036)
            _3120 <= _1055;
        else
            _3120 <= _231;
    end
    assign _3124 = 9'b100011010;
    assign _3125 = _1062 == _3124;
    assign _3126 = _1059 & _3125;
    assign _3130 = _3126 ? _515 : _3129;
    assign _3132 = _1047 ? _1055 : _3130;
    assign _232 = _3132;
    always @(posedge _1038) begin
        if (_1036)
            _3129 <= _1055;
        else
            _3129 <= _232;
    end
    assign _3133 = 9'b100011001;
    assign _3134 = _1062 == _3133;
    assign _3135 = _1059 & _3134;
    assign _3139 = _3135 ? _515 : _3138;
    assign _3141 = _1047 ? _1055 : _3139;
    assign _233 = _3141;
    always @(posedge _1038) begin
        if (_1036)
            _3138 <= _1055;
        else
            _3138 <= _233;
    end
    assign _3142 = 9'b100011000;
    assign _3143 = _1062 == _3142;
    assign _3144 = _1059 & _3143;
    assign _3148 = _3144 ? _515 : _3147;
    assign _3150 = _1047 ? _1055 : _3148;
    assign _234 = _3150;
    always @(posedge _1038) begin
        if (_1036)
            _3147 <= _1055;
        else
            _3147 <= _234;
    end
    assign _3151 = 9'b100010111;
    assign _3152 = _1062 == _3151;
    assign _3153 = _1059 & _3152;
    assign _3157 = _3153 ? _515 : _3156;
    assign _3159 = _1047 ? _1055 : _3157;
    assign _235 = _3159;
    always @(posedge _1038) begin
        if (_1036)
            _3156 <= _1055;
        else
            _3156 <= _235;
    end
    assign _3160 = 9'b100010110;
    assign _3161 = _1062 == _3160;
    assign _3162 = _1059 & _3161;
    assign _3166 = _3162 ? _515 : _3165;
    assign _3168 = _1047 ? _1055 : _3166;
    assign _236 = _3168;
    always @(posedge _1038) begin
        if (_1036)
            _3165 <= _1055;
        else
            _3165 <= _236;
    end
    assign _3169 = 9'b100010101;
    assign _3170 = _1062 == _3169;
    assign _3171 = _1059 & _3170;
    assign _3175 = _3171 ? _515 : _3174;
    assign _3177 = _1047 ? _1055 : _3175;
    assign _237 = _3177;
    always @(posedge _1038) begin
        if (_1036)
            _3174 <= _1055;
        else
            _3174 <= _237;
    end
    assign _3178 = 9'b100010100;
    assign _3179 = _1062 == _3178;
    assign _3180 = _1059 & _3179;
    assign _3184 = _3180 ? _515 : _3183;
    assign _3186 = _1047 ? _1055 : _3184;
    assign _238 = _3186;
    always @(posedge _1038) begin
        if (_1036)
            _3183 <= _1055;
        else
            _3183 <= _238;
    end
    assign _3187 = 9'b100010011;
    assign _3188 = _1062 == _3187;
    assign _3189 = _1059 & _3188;
    assign _3193 = _3189 ? _515 : _3192;
    assign _3195 = _1047 ? _1055 : _3193;
    assign _239 = _3195;
    always @(posedge _1038) begin
        if (_1036)
            _3192 <= _1055;
        else
            _3192 <= _239;
    end
    assign _3196 = 9'b100010010;
    assign _3197 = _1062 == _3196;
    assign _3198 = _1059 & _3197;
    assign _3202 = _3198 ? _515 : _3201;
    assign _3204 = _1047 ? _1055 : _3202;
    assign _240 = _3204;
    always @(posedge _1038) begin
        if (_1036)
            _3201 <= _1055;
        else
            _3201 <= _240;
    end
    assign _3205 = 9'b100010001;
    assign _3206 = _1062 == _3205;
    assign _3207 = _1059 & _3206;
    assign _3211 = _3207 ? _515 : _3210;
    assign _3213 = _1047 ? _1055 : _3211;
    assign _241 = _3213;
    always @(posedge _1038) begin
        if (_1036)
            _3210 <= _1055;
        else
            _3210 <= _241;
    end
    assign _3214 = 9'b100010000;
    assign _3215 = _1062 == _3214;
    assign _3216 = _1059 & _3215;
    assign _3220 = _3216 ? _515 : _3219;
    assign _3222 = _1047 ? _1055 : _3220;
    assign _242 = _3222;
    always @(posedge _1038) begin
        if (_1036)
            _3219 <= _1055;
        else
            _3219 <= _242;
    end
    assign _3223 = 9'b100001111;
    assign _3224 = _1062 == _3223;
    assign _3225 = _1059 & _3224;
    assign _3229 = _3225 ? _515 : _3228;
    assign _3231 = _1047 ? _1055 : _3229;
    assign _243 = _3231;
    always @(posedge _1038) begin
        if (_1036)
            _3228 <= _1055;
        else
            _3228 <= _243;
    end
    assign _3232 = 9'b100001110;
    assign _3233 = _1062 == _3232;
    assign _3234 = _1059 & _3233;
    assign _3238 = _3234 ? _515 : _3237;
    assign _3240 = _1047 ? _1055 : _3238;
    assign _244 = _3240;
    always @(posedge _1038) begin
        if (_1036)
            _3237 <= _1055;
        else
            _3237 <= _244;
    end
    assign _3241 = 9'b100001101;
    assign _3242 = _1062 == _3241;
    assign _3243 = _1059 & _3242;
    assign _3247 = _3243 ? _515 : _3246;
    assign _3249 = _1047 ? _1055 : _3247;
    assign _245 = _3249;
    always @(posedge _1038) begin
        if (_1036)
            _3246 <= _1055;
        else
            _3246 <= _245;
    end
    assign _3250 = 9'b100001100;
    assign _3251 = _1062 == _3250;
    assign _3252 = _1059 & _3251;
    assign _3256 = _3252 ? _515 : _3255;
    assign _3258 = _1047 ? _1055 : _3256;
    assign _246 = _3258;
    always @(posedge _1038) begin
        if (_1036)
            _3255 <= _1055;
        else
            _3255 <= _246;
    end
    assign _3259 = 9'b100001011;
    assign _3260 = _1062 == _3259;
    assign _3261 = _1059 & _3260;
    assign _3265 = _3261 ? _515 : _3264;
    assign _3267 = _1047 ? _1055 : _3265;
    assign _247 = _3267;
    always @(posedge _1038) begin
        if (_1036)
            _3264 <= _1055;
        else
            _3264 <= _247;
    end
    assign _3268 = 9'b100001010;
    assign _3269 = _1062 == _3268;
    assign _3270 = _1059 & _3269;
    assign _3274 = _3270 ? _515 : _3273;
    assign _3276 = _1047 ? _1055 : _3274;
    assign _248 = _3276;
    always @(posedge _1038) begin
        if (_1036)
            _3273 <= _1055;
        else
            _3273 <= _248;
    end
    assign _3277 = 9'b100001001;
    assign _3278 = _1062 == _3277;
    assign _3279 = _1059 & _3278;
    assign _3283 = _3279 ? _515 : _3282;
    assign _3285 = _1047 ? _1055 : _3283;
    assign _249 = _3285;
    always @(posedge _1038) begin
        if (_1036)
            _3282 <= _1055;
        else
            _3282 <= _249;
    end
    assign _3286 = 9'b100001000;
    assign _3287 = _1062 == _3286;
    assign _3288 = _1059 & _3287;
    assign _3292 = _3288 ? _515 : _3291;
    assign _3294 = _1047 ? _1055 : _3292;
    assign _250 = _3294;
    always @(posedge _1038) begin
        if (_1036)
            _3291 <= _1055;
        else
            _3291 <= _250;
    end
    assign _3295 = 9'b100000111;
    assign _3296 = _1062 == _3295;
    assign _3297 = _1059 & _3296;
    assign _3301 = _3297 ? _515 : _3300;
    assign _3303 = _1047 ? _1055 : _3301;
    assign _251 = _3303;
    always @(posedge _1038) begin
        if (_1036)
            _3300 <= _1055;
        else
            _3300 <= _251;
    end
    assign _3304 = 9'b100000110;
    assign _3305 = _1062 == _3304;
    assign _3306 = _1059 & _3305;
    assign _3310 = _3306 ? _515 : _3309;
    assign _3312 = _1047 ? _1055 : _3310;
    assign _252 = _3312;
    always @(posedge _1038) begin
        if (_1036)
            _3309 <= _1055;
        else
            _3309 <= _252;
    end
    assign _3313 = 9'b100000101;
    assign _3314 = _1062 == _3313;
    assign _3315 = _1059 & _3314;
    assign _3319 = _3315 ? _515 : _3318;
    assign _3321 = _1047 ? _1055 : _3319;
    assign _253 = _3321;
    always @(posedge _1038) begin
        if (_1036)
            _3318 <= _1055;
        else
            _3318 <= _253;
    end
    assign _3322 = 9'b100000100;
    assign _3323 = _1062 == _3322;
    assign _3324 = _1059 & _3323;
    assign _3328 = _3324 ? _515 : _3327;
    assign _3330 = _1047 ? _1055 : _3328;
    assign _254 = _3330;
    always @(posedge _1038) begin
        if (_1036)
            _3327 <= _1055;
        else
            _3327 <= _254;
    end
    assign _3331 = 9'b100000011;
    assign _3332 = _1062 == _3331;
    assign _3333 = _1059 & _3332;
    assign _3337 = _3333 ? _515 : _3336;
    assign _3339 = _1047 ? _1055 : _3337;
    assign _255 = _3339;
    always @(posedge _1038) begin
        if (_1036)
            _3336 <= _1055;
        else
            _3336 <= _255;
    end
    assign _3340 = 9'b100000010;
    assign _3341 = _1062 == _3340;
    assign _3342 = _1059 & _3341;
    assign _3346 = _3342 ? _515 : _3345;
    assign _3348 = _1047 ? _1055 : _3346;
    assign _256 = _3348;
    always @(posedge _1038) begin
        if (_1036)
            _3345 <= _1055;
        else
            _3345 <= _256;
    end
    assign _3349 = 9'b100000001;
    assign _3350 = _1062 == _3349;
    assign _3351 = _1059 & _3350;
    assign _3355 = _3351 ? _515 : _3354;
    assign _3357 = _1047 ? _1055 : _3355;
    assign _257 = _3357;
    always @(posedge _1038) begin
        if (_1036)
            _3354 <= _1055;
        else
            _3354 <= _257;
    end
    assign _3358 = 9'b100000000;
    assign _3359 = _1062 == _3358;
    assign _3360 = _1059 & _3359;
    assign _3364 = _3360 ? _515 : _3363;
    assign _3366 = _1047 ? _1055 : _3364;
    assign _258 = _3366;
    always @(posedge _1038) begin
        if (_1036)
            _3363 <= _1055;
        else
            _3363 <= _258;
    end
    assign _3367 = 9'b011111111;
    assign _3368 = _1062 == _3367;
    assign _3369 = _1059 & _3368;
    assign _3373 = _3369 ? _515 : _3372;
    assign _3375 = _1047 ? _1055 : _3373;
    assign _259 = _3375;
    always @(posedge _1038) begin
        if (_1036)
            _3372 <= _1055;
        else
            _3372 <= _259;
    end
    assign _3376 = 9'b011111110;
    assign _3377 = _1062 == _3376;
    assign _3378 = _1059 & _3377;
    assign _3382 = _3378 ? _515 : _3381;
    assign _3384 = _1047 ? _1055 : _3382;
    assign _260 = _3384;
    always @(posedge _1038) begin
        if (_1036)
            _3381 <= _1055;
        else
            _3381 <= _260;
    end
    assign _3385 = 9'b011111101;
    assign _3386 = _1062 == _3385;
    assign _3387 = _1059 & _3386;
    assign _3391 = _3387 ? _515 : _3390;
    assign _3393 = _1047 ? _1055 : _3391;
    assign _261 = _3393;
    always @(posedge _1038) begin
        if (_1036)
            _3390 <= _1055;
        else
            _3390 <= _261;
    end
    assign _3394 = 9'b011111100;
    assign _3395 = _1062 == _3394;
    assign _3396 = _1059 & _3395;
    assign _3400 = _3396 ? _515 : _3399;
    assign _3402 = _1047 ? _1055 : _3400;
    assign _262 = _3402;
    always @(posedge _1038) begin
        if (_1036)
            _3399 <= _1055;
        else
            _3399 <= _262;
    end
    assign _3403 = 9'b011111011;
    assign _3404 = _1062 == _3403;
    assign _3405 = _1059 & _3404;
    assign _3409 = _3405 ? _515 : _3408;
    assign _3411 = _1047 ? _1055 : _3409;
    assign _263 = _3411;
    always @(posedge _1038) begin
        if (_1036)
            _3408 <= _1055;
        else
            _3408 <= _263;
    end
    assign _3412 = 9'b011111010;
    assign _3413 = _1062 == _3412;
    assign _3414 = _1059 & _3413;
    assign _3418 = _3414 ? _515 : _3417;
    assign _3420 = _1047 ? _1055 : _3418;
    assign _264 = _3420;
    always @(posedge _1038) begin
        if (_1036)
            _3417 <= _1055;
        else
            _3417 <= _264;
    end
    assign _3421 = 9'b011111001;
    assign _3422 = _1062 == _3421;
    assign _3423 = _1059 & _3422;
    assign _3427 = _3423 ? _515 : _3426;
    assign _3429 = _1047 ? _1055 : _3427;
    assign _265 = _3429;
    always @(posedge _1038) begin
        if (_1036)
            _3426 <= _1055;
        else
            _3426 <= _265;
    end
    assign _3430 = 9'b011111000;
    assign _3431 = _1062 == _3430;
    assign _3432 = _1059 & _3431;
    assign _3436 = _3432 ? _515 : _3435;
    assign _3438 = _1047 ? _1055 : _3436;
    assign _266 = _3438;
    always @(posedge _1038) begin
        if (_1036)
            _3435 <= _1055;
        else
            _3435 <= _266;
    end
    assign _3439 = 9'b011110111;
    assign _3440 = _1062 == _3439;
    assign _3441 = _1059 & _3440;
    assign _3445 = _3441 ? _515 : _3444;
    assign _3447 = _1047 ? _1055 : _3445;
    assign _267 = _3447;
    always @(posedge _1038) begin
        if (_1036)
            _3444 <= _1055;
        else
            _3444 <= _267;
    end
    assign _3448 = 9'b011110110;
    assign _3449 = _1062 == _3448;
    assign _3450 = _1059 & _3449;
    assign _3454 = _3450 ? _515 : _3453;
    assign _3456 = _1047 ? _1055 : _3454;
    assign _268 = _3456;
    always @(posedge _1038) begin
        if (_1036)
            _3453 <= _1055;
        else
            _3453 <= _268;
    end
    assign _3457 = 9'b011110101;
    assign _3458 = _1062 == _3457;
    assign _3459 = _1059 & _3458;
    assign _3463 = _3459 ? _515 : _3462;
    assign _3465 = _1047 ? _1055 : _3463;
    assign _269 = _3465;
    always @(posedge _1038) begin
        if (_1036)
            _3462 <= _1055;
        else
            _3462 <= _269;
    end
    assign _3466 = 9'b011110100;
    assign _3467 = _1062 == _3466;
    assign _3468 = _1059 & _3467;
    assign _3472 = _3468 ? _515 : _3471;
    assign _3474 = _1047 ? _1055 : _3472;
    assign _270 = _3474;
    always @(posedge _1038) begin
        if (_1036)
            _3471 <= _1055;
        else
            _3471 <= _270;
    end
    assign _3475 = 9'b011110011;
    assign _3476 = _1062 == _3475;
    assign _3477 = _1059 & _3476;
    assign _3481 = _3477 ? _515 : _3480;
    assign _3483 = _1047 ? _1055 : _3481;
    assign _271 = _3483;
    always @(posedge _1038) begin
        if (_1036)
            _3480 <= _1055;
        else
            _3480 <= _271;
    end
    assign _3484 = 9'b011110010;
    assign _3485 = _1062 == _3484;
    assign _3486 = _1059 & _3485;
    assign _3490 = _3486 ? _515 : _3489;
    assign _3492 = _1047 ? _1055 : _3490;
    assign _272 = _3492;
    always @(posedge _1038) begin
        if (_1036)
            _3489 <= _1055;
        else
            _3489 <= _272;
    end
    assign _3493 = 9'b011110001;
    assign _3494 = _1062 == _3493;
    assign _3495 = _1059 & _3494;
    assign _3499 = _3495 ? _515 : _3498;
    assign _3501 = _1047 ? _1055 : _3499;
    assign _273 = _3501;
    always @(posedge _1038) begin
        if (_1036)
            _3498 <= _1055;
        else
            _3498 <= _273;
    end
    assign _3502 = 9'b011110000;
    assign _3503 = _1062 == _3502;
    assign _3504 = _1059 & _3503;
    assign _3508 = _3504 ? _515 : _3507;
    assign _3510 = _1047 ? _1055 : _3508;
    assign _274 = _3510;
    always @(posedge _1038) begin
        if (_1036)
            _3507 <= _1055;
        else
            _3507 <= _274;
    end
    assign _3511 = 9'b011101111;
    assign _3512 = _1062 == _3511;
    assign _3513 = _1059 & _3512;
    assign _3517 = _3513 ? _515 : _3516;
    assign _3519 = _1047 ? _1055 : _3517;
    assign _275 = _3519;
    always @(posedge _1038) begin
        if (_1036)
            _3516 <= _1055;
        else
            _3516 <= _275;
    end
    assign _3520 = 9'b011101110;
    assign _3521 = _1062 == _3520;
    assign _3522 = _1059 & _3521;
    assign _3526 = _3522 ? _515 : _3525;
    assign _3528 = _1047 ? _1055 : _3526;
    assign _276 = _3528;
    always @(posedge _1038) begin
        if (_1036)
            _3525 <= _1055;
        else
            _3525 <= _276;
    end
    assign _3529 = 9'b011101101;
    assign _3530 = _1062 == _3529;
    assign _3531 = _1059 & _3530;
    assign _3535 = _3531 ? _515 : _3534;
    assign _3537 = _1047 ? _1055 : _3535;
    assign _277 = _3537;
    always @(posedge _1038) begin
        if (_1036)
            _3534 <= _1055;
        else
            _3534 <= _277;
    end
    assign _3538 = 9'b011101100;
    assign _3539 = _1062 == _3538;
    assign _3540 = _1059 & _3539;
    assign _3544 = _3540 ? _515 : _3543;
    assign _3546 = _1047 ? _1055 : _3544;
    assign _278 = _3546;
    always @(posedge _1038) begin
        if (_1036)
            _3543 <= _1055;
        else
            _3543 <= _278;
    end
    assign _3547 = 9'b011101011;
    assign _3548 = _1062 == _3547;
    assign _3549 = _1059 & _3548;
    assign _3553 = _3549 ? _515 : _3552;
    assign _3555 = _1047 ? _1055 : _3553;
    assign _279 = _3555;
    always @(posedge _1038) begin
        if (_1036)
            _3552 <= _1055;
        else
            _3552 <= _279;
    end
    assign _3556 = 9'b011101010;
    assign _3557 = _1062 == _3556;
    assign _3558 = _1059 & _3557;
    assign _3562 = _3558 ? _515 : _3561;
    assign _3564 = _1047 ? _1055 : _3562;
    assign _280 = _3564;
    always @(posedge _1038) begin
        if (_1036)
            _3561 <= _1055;
        else
            _3561 <= _280;
    end
    assign _3565 = 9'b011101001;
    assign _3566 = _1062 == _3565;
    assign _3567 = _1059 & _3566;
    assign _3571 = _3567 ? _515 : _3570;
    assign _3573 = _1047 ? _1055 : _3571;
    assign _281 = _3573;
    always @(posedge _1038) begin
        if (_1036)
            _3570 <= _1055;
        else
            _3570 <= _281;
    end
    assign _3574 = 9'b011101000;
    assign _3575 = _1062 == _3574;
    assign _3576 = _1059 & _3575;
    assign _3580 = _3576 ? _515 : _3579;
    assign _3582 = _1047 ? _1055 : _3580;
    assign _282 = _3582;
    always @(posedge _1038) begin
        if (_1036)
            _3579 <= _1055;
        else
            _3579 <= _282;
    end
    assign _3583 = 9'b011100111;
    assign _3584 = _1062 == _3583;
    assign _3585 = _1059 & _3584;
    assign _3589 = _3585 ? _515 : _3588;
    assign _3591 = _1047 ? _1055 : _3589;
    assign _283 = _3591;
    always @(posedge _1038) begin
        if (_1036)
            _3588 <= _1055;
        else
            _3588 <= _283;
    end
    assign _3592 = 9'b011100110;
    assign _3593 = _1062 == _3592;
    assign _3594 = _1059 & _3593;
    assign _3598 = _3594 ? _515 : _3597;
    assign _3600 = _1047 ? _1055 : _3598;
    assign _284 = _3600;
    always @(posedge _1038) begin
        if (_1036)
            _3597 <= _1055;
        else
            _3597 <= _284;
    end
    assign _3601 = 9'b011100101;
    assign _3602 = _1062 == _3601;
    assign _3603 = _1059 & _3602;
    assign _3607 = _3603 ? _515 : _3606;
    assign _3609 = _1047 ? _1055 : _3607;
    assign _285 = _3609;
    always @(posedge _1038) begin
        if (_1036)
            _3606 <= _1055;
        else
            _3606 <= _285;
    end
    assign _3610 = 9'b011100100;
    assign _3611 = _1062 == _3610;
    assign _3612 = _1059 & _3611;
    assign _3616 = _3612 ? _515 : _3615;
    assign _3618 = _1047 ? _1055 : _3616;
    assign _286 = _3618;
    always @(posedge _1038) begin
        if (_1036)
            _3615 <= _1055;
        else
            _3615 <= _286;
    end
    assign _3619 = 9'b011100011;
    assign _3620 = _1062 == _3619;
    assign _3621 = _1059 & _3620;
    assign _3625 = _3621 ? _515 : _3624;
    assign _3627 = _1047 ? _1055 : _3625;
    assign _287 = _3627;
    always @(posedge _1038) begin
        if (_1036)
            _3624 <= _1055;
        else
            _3624 <= _287;
    end
    assign _3628 = 9'b011100010;
    assign _3629 = _1062 == _3628;
    assign _3630 = _1059 & _3629;
    assign _3634 = _3630 ? _515 : _3633;
    assign _3636 = _1047 ? _1055 : _3634;
    assign _288 = _3636;
    always @(posedge _1038) begin
        if (_1036)
            _3633 <= _1055;
        else
            _3633 <= _288;
    end
    assign _3637 = 9'b011100001;
    assign _3638 = _1062 == _3637;
    assign _3639 = _1059 & _3638;
    assign _3643 = _3639 ? _515 : _3642;
    assign _3645 = _1047 ? _1055 : _3643;
    assign _289 = _3645;
    always @(posedge _1038) begin
        if (_1036)
            _3642 <= _1055;
        else
            _3642 <= _289;
    end
    assign _3646 = 9'b011100000;
    assign _3647 = _1062 == _3646;
    assign _3648 = _1059 & _3647;
    assign _3652 = _3648 ? _515 : _3651;
    assign _3654 = _1047 ? _1055 : _3652;
    assign _290 = _3654;
    always @(posedge _1038) begin
        if (_1036)
            _3651 <= _1055;
        else
            _3651 <= _290;
    end
    assign _3655 = 9'b011011111;
    assign _3656 = _1062 == _3655;
    assign _3657 = _1059 & _3656;
    assign _3661 = _3657 ? _515 : _3660;
    assign _3663 = _1047 ? _1055 : _3661;
    assign _291 = _3663;
    always @(posedge _1038) begin
        if (_1036)
            _3660 <= _1055;
        else
            _3660 <= _291;
    end
    assign _3664 = 9'b011011110;
    assign _3665 = _1062 == _3664;
    assign _3666 = _1059 & _3665;
    assign _3670 = _3666 ? _515 : _3669;
    assign _3672 = _1047 ? _1055 : _3670;
    assign _292 = _3672;
    always @(posedge _1038) begin
        if (_1036)
            _3669 <= _1055;
        else
            _3669 <= _292;
    end
    assign _3673 = 9'b011011101;
    assign _3674 = _1062 == _3673;
    assign _3675 = _1059 & _3674;
    assign _3679 = _3675 ? _515 : _3678;
    assign _3681 = _1047 ? _1055 : _3679;
    assign _293 = _3681;
    always @(posedge _1038) begin
        if (_1036)
            _3678 <= _1055;
        else
            _3678 <= _293;
    end
    assign _3682 = 9'b011011100;
    assign _3683 = _1062 == _3682;
    assign _3684 = _1059 & _3683;
    assign _3688 = _3684 ? _515 : _3687;
    assign _3690 = _1047 ? _1055 : _3688;
    assign _294 = _3690;
    always @(posedge _1038) begin
        if (_1036)
            _3687 <= _1055;
        else
            _3687 <= _294;
    end
    assign _3691 = 9'b011011011;
    assign _3692 = _1062 == _3691;
    assign _3693 = _1059 & _3692;
    assign _3697 = _3693 ? _515 : _3696;
    assign _3699 = _1047 ? _1055 : _3697;
    assign _295 = _3699;
    always @(posedge _1038) begin
        if (_1036)
            _3696 <= _1055;
        else
            _3696 <= _295;
    end
    assign _3700 = 9'b011011010;
    assign _3701 = _1062 == _3700;
    assign _3702 = _1059 & _3701;
    assign _3706 = _3702 ? _515 : _3705;
    assign _3708 = _1047 ? _1055 : _3706;
    assign _296 = _3708;
    always @(posedge _1038) begin
        if (_1036)
            _3705 <= _1055;
        else
            _3705 <= _296;
    end
    assign _3709 = 9'b011011001;
    assign _3710 = _1062 == _3709;
    assign _3711 = _1059 & _3710;
    assign _3715 = _3711 ? _515 : _3714;
    assign _3717 = _1047 ? _1055 : _3715;
    assign _297 = _3717;
    always @(posedge _1038) begin
        if (_1036)
            _3714 <= _1055;
        else
            _3714 <= _297;
    end
    assign _3718 = 9'b011011000;
    assign _3719 = _1062 == _3718;
    assign _3720 = _1059 & _3719;
    assign _3724 = _3720 ? _515 : _3723;
    assign _3726 = _1047 ? _1055 : _3724;
    assign _298 = _3726;
    always @(posedge _1038) begin
        if (_1036)
            _3723 <= _1055;
        else
            _3723 <= _298;
    end
    assign _3727 = 9'b011010111;
    assign _3728 = _1062 == _3727;
    assign _3729 = _1059 & _3728;
    assign _3733 = _3729 ? _515 : _3732;
    assign _3735 = _1047 ? _1055 : _3733;
    assign _299 = _3735;
    always @(posedge _1038) begin
        if (_1036)
            _3732 <= _1055;
        else
            _3732 <= _299;
    end
    assign _3736 = 9'b011010110;
    assign _3737 = _1062 == _3736;
    assign _3738 = _1059 & _3737;
    assign _3742 = _3738 ? _515 : _3741;
    assign _3744 = _1047 ? _1055 : _3742;
    assign _300 = _3744;
    always @(posedge _1038) begin
        if (_1036)
            _3741 <= _1055;
        else
            _3741 <= _300;
    end
    assign _3745 = 9'b011010101;
    assign _3746 = _1062 == _3745;
    assign _3747 = _1059 & _3746;
    assign _3751 = _3747 ? _515 : _3750;
    assign _3753 = _1047 ? _1055 : _3751;
    assign _301 = _3753;
    always @(posedge _1038) begin
        if (_1036)
            _3750 <= _1055;
        else
            _3750 <= _301;
    end
    assign _3754 = 9'b011010100;
    assign _3755 = _1062 == _3754;
    assign _3756 = _1059 & _3755;
    assign _3760 = _3756 ? _515 : _3759;
    assign _3762 = _1047 ? _1055 : _3760;
    assign _302 = _3762;
    always @(posedge _1038) begin
        if (_1036)
            _3759 <= _1055;
        else
            _3759 <= _302;
    end
    assign _3763 = 9'b011010011;
    assign _3764 = _1062 == _3763;
    assign _3765 = _1059 & _3764;
    assign _3769 = _3765 ? _515 : _3768;
    assign _3771 = _1047 ? _1055 : _3769;
    assign _303 = _3771;
    always @(posedge _1038) begin
        if (_1036)
            _3768 <= _1055;
        else
            _3768 <= _303;
    end
    assign _3772 = 9'b011010010;
    assign _3773 = _1062 == _3772;
    assign _3774 = _1059 & _3773;
    assign _3778 = _3774 ? _515 : _3777;
    assign _3780 = _1047 ? _1055 : _3778;
    assign _304 = _3780;
    always @(posedge _1038) begin
        if (_1036)
            _3777 <= _1055;
        else
            _3777 <= _304;
    end
    assign _3781 = 9'b011010001;
    assign _3782 = _1062 == _3781;
    assign _3783 = _1059 & _3782;
    assign _3787 = _3783 ? _515 : _3786;
    assign _3789 = _1047 ? _1055 : _3787;
    assign _305 = _3789;
    always @(posedge _1038) begin
        if (_1036)
            _3786 <= _1055;
        else
            _3786 <= _305;
    end
    assign _3790 = 9'b011010000;
    assign _3791 = _1062 == _3790;
    assign _3792 = _1059 & _3791;
    assign _3796 = _3792 ? _515 : _3795;
    assign _3798 = _1047 ? _1055 : _3796;
    assign _306 = _3798;
    always @(posedge _1038) begin
        if (_1036)
            _3795 <= _1055;
        else
            _3795 <= _306;
    end
    assign _3799 = 9'b011001111;
    assign _3800 = _1062 == _3799;
    assign _3801 = _1059 & _3800;
    assign _3805 = _3801 ? _515 : _3804;
    assign _3807 = _1047 ? _1055 : _3805;
    assign _307 = _3807;
    always @(posedge _1038) begin
        if (_1036)
            _3804 <= _1055;
        else
            _3804 <= _307;
    end
    assign _3808 = 9'b011001110;
    assign _3809 = _1062 == _3808;
    assign _3810 = _1059 & _3809;
    assign _3814 = _3810 ? _515 : _3813;
    assign _3816 = _1047 ? _1055 : _3814;
    assign _308 = _3816;
    always @(posedge _1038) begin
        if (_1036)
            _3813 <= _1055;
        else
            _3813 <= _308;
    end
    assign _3817 = 9'b011001101;
    assign _3818 = _1062 == _3817;
    assign _3819 = _1059 & _3818;
    assign _3823 = _3819 ? _515 : _3822;
    assign _3825 = _1047 ? _1055 : _3823;
    assign _309 = _3825;
    always @(posedge _1038) begin
        if (_1036)
            _3822 <= _1055;
        else
            _3822 <= _309;
    end
    assign _3826 = 9'b011001100;
    assign _3827 = _1062 == _3826;
    assign _3828 = _1059 & _3827;
    assign _3832 = _3828 ? _515 : _3831;
    assign _3834 = _1047 ? _1055 : _3832;
    assign _310 = _3834;
    always @(posedge _1038) begin
        if (_1036)
            _3831 <= _1055;
        else
            _3831 <= _310;
    end
    assign _3835 = 9'b011001011;
    assign _3836 = _1062 == _3835;
    assign _3837 = _1059 & _3836;
    assign _3841 = _3837 ? _515 : _3840;
    assign _3843 = _1047 ? _1055 : _3841;
    assign _311 = _3843;
    always @(posedge _1038) begin
        if (_1036)
            _3840 <= _1055;
        else
            _3840 <= _311;
    end
    assign _3844 = 9'b011001010;
    assign _3845 = _1062 == _3844;
    assign _3846 = _1059 & _3845;
    assign _3850 = _3846 ? _515 : _3849;
    assign _3852 = _1047 ? _1055 : _3850;
    assign _312 = _3852;
    always @(posedge _1038) begin
        if (_1036)
            _3849 <= _1055;
        else
            _3849 <= _312;
    end
    assign _3853 = 9'b011001001;
    assign _3854 = _1062 == _3853;
    assign _3855 = _1059 & _3854;
    assign _3859 = _3855 ? _515 : _3858;
    assign _3861 = _1047 ? _1055 : _3859;
    assign _313 = _3861;
    always @(posedge _1038) begin
        if (_1036)
            _3858 <= _1055;
        else
            _3858 <= _313;
    end
    assign _3862 = 9'b011001000;
    assign _3863 = _1062 == _3862;
    assign _3864 = _1059 & _3863;
    assign _3868 = _3864 ? _515 : _3867;
    assign _3870 = _1047 ? _1055 : _3868;
    assign _314 = _3870;
    always @(posedge _1038) begin
        if (_1036)
            _3867 <= _1055;
        else
            _3867 <= _314;
    end
    assign _3871 = 9'b011000111;
    assign _3872 = _1062 == _3871;
    assign _3873 = _1059 & _3872;
    assign _3877 = _3873 ? _515 : _3876;
    assign _3879 = _1047 ? _1055 : _3877;
    assign _315 = _3879;
    always @(posedge _1038) begin
        if (_1036)
            _3876 <= _1055;
        else
            _3876 <= _315;
    end
    assign _3880 = 9'b011000110;
    assign _3881 = _1062 == _3880;
    assign _3882 = _1059 & _3881;
    assign _3886 = _3882 ? _515 : _3885;
    assign _3888 = _1047 ? _1055 : _3886;
    assign _316 = _3888;
    always @(posedge _1038) begin
        if (_1036)
            _3885 <= _1055;
        else
            _3885 <= _316;
    end
    assign _3889 = 9'b011000101;
    assign _3890 = _1062 == _3889;
    assign _3891 = _1059 & _3890;
    assign _3895 = _3891 ? _515 : _3894;
    assign _3897 = _1047 ? _1055 : _3895;
    assign _317 = _3897;
    always @(posedge _1038) begin
        if (_1036)
            _3894 <= _1055;
        else
            _3894 <= _317;
    end
    assign _3898 = 9'b011000100;
    assign _3899 = _1062 == _3898;
    assign _3900 = _1059 & _3899;
    assign _3904 = _3900 ? _515 : _3903;
    assign _3906 = _1047 ? _1055 : _3904;
    assign _318 = _3906;
    always @(posedge _1038) begin
        if (_1036)
            _3903 <= _1055;
        else
            _3903 <= _318;
    end
    assign _3907 = 9'b011000011;
    assign _3908 = _1062 == _3907;
    assign _3909 = _1059 & _3908;
    assign _3913 = _3909 ? _515 : _3912;
    assign _3915 = _1047 ? _1055 : _3913;
    assign _319 = _3915;
    always @(posedge _1038) begin
        if (_1036)
            _3912 <= _1055;
        else
            _3912 <= _319;
    end
    assign _3916 = 9'b011000010;
    assign _3917 = _1062 == _3916;
    assign _3918 = _1059 & _3917;
    assign _3922 = _3918 ? _515 : _3921;
    assign _3924 = _1047 ? _1055 : _3922;
    assign _320 = _3924;
    always @(posedge _1038) begin
        if (_1036)
            _3921 <= _1055;
        else
            _3921 <= _320;
    end
    assign _3925 = 9'b011000001;
    assign _3926 = _1062 == _3925;
    assign _3927 = _1059 & _3926;
    assign _3931 = _3927 ? _515 : _3930;
    assign _3933 = _1047 ? _1055 : _3931;
    assign _321 = _3933;
    always @(posedge _1038) begin
        if (_1036)
            _3930 <= _1055;
        else
            _3930 <= _321;
    end
    assign _3934 = 9'b011000000;
    assign _3935 = _1062 == _3934;
    assign _3936 = _1059 & _3935;
    assign _3940 = _3936 ? _515 : _3939;
    assign _3942 = _1047 ? _1055 : _3940;
    assign _322 = _3942;
    always @(posedge _1038) begin
        if (_1036)
            _3939 <= _1055;
        else
            _3939 <= _322;
    end
    assign _3943 = 9'b010111111;
    assign _3944 = _1062 == _3943;
    assign _3945 = _1059 & _3944;
    assign _3949 = _3945 ? _515 : _3948;
    assign _3951 = _1047 ? _1055 : _3949;
    assign _323 = _3951;
    always @(posedge _1038) begin
        if (_1036)
            _3948 <= _1055;
        else
            _3948 <= _323;
    end
    assign _3952 = 9'b010111110;
    assign _3953 = _1062 == _3952;
    assign _3954 = _1059 & _3953;
    assign _3958 = _3954 ? _515 : _3957;
    assign _3960 = _1047 ? _1055 : _3958;
    assign _324 = _3960;
    always @(posedge _1038) begin
        if (_1036)
            _3957 <= _1055;
        else
            _3957 <= _324;
    end
    assign _3961 = 9'b010111101;
    assign _3962 = _1062 == _3961;
    assign _3963 = _1059 & _3962;
    assign _3967 = _3963 ? _515 : _3966;
    assign _3969 = _1047 ? _1055 : _3967;
    assign _325 = _3969;
    always @(posedge _1038) begin
        if (_1036)
            _3966 <= _1055;
        else
            _3966 <= _325;
    end
    assign _3970 = 9'b010111100;
    assign _3971 = _1062 == _3970;
    assign _3972 = _1059 & _3971;
    assign _3976 = _3972 ? _515 : _3975;
    assign _3978 = _1047 ? _1055 : _3976;
    assign _326 = _3978;
    always @(posedge _1038) begin
        if (_1036)
            _3975 <= _1055;
        else
            _3975 <= _326;
    end
    assign _3979 = 9'b010111011;
    assign _3980 = _1062 == _3979;
    assign _3981 = _1059 & _3980;
    assign _3985 = _3981 ? _515 : _3984;
    assign _3987 = _1047 ? _1055 : _3985;
    assign _327 = _3987;
    always @(posedge _1038) begin
        if (_1036)
            _3984 <= _1055;
        else
            _3984 <= _327;
    end
    assign _3988 = 9'b010111010;
    assign _3989 = _1062 == _3988;
    assign _3990 = _1059 & _3989;
    assign _3994 = _3990 ? _515 : _3993;
    assign _3996 = _1047 ? _1055 : _3994;
    assign _328 = _3996;
    always @(posedge _1038) begin
        if (_1036)
            _3993 <= _1055;
        else
            _3993 <= _328;
    end
    assign _3997 = 9'b010111001;
    assign _3998 = _1062 == _3997;
    assign _3999 = _1059 & _3998;
    assign _4003 = _3999 ? _515 : _4002;
    assign _4005 = _1047 ? _1055 : _4003;
    assign _329 = _4005;
    always @(posedge _1038) begin
        if (_1036)
            _4002 <= _1055;
        else
            _4002 <= _329;
    end
    assign _4006 = 9'b010111000;
    assign _4007 = _1062 == _4006;
    assign _4008 = _1059 & _4007;
    assign _4012 = _4008 ? _515 : _4011;
    assign _4014 = _1047 ? _1055 : _4012;
    assign _330 = _4014;
    always @(posedge _1038) begin
        if (_1036)
            _4011 <= _1055;
        else
            _4011 <= _330;
    end
    assign _4015 = 9'b010110111;
    assign _4016 = _1062 == _4015;
    assign _4017 = _1059 & _4016;
    assign _4021 = _4017 ? _515 : _4020;
    assign _4023 = _1047 ? _1055 : _4021;
    assign _331 = _4023;
    always @(posedge _1038) begin
        if (_1036)
            _4020 <= _1055;
        else
            _4020 <= _331;
    end
    assign _4024 = 9'b010110110;
    assign _4025 = _1062 == _4024;
    assign _4026 = _1059 & _4025;
    assign _4030 = _4026 ? _515 : _4029;
    assign _4032 = _1047 ? _1055 : _4030;
    assign _332 = _4032;
    always @(posedge _1038) begin
        if (_1036)
            _4029 <= _1055;
        else
            _4029 <= _332;
    end
    assign _4033 = 9'b010110101;
    assign _4034 = _1062 == _4033;
    assign _4035 = _1059 & _4034;
    assign _4039 = _4035 ? _515 : _4038;
    assign _4041 = _1047 ? _1055 : _4039;
    assign _333 = _4041;
    always @(posedge _1038) begin
        if (_1036)
            _4038 <= _1055;
        else
            _4038 <= _333;
    end
    assign _4042 = 9'b010110100;
    assign _4043 = _1062 == _4042;
    assign _4044 = _1059 & _4043;
    assign _4048 = _4044 ? _515 : _4047;
    assign _4050 = _1047 ? _1055 : _4048;
    assign _334 = _4050;
    always @(posedge _1038) begin
        if (_1036)
            _4047 <= _1055;
        else
            _4047 <= _334;
    end
    assign _4051 = 9'b010110011;
    assign _4052 = _1062 == _4051;
    assign _4053 = _1059 & _4052;
    assign _4057 = _4053 ? _515 : _4056;
    assign _4059 = _1047 ? _1055 : _4057;
    assign _335 = _4059;
    always @(posedge _1038) begin
        if (_1036)
            _4056 <= _1055;
        else
            _4056 <= _335;
    end
    assign _4060 = 9'b010110010;
    assign _4061 = _1062 == _4060;
    assign _4062 = _1059 & _4061;
    assign _4066 = _4062 ? _515 : _4065;
    assign _4068 = _1047 ? _1055 : _4066;
    assign _336 = _4068;
    always @(posedge _1038) begin
        if (_1036)
            _4065 <= _1055;
        else
            _4065 <= _336;
    end
    assign _4069 = 9'b010110001;
    assign _4070 = _1062 == _4069;
    assign _4071 = _1059 & _4070;
    assign _4075 = _4071 ? _515 : _4074;
    assign _4077 = _1047 ? _1055 : _4075;
    assign _337 = _4077;
    always @(posedge _1038) begin
        if (_1036)
            _4074 <= _1055;
        else
            _4074 <= _337;
    end
    assign _4078 = 9'b010110000;
    assign _4079 = _1062 == _4078;
    assign _4080 = _1059 & _4079;
    assign _4084 = _4080 ? _515 : _4083;
    assign _4086 = _1047 ? _1055 : _4084;
    assign _338 = _4086;
    always @(posedge _1038) begin
        if (_1036)
            _4083 <= _1055;
        else
            _4083 <= _338;
    end
    assign _4087 = 9'b010101111;
    assign _4088 = _1062 == _4087;
    assign _4089 = _1059 & _4088;
    assign _4093 = _4089 ? _515 : _4092;
    assign _4095 = _1047 ? _1055 : _4093;
    assign _339 = _4095;
    always @(posedge _1038) begin
        if (_1036)
            _4092 <= _1055;
        else
            _4092 <= _339;
    end
    assign _4096 = 9'b010101110;
    assign _4097 = _1062 == _4096;
    assign _4098 = _1059 & _4097;
    assign _4102 = _4098 ? _515 : _4101;
    assign _4104 = _1047 ? _1055 : _4102;
    assign _340 = _4104;
    always @(posedge _1038) begin
        if (_1036)
            _4101 <= _1055;
        else
            _4101 <= _340;
    end
    assign _4105 = 9'b010101101;
    assign _4106 = _1062 == _4105;
    assign _4107 = _1059 & _4106;
    assign _4111 = _4107 ? _515 : _4110;
    assign _4113 = _1047 ? _1055 : _4111;
    assign _341 = _4113;
    always @(posedge _1038) begin
        if (_1036)
            _4110 <= _1055;
        else
            _4110 <= _341;
    end
    assign _4114 = 9'b010101100;
    assign _4115 = _1062 == _4114;
    assign _4116 = _1059 & _4115;
    assign _4120 = _4116 ? _515 : _4119;
    assign _4122 = _1047 ? _1055 : _4120;
    assign _342 = _4122;
    always @(posedge _1038) begin
        if (_1036)
            _4119 <= _1055;
        else
            _4119 <= _342;
    end
    assign _4123 = 9'b010101011;
    assign _4124 = _1062 == _4123;
    assign _4125 = _1059 & _4124;
    assign _4129 = _4125 ? _515 : _4128;
    assign _4131 = _1047 ? _1055 : _4129;
    assign _343 = _4131;
    always @(posedge _1038) begin
        if (_1036)
            _4128 <= _1055;
        else
            _4128 <= _343;
    end
    assign _4132 = 9'b010101010;
    assign _4133 = _1062 == _4132;
    assign _4134 = _1059 & _4133;
    assign _4138 = _4134 ? _515 : _4137;
    assign _4140 = _1047 ? _1055 : _4138;
    assign _344 = _4140;
    always @(posedge _1038) begin
        if (_1036)
            _4137 <= _1055;
        else
            _4137 <= _344;
    end
    assign _4141 = 9'b010101001;
    assign _4142 = _1062 == _4141;
    assign _4143 = _1059 & _4142;
    assign _4147 = _4143 ? _515 : _4146;
    assign _4149 = _1047 ? _1055 : _4147;
    assign _345 = _4149;
    always @(posedge _1038) begin
        if (_1036)
            _4146 <= _1055;
        else
            _4146 <= _345;
    end
    assign _4150 = 9'b010101000;
    assign _4151 = _1062 == _4150;
    assign _4152 = _1059 & _4151;
    assign _4156 = _4152 ? _515 : _4155;
    assign _4158 = _1047 ? _1055 : _4156;
    assign _346 = _4158;
    always @(posedge _1038) begin
        if (_1036)
            _4155 <= _1055;
        else
            _4155 <= _346;
    end
    assign _4159 = 9'b010100111;
    assign _4160 = _1062 == _4159;
    assign _4161 = _1059 & _4160;
    assign _4165 = _4161 ? _515 : _4164;
    assign _4167 = _1047 ? _1055 : _4165;
    assign _347 = _4167;
    always @(posedge _1038) begin
        if (_1036)
            _4164 <= _1055;
        else
            _4164 <= _347;
    end
    assign _4168 = 9'b010100110;
    assign _4169 = _1062 == _4168;
    assign _4170 = _1059 & _4169;
    assign _4174 = _4170 ? _515 : _4173;
    assign _4176 = _1047 ? _1055 : _4174;
    assign _348 = _4176;
    always @(posedge _1038) begin
        if (_1036)
            _4173 <= _1055;
        else
            _4173 <= _348;
    end
    assign _4177 = 9'b010100101;
    assign _4178 = _1062 == _4177;
    assign _4179 = _1059 & _4178;
    assign _4183 = _4179 ? _515 : _4182;
    assign _4185 = _1047 ? _1055 : _4183;
    assign _349 = _4185;
    always @(posedge _1038) begin
        if (_1036)
            _4182 <= _1055;
        else
            _4182 <= _349;
    end
    assign _4186 = 9'b010100100;
    assign _4187 = _1062 == _4186;
    assign _4188 = _1059 & _4187;
    assign _4192 = _4188 ? _515 : _4191;
    assign _4194 = _1047 ? _1055 : _4192;
    assign _350 = _4194;
    always @(posedge _1038) begin
        if (_1036)
            _4191 <= _1055;
        else
            _4191 <= _350;
    end
    assign _4195 = 9'b010100011;
    assign _4196 = _1062 == _4195;
    assign _4197 = _1059 & _4196;
    assign _4201 = _4197 ? _515 : _4200;
    assign _4203 = _1047 ? _1055 : _4201;
    assign _351 = _4203;
    always @(posedge _1038) begin
        if (_1036)
            _4200 <= _1055;
        else
            _4200 <= _351;
    end
    assign _4204 = 9'b010100010;
    assign _4205 = _1062 == _4204;
    assign _4206 = _1059 & _4205;
    assign _4210 = _4206 ? _515 : _4209;
    assign _4212 = _1047 ? _1055 : _4210;
    assign _352 = _4212;
    always @(posedge _1038) begin
        if (_1036)
            _4209 <= _1055;
        else
            _4209 <= _352;
    end
    assign _4213 = 9'b010100001;
    assign _4214 = _1062 == _4213;
    assign _4215 = _1059 & _4214;
    assign _4219 = _4215 ? _515 : _4218;
    assign _4221 = _1047 ? _1055 : _4219;
    assign _353 = _4221;
    always @(posedge _1038) begin
        if (_1036)
            _4218 <= _1055;
        else
            _4218 <= _353;
    end
    assign _4222 = 9'b010100000;
    assign _4223 = _1062 == _4222;
    assign _4224 = _1059 & _4223;
    assign _4228 = _4224 ? _515 : _4227;
    assign _4230 = _1047 ? _1055 : _4228;
    assign _354 = _4230;
    always @(posedge _1038) begin
        if (_1036)
            _4227 <= _1055;
        else
            _4227 <= _354;
    end
    assign _4231 = 9'b010011111;
    assign _4232 = _1062 == _4231;
    assign _4233 = _1059 & _4232;
    assign _4237 = _4233 ? _515 : _4236;
    assign _4239 = _1047 ? _1055 : _4237;
    assign _355 = _4239;
    always @(posedge _1038) begin
        if (_1036)
            _4236 <= _1055;
        else
            _4236 <= _355;
    end
    assign _4240 = 9'b010011110;
    assign _4241 = _1062 == _4240;
    assign _4242 = _1059 & _4241;
    assign _4246 = _4242 ? _515 : _4245;
    assign _4248 = _1047 ? _1055 : _4246;
    assign _356 = _4248;
    always @(posedge _1038) begin
        if (_1036)
            _4245 <= _1055;
        else
            _4245 <= _356;
    end
    assign _4249 = 9'b010011101;
    assign _4250 = _1062 == _4249;
    assign _4251 = _1059 & _4250;
    assign _4255 = _4251 ? _515 : _4254;
    assign _4257 = _1047 ? _1055 : _4255;
    assign _357 = _4257;
    always @(posedge _1038) begin
        if (_1036)
            _4254 <= _1055;
        else
            _4254 <= _357;
    end
    assign _4258 = 9'b010011100;
    assign _4259 = _1062 == _4258;
    assign _4260 = _1059 & _4259;
    assign _4264 = _4260 ? _515 : _4263;
    assign _4266 = _1047 ? _1055 : _4264;
    assign _358 = _4266;
    always @(posedge _1038) begin
        if (_1036)
            _4263 <= _1055;
        else
            _4263 <= _358;
    end
    assign _4267 = 9'b010011011;
    assign _4268 = _1062 == _4267;
    assign _4269 = _1059 & _4268;
    assign _4273 = _4269 ? _515 : _4272;
    assign _4275 = _1047 ? _1055 : _4273;
    assign _359 = _4275;
    always @(posedge _1038) begin
        if (_1036)
            _4272 <= _1055;
        else
            _4272 <= _359;
    end
    assign _4276 = 9'b010011010;
    assign _4277 = _1062 == _4276;
    assign _4278 = _1059 & _4277;
    assign _4282 = _4278 ? _515 : _4281;
    assign _4284 = _1047 ? _1055 : _4282;
    assign _360 = _4284;
    always @(posedge _1038) begin
        if (_1036)
            _4281 <= _1055;
        else
            _4281 <= _360;
    end
    assign _4285 = 9'b010011001;
    assign _4286 = _1062 == _4285;
    assign _4287 = _1059 & _4286;
    assign _4291 = _4287 ? _515 : _4290;
    assign _4293 = _1047 ? _1055 : _4291;
    assign _361 = _4293;
    always @(posedge _1038) begin
        if (_1036)
            _4290 <= _1055;
        else
            _4290 <= _361;
    end
    assign _4294 = 9'b010011000;
    assign _4295 = _1062 == _4294;
    assign _4296 = _1059 & _4295;
    assign _4300 = _4296 ? _515 : _4299;
    assign _4302 = _1047 ? _1055 : _4300;
    assign _362 = _4302;
    always @(posedge _1038) begin
        if (_1036)
            _4299 <= _1055;
        else
            _4299 <= _362;
    end
    assign _4303 = 9'b010010111;
    assign _4304 = _1062 == _4303;
    assign _4305 = _1059 & _4304;
    assign _4309 = _4305 ? _515 : _4308;
    assign _4311 = _1047 ? _1055 : _4309;
    assign _363 = _4311;
    always @(posedge _1038) begin
        if (_1036)
            _4308 <= _1055;
        else
            _4308 <= _363;
    end
    assign _4312 = 9'b010010110;
    assign _4313 = _1062 == _4312;
    assign _4314 = _1059 & _4313;
    assign _4318 = _4314 ? _515 : _4317;
    assign _4320 = _1047 ? _1055 : _4318;
    assign _364 = _4320;
    always @(posedge _1038) begin
        if (_1036)
            _4317 <= _1055;
        else
            _4317 <= _364;
    end
    assign _4321 = 9'b010010101;
    assign _4322 = _1062 == _4321;
    assign _4323 = _1059 & _4322;
    assign _4327 = _4323 ? _515 : _4326;
    assign _4329 = _1047 ? _1055 : _4327;
    assign _365 = _4329;
    always @(posedge _1038) begin
        if (_1036)
            _4326 <= _1055;
        else
            _4326 <= _365;
    end
    assign _4330 = 9'b010010100;
    assign _4331 = _1062 == _4330;
    assign _4332 = _1059 & _4331;
    assign _4336 = _4332 ? _515 : _4335;
    assign _4338 = _1047 ? _1055 : _4336;
    assign _366 = _4338;
    always @(posedge _1038) begin
        if (_1036)
            _4335 <= _1055;
        else
            _4335 <= _366;
    end
    assign _4339 = 9'b010010011;
    assign _4340 = _1062 == _4339;
    assign _4341 = _1059 & _4340;
    assign _4345 = _4341 ? _515 : _4344;
    assign _4347 = _1047 ? _1055 : _4345;
    assign _367 = _4347;
    always @(posedge _1038) begin
        if (_1036)
            _4344 <= _1055;
        else
            _4344 <= _367;
    end
    assign _4348 = 9'b010010010;
    assign _4349 = _1062 == _4348;
    assign _4350 = _1059 & _4349;
    assign _4354 = _4350 ? _515 : _4353;
    assign _4356 = _1047 ? _1055 : _4354;
    assign _368 = _4356;
    always @(posedge _1038) begin
        if (_1036)
            _4353 <= _1055;
        else
            _4353 <= _368;
    end
    assign _4357 = 9'b010010001;
    assign _4358 = _1062 == _4357;
    assign _4359 = _1059 & _4358;
    assign _4363 = _4359 ? _515 : _4362;
    assign _4365 = _1047 ? _1055 : _4363;
    assign _369 = _4365;
    always @(posedge _1038) begin
        if (_1036)
            _4362 <= _1055;
        else
            _4362 <= _369;
    end
    assign _4366 = 9'b010010000;
    assign _4367 = _1062 == _4366;
    assign _4368 = _1059 & _4367;
    assign _4372 = _4368 ? _515 : _4371;
    assign _4374 = _1047 ? _1055 : _4372;
    assign _370 = _4374;
    always @(posedge _1038) begin
        if (_1036)
            _4371 <= _1055;
        else
            _4371 <= _370;
    end
    assign _4375 = 9'b010001111;
    assign _4376 = _1062 == _4375;
    assign _4377 = _1059 & _4376;
    assign _4381 = _4377 ? _515 : _4380;
    assign _4383 = _1047 ? _1055 : _4381;
    assign _371 = _4383;
    always @(posedge _1038) begin
        if (_1036)
            _4380 <= _1055;
        else
            _4380 <= _371;
    end
    assign _4384 = 9'b010001110;
    assign _4385 = _1062 == _4384;
    assign _4386 = _1059 & _4385;
    assign _4390 = _4386 ? _515 : _4389;
    assign _4392 = _1047 ? _1055 : _4390;
    assign _372 = _4392;
    always @(posedge _1038) begin
        if (_1036)
            _4389 <= _1055;
        else
            _4389 <= _372;
    end
    assign _4393 = 9'b010001101;
    assign _4394 = _1062 == _4393;
    assign _4395 = _1059 & _4394;
    assign _4399 = _4395 ? _515 : _4398;
    assign _4401 = _1047 ? _1055 : _4399;
    assign _373 = _4401;
    always @(posedge _1038) begin
        if (_1036)
            _4398 <= _1055;
        else
            _4398 <= _373;
    end
    assign _4402 = 9'b010001100;
    assign _4403 = _1062 == _4402;
    assign _4404 = _1059 & _4403;
    assign _4408 = _4404 ? _515 : _4407;
    assign _4410 = _1047 ? _1055 : _4408;
    assign _374 = _4410;
    always @(posedge _1038) begin
        if (_1036)
            _4407 <= _1055;
        else
            _4407 <= _374;
    end
    assign _4411 = 9'b010001011;
    assign _4412 = _1062 == _4411;
    assign _4413 = _1059 & _4412;
    assign _4417 = _4413 ? _515 : _4416;
    assign _4419 = _1047 ? _1055 : _4417;
    assign _375 = _4419;
    always @(posedge _1038) begin
        if (_1036)
            _4416 <= _1055;
        else
            _4416 <= _375;
    end
    assign _4420 = 9'b010001010;
    assign _4421 = _1062 == _4420;
    assign _4422 = _1059 & _4421;
    assign _4426 = _4422 ? _515 : _4425;
    assign _4428 = _1047 ? _1055 : _4426;
    assign _376 = _4428;
    always @(posedge _1038) begin
        if (_1036)
            _4425 <= _1055;
        else
            _4425 <= _376;
    end
    assign _4429 = 9'b010001001;
    assign _4430 = _1062 == _4429;
    assign _4431 = _1059 & _4430;
    assign _4435 = _4431 ? _515 : _4434;
    assign _4437 = _1047 ? _1055 : _4435;
    assign _377 = _4437;
    always @(posedge _1038) begin
        if (_1036)
            _4434 <= _1055;
        else
            _4434 <= _377;
    end
    assign _4438 = 9'b010001000;
    assign _4439 = _1062 == _4438;
    assign _4440 = _1059 & _4439;
    assign _4444 = _4440 ? _515 : _4443;
    assign _4446 = _1047 ? _1055 : _4444;
    assign _378 = _4446;
    always @(posedge _1038) begin
        if (_1036)
            _4443 <= _1055;
        else
            _4443 <= _378;
    end
    assign _4447 = 9'b010000111;
    assign _4448 = _1062 == _4447;
    assign _4449 = _1059 & _4448;
    assign _4453 = _4449 ? _515 : _4452;
    assign _4455 = _1047 ? _1055 : _4453;
    assign _379 = _4455;
    always @(posedge _1038) begin
        if (_1036)
            _4452 <= _1055;
        else
            _4452 <= _379;
    end
    assign _4456 = 9'b010000110;
    assign _4457 = _1062 == _4456;
    assign _4458 = _1059 & _4457;
    assign _4462 = _4458 ? _515 : _4461;
    assign _4464 = _1047 ? _1055 : _4462;
    assign _380 = _4464;
    always @(posedge _1038) begin
        if (_1036)
            _4461 <= _1055;
        else
            _4461 <= _380;
    end
    assign _4465 = 9'b010000101;
    assign _4466 = _1062 == _4465;
    assign _4467 = _1059 & _4466;
    assign _4471 = _4467 ? _515 : _4470;
    assign _4473 = _1047 ? _1055 : _4471;
    assign _381 = _4473;
    always @(posedge _1038) begin
        if (_1036)
            _4470 <= _1055;
        else
            _4470 <= _381;
    end
    assign _4474 = 9'b010000100;
    assign _4475 = _1062 == _4474;
    assign _4476 = _1059 & _4475;
    assign _4480 = _4476 ? _515 : _4479;
    assign _4482 = _1047 ? _1055 : _4480;
    assign _382 = _4482;
    always @(posedge _1038) begin
        if (_1036)
            _4479 <= _1055;
        else
            _4479 <= _382;
    end
    assign _4483 = 9'b010000011;
    assign _4484 = _1062 == _4483;
    assign _4485 = _1059 & _4484;
    assign _4489 = _4485 ? _515 : _4488;
    assign _4491 = _1047 ? _1055 : _4489;
    assign _383 = _4491;
    always @(posedge _1038) begin
        if (_1036)
            _4488 <= _1055;
        else
            _4488 <= _383;
    end
    assign _4492 = 9'b010000010;
    assign _4493 = _1062 == _4492;
    assign _4494 = _1059 & _4493;
    assign _4498 = _4494 ? _515 : _4497;
    assign _4500 = _1047 ? _1055 : _4498;
    assign _384 = _4500;
    always @(posedge _1038) begin
        if (_1036)
            _4497 <= _1055;
        else
            _4497 <= _384;
    end
    assign _4501 = 9'b010000001;
    assign _4502 = _1062 == _4501;
    assign _4503 = _1059 & _4502;
    assign _4507 = _4503 ? _515 : _4506;
    assign _4509 = _1047 ? _1055 : _4507;
    assign _385 = _4509;
    always @(posedge _1038) begin
        if (_1036)
            _4506 <= _1055;
        else
            _4506 <= _385;
    end
    assign _4510 = 9'b010000000;
    assign _4511 = _1062 == _4510;
    assign _4512 = _1059 & _4511;
    assign _4516 = _4512 ? _515 : _4515;
    assign _4518 = _1047 ? _1055 : _4516;
    assign _386 = _4518;
    always @(posedge _1038) begin
        if (_1036)
            _4515 <= _1055;
        else
            _4515 <= _386;
    end
    assign _4519 = 9'b001111111;
    assign _4520 = _1062 == _4519;
    assign _4521 = _1059 & _4520;
    assign _4525 = _4521 ? _515 : _4524;
    assign _4527 = _1047 ? _1055 : _4525;
    assign _387 = _4527;
    always @(posedge _1038) begin
        if (_1036)
            _4524 <= _1055;
        else
            _4524 <= _387;
    end
    assign _4528 = 9'b001111110;
    assign _4529 = _1062 == _4528;
    assign _4530 = _1059 & _4529;
    assign _4534 = _4530 ? _515 : _4533;
    assign _4536 = _1047 ? _1055 : _4534;
    assign _388 = _4536;
    always @(posedge _1038) begin
        if (_1036)
            _4533 <= _1055;
        else
            _4533 <= _388;
    end
    assign _4537 = 9'b001111101;
    assign _4538 = _1062 == _4537;
    assign _4539 = _1059 & _4538;
    assign _4543 = _4539 ? _515 : _4542;
    assign _4545 = _1047 ? _1055 : _4543;
    assign _389 = _4545;
    always @(posedge _1038) begin
        if (_1036)
            _4542 <= _1055;
        else
            _4542 <= _389;
    end
    assign _4546 = 9'b001111100;
    assign _4547 = _1062 == _4546;
    assign _4548 = _1059 & _4547;
    assign _4552 = _4548 ? _515 : _4551;
    assign _4554 = _1047 ? _1055 : _4552;
    assign _390 = _4554;
    always @(posedge _1038) begin
        if (_1036)
            _4551 <= _1055;
        else
            _4551 <= _390;
    end
    assign _4555 = 9'b001111011;
    assign _4556 = _1062 == _4555;
    assign _4557 = _1059 & _4556;
    assign _4561 = _4557 ? _515 : _4560;
    assign _4563 = _1047 ? _1055 : _4561;
    assign _391 = _4563;
    always @(posedge _1038) begin
        if (_1036)
            _4560 <= _1055;
        else
            _4560 <= _391;
    end
    assign _4564 = 9'b001111010;
    assign _4565 = _1062 == _4564;
    assign _4566 = _1059 & _4565;
    assign _4570 = _4566 ? _515 : _4569;
    assign _4572 = _1047 ? _1055 : _4570;
    assign _392 = _4572;
    always @(posedge _1038) begin
        if (_1036)
            _4569 <= _1055;
        else
            _4569 <= _392;
    end
    assign _4573 = 9'b001111001;
    assign _4574 = _1062 == _4573;
    assign _4575 = _1059 & _4574;
    assign _4579 = _4575 ? _515 : _4578;
    assign _4581 = _1047 ? _1055 : _4579;
    assign _393 = _4581;
    always @(posedge _1038) begin
        if (_1036)
            _4578 <= _1055;
        else
            _4578 <= _393;
    end
    assign _4582 = 9'b001111000;
    assign _4583 = _1062 == _4582;
    assign _4584 = _1059 & _4583;
    assign _4588 = _4584 ? _515 : _4587;
    assign _4590 = _1047 ? _1055 : _4588;
    assign _394 = _4590;
    always @(posedge _1038) begin
        if (_1036)
            _4587 <= _1055;
        else
            _4587 <= _394;
    end
    assign _4591 = 9'b001110111;
    assign _4592 = _1062 == _4591;
    assign _4593 = _1059 & _4592;
    assign _4597 = _4593 ? _515 : _4596;
    assign _4599 = _1047 ? _1055 : _4597;
    assign _395 = _4599;
    always @(posedge _1038) begin
        if (_1036)
            _4596 <= _1055;
        else
            _4596 <= _395;
    end
    assign _4600 = 9'b001110110;
    assign _4601 = _1062 == _4600;
    assign _4602 = _1059 & _4601;
    assign _4606 = _4602 ? _515 : _4605;
    assign _4608 = _1047 ? _1055 : _4606;
    assign _396 = _4608;
    always @(posedge _1038) begin
        if (_1036)
            _4605 <= _1055;
        else
            _4605 <= _396;
    end
    assign _4609 = 9'b001110101;
    assign _4610 = _1062 == _4609;
    assign _4611 = _1059 & _4610;
    assign _4615 = _4611 ? _515 : _4614;
    assign _4617 = _1047 ? _1055 : _4615;
    assign _397 = _4617;
    always @(posedge _1038) begin
        if (_1036)
            _4614 <= _1055;
        else
            _4614 <= _397;
    end
    assign _4618 = 9'b001110100;
    assign _4619 = _1062 == _4618;
    assign _4620 = _1059 & _4619;
    assign _4624 = _4620 ? _515 : _4623;
    assign _4626 = _1047 ? _1055 : _4624;
    assign _398 = _4626;
    always @(posedge _1038) begin
        if (_1036)
            _4623 <= _1055;
        else
            _4623 <= _398;
    end
    assign _4627 = 9'b001110011;
    assign _4628 = _1062 == _4627;
    assign _4629 = _1059 & _4628;
    assign _4633 = _4629 ? _515 : _4632;
    assign _4635 = _1047 ? _1055 : _4633;
    assign _399 = _4635;
    always @(posedge _1038) begin
        if (_1036)
            _4632 <= _1055;
        else
            _4632 <= _399;
    end
    assign _4636 = 9'b001110010;
    assign _4637 = _1062 == _4636;
    assign _4638 = _1059 & _4637;
    assign _4642 = _4638 ? _515 : _4641;
    assign _4644 = _1047 ? _1055 : _4642;
    assign _400 = _4644;
    always @(posedge _1038) begin
        if (_1036)
            _4641 <= _1055;
        else
            _4641 <= _400;
    end
    assign _4645 = 9'b001110001;
    assign _4646 = _1062 == _4645;
    assign _4647 = _1059 & _4646;
    assign _4651 = _4647 ? _515 : _4650;
    assign _4653 = _1047 ? _1055 : _4651;
    assign _401 = _4653;
    always @(posedge _1038) begin
        if (_1036)
            _4650 <= _1055;
        else
            _4650 <= _401;
    end
    assign _4654 = 9'b001110000;
    assign _4655 = _1062 == _4654;
    assign _4656 = _1059 & _4655;
    assign _4660 = _4656 ? _515 : _4659;
    assign _4662 = _1047 ? _1055 : _4660;
    assign _402 = _4662;
    always @(posedge _1038) begin
        if (_1036)
            _4659 <= _1055;
        else
            _4659 <= _402;
    end
    assign _4663 = 9'b001101111;
    assign _4664 = _1062 == _4663;
    assign _4665 = _1059 & _4664;
    assign _4669 = _4665 ? _515 : _4668;
    assign _4671 = _1047 ? _1055 : _4669;
    assign _403 = _4671;
    always @(posedge _1038) begin
        if (_1036)
            _4668 <= _1055;
        else
            _4668 <= _403;
    end
    assign _4672 = 9'b001101110;
    assign _4673 = _1062 == _4672;
    assign _4674 = _1059 & _4673;
    assign _4678 = _4674 ? _515 : _4677;
    assign _4680 = _1047 ? _1055 : _4678;
    assign _404 = _4680;
    always @(posedge _1038) begin
        if (_1036)
            _4677 <= _1055;
        else
            _4677 <= _404;
    end
    assign _4681 = 9'b001101101;
    assign _4682 = _1062 == _4681;
    assign _4683 = _1059 & _4682;
    assign _4687 = _4683 ? _515 : _4686;
    assign _4689 = _1047 ? _1055 : _4687;
    assign _405 = _4689;
    always @(posedge _1038) begin
        if (_1036)
            _4686 <= _1055;
        else
            _4686 <= _405;
    end
    assign _4690 = 9'b001101100;
    assign _4691 = _1062 == _4690;
    assign _4692 = _1059 & _4691;
    assign _4696 = _4692 ? _515 : _4695;
    assign _4698 = _1047 ? _1055 : _4696;
    assign _406 = _4698;
    always @(posedge _1038) begin
        if (_1036)
            _4695 <= _1055;
        else
            _4695 <= _406;
    end
    assign _4699 = 9'b001101011;
    assign _4700 = _1062 == _4699;
    assign _4701 = _1059 & _4700;
    assign _4705 = _4701 ? _515 : _4704;
    assign _4707 = _1047 ? _1055 : _4705;
    assign _407 = _4707;
    always @(posedge _1038) begin
        if (_1036)
            _4704 <= _1055;
        else
            _4704 <= _407;
    end
    assign _4708 = 9'b001101010;
    assign _4709 = _1062 == _4708;
    assign _4710 = _1059 & _4709;
    assign _4714 = _4710 ? _515 : _4713;
    assign _4716 = _1047 ? _1055 : _4714;
    assign _408 = _4716;
    always @(posedge _1038) begin
        if (_1036)
            _4713 <= _1055;
        else
            _4713 <= _408;
    end
    assign _4717 = 9'b001101001;
    assign _4718 = _1062 == _4717;
    assign _4719 = _1059 & _4718;
    assign _4723 = _4719 ? _515 : _4722;
    assign _4725 = _1047 ? _1055 : _4723;
    assign _409 = _4725;
    always @(posedge _1038) begin
        if (_1036)
            _4722 <= _1055;
        else
            _4722 <= _409;
    end
    assign _4726 = 9'b001101000;
    assign _4727 = _1062 == _4726;
    assign _4728 = _1059 & _4727;
    assign _4732 = _4728 ? _515 : _4731;
    assign _4734 = _1047 ? _1055 : _4732;
    assign _410 = _4734;
    always @(posedge _1038) begin
        if (_1036)
            _4731 <= _1055;
        else
            _4731 <= _410;
    end
    assign _4735 = 9'b001100111;
    assign _4736 = _1062 == _4735;
    assign _4737 = _1059 & _4736;
    assign _4741 = _4737 ? _515 : _4740;
    assign _4743 = _1047 ? _1055 : _4741;
    assign _411 = _4743;
    always @(posedge _1038) begin
        if (_1036)
            _4740 <= _1055;
        else
            _4740 <= _411;
    end
    assign _4744 = 9'b001100110;
    assign _4745 = _1062 == _4744;
    assign _4746 = _1059 & _4745;
    assign _4750 = _4746 ? _515 : _4749;
    assign _4752 = _1047 ? _1055 : _4750;
    assign _412 = _4752;
    always @(posedge _1038) begin
        if (_1036)
            _4749 <= _1055;
        else
            _4749 <= _412;
    end
    assign _4753 = 9'b001100101;
    assign _4754 = _1062 == _4753;
    assign _4755 = _1059 & _4754;
    assign _4759 = _4755 ? _515 : _4758;
    assign _4761 = _1047 ? _1055 : _4759;
    assign _413 = _4761;
    always @(posedge _1038) begin
        if (_1036)
            _4758 <= _1055;
        else
            _4758 <= _413;
    end
    assign _4762 = 9'b001100100;
    assign _4763 = _1062 == _4762;
    assign _4764 = _1059 & _4763;
    assign _4768 = _4764 ? _515 : _4767;
    assign _4770 = _1047 ? _1055 : _4768;
    assign _414 = _4770;
    always @(posedge _1038) begin
        if (_1036)
            _4767 <= _1055;
        else
            _4767 <= _414;
    end
    assign _4771 = 9'b001100011;
    assign _4772 = _1062 == _4771;
    assign _4773 = _1059 & _4772;
    assign _4777 = _4773 ? _515 : _4776;
    assign _4779 = _1047 ? _1055 : _4777;
    assign _415 = _4779;
    always @(posedge _1038) begin
        if (_1036)
            _4776 <= _1055;
        else
            _4776 <= _415;
    end
    assign _4780 = 9'b001100010;
    assign _4781 = _1062 == _4780;
    assign _4782 = _1059 & _4781;
    assign _4786 = _4782 ? _515 : _4785;
    assign _4788 = _1047 ? _1055 : _4786;
    assign _416 = _4788;
    always @(posedge _1038) begin
        if (_1036)
            _4785 <= _1055;
        else
            _4785 <= _416;
    end
    assign _4789 = 9'b001100001;
    assign _4790 = _1062 == _4789;
    assign _4791 = _1059 & _4790;
    assign _4795 = _4791 ? _515 : _4794;
    assign _4797 = _1047 ? _1055 : _4795;
    assign _417 = _4797;
    always @(posedge _1038) begin
        if (_1036)
            _4794 <= _1055;
        else
            _4794 <= _417;
    end
    assign _4798 = 9'b001100000;
    assign _4799 = _1062 == _4798;
    assign _4800 = _1059 & _4799;
    assign _4804 = _4800 ? _515 : _4803;
    assign _4806 = _1047 ? _1055 : _4804;
    assign _418 = _4806;
    always @(posedge _1038) begin
        if (_1036)
            _4803 <= _1055;
        else
            _4803 <= _418;
    end
    assign _4807 = 9'b001011111;
    assign _4808 = _1062 == _4807;
    assign _4809 = _1059 & _4808;
    assign _4813 = _4809 ? _515 : _4812;
    assign _4815 = _1047 ? _1055 : _4813;
    assign _419 = _4815;
    always @(posedge _1038) begin
        if (_1036)
            _4812 <= _1055;
        else
            _4812 <= _419;
    end
    assign _4816 = 9'b001011110;
    assign _4817 = _1062 == _4816;
    assign _4818 = _1059 & _4817;
    assign _4822 = _4818 ? _515 : _4821;
    assign _4824 = _1047 ? _1055 : _4822;
    assign _420 = _4824;
    always @(posedge _1038) begin
        if (_1036)
            _4821 <= _1055;
        else
            _4821 <= _420;
    end
    assign _4825 = 9'b001011101;
    assign _4826 = _1062 == _4825;
    assign _4827 = _1059 & _4826;
    assign _4831 = _4827 ? _515 : _4830;
    assign _4833 = _1047 ? _1055 : _4831;
    assign _421 = _4833;
    always @(posedge _1038) begin
        if (_1036)
            _4830 <= _1055;
        else
            _4830 <= _421;
    end
    assign _4834 = 9'b001011100;
    assign _4835 = _1062 == _4834;
    assign _4836 = _1059 & _4835;
    assign _4840 = _4836 ? _515 : _4839;
    assign _4842 = _1047 ? _1055 : _4840;
    assign _422 = _4842;
    always @(posedge _1038) begin
        if (_1036)
            _4839 <= _1055;
        else
            _4839 <= _422;
    end
    assign _4843 = 9'b001011011;
    assign _4844 = _1062 == _4843;
    assign _4845 = _1059 & _4844;
    assign _4849 = _4845 ? _515 : _4848;
    assign _4851 = _1047 ? _1055 : _4849;
    assign _423 = _4851;
    always @(posedge _1038) begin
        if (_1036)
            _4848 <= _1055;
        else
            _4848 <= _423;
    end
    assign _4852 = 9'b001011010;
    assign _4853 = _1062 == _4852;
    assign _4854 = _1059 & _4853;
    assign _4858 = _4854 ? _515 : _4857;
    assign _4860 = _1047 ? _1055 : _4858;
    assign _424 = _4860;
    always @(posedge _1038) begin
        if (_1036)
            _4857 <= _1055;
        else
            _4857 <= _424;
    end
    assign _4861 = 9'b001011001;
    assign _4862 = _1062 == _4861;
    assign _4863 = _1059 & _4862;
    assign _4867 = _4863 ? _515 : _4866;
    assign _4869 = _1047 ? _1055 : _4867;
    assign _425 = _4869;
    always @(posedge _1038) begin
        if (_1036)
            _4866 <= _1055;
        else
            _4866 <= _425;
    end
    assign _4870 = 9'b001011000;
    assign _4871 = _1062 == _4870;
    assign _4872 = _1059 & _4871;
    assign _4876 = _4872 ? _515 : _4875;
    assign _4878 = _1047 ? _1055 : _4876;
    assign _426 = _4878;
    always @(posedge _1038) begin
        if (_1036)
            _4875 <= _1055;
        else
            _4875 <= _426;
    end
    assign _4879 = 9'b001010111;
    assign _4880 = _1062 == _4879;
    assign _4881 = _1059 & _4880;
    assign _4885 = _4881 ? _515 : _4884;
    assign _4887 = _1047 ? _1055 : _4885;
    assign _427 = _4887;
    always @(posedge _1038) begin
        if (_1036)
            _4884 <= _1055;
        else
            _4884 <= _427;
    end
    assign _4888 = 9'b001010110;
    assign _4889 = _1062 == _4888;
    assign _4890 = _1059 & _4889;
    assign _4894 = _4890 ? _515 : _4893;
    assign _4896 = _1047 ? _1055 : _4894;
    assign _428 = _4896;
    always @(posedge _1038) begin
        if (_1036)
            _4893 <= _1055;
        else
            _4893 <= _428;
    end
    assign _4897 = 9'b001010101;
    assign _4898 = _1062 == _4897;
    assign _4899 = _1059 & _4898;
    assign _4903 = _4899 ? _515 : _4902;
    assign _4905 = _1047 ? _1055 : _4903;
    assign _429 = _4905;
    always @(posedge _1038) begin
        if (_1036)
            _4902 <= _1055;
        else
            _4902 <= _429;
    end
    assign _4906 = 9'b001010100;
    assign _4907 = _1062 == _4906;
    assign _4908 = _1059 & _4907;
    assign _4912 = _4908 ? _515 : _4911;
    assign _4914 = _1047 ? _1055 : _4912;
    assign _430 = _4914;
    always @(posedge _1038) begin
        if (_1036)
            _4911 <= _1055;
        else
            _4911 <= _430;
    end
    assign _4915 = 9'b001010011;
    assign _4916 = _1062 == _4915;
    assign _4917 = _1059 & _4916;
    assign _4921 = _4917 ? _515 : _4920;
    assign _4923 = _1047 ? _1055 : _4921;
    assign _431 = _4923;
    always @(posedge _1038) begin
        if (_1036)
            _4920 <= _1055;
        else
            _4920 <= _431;
    end
    assign _4924 = 9'b001010010;
    assign _4925 = _1062 == _4924;
    assign _4926 = _1059 & _4925;
    assign _4930 = _4926 ? _515 : _4929;
    assign _4932 = _1047 ? _1055 : _4930;
    assign _432 = _4932;
    always @(posedge _1038) begin
        if (_1036)
            _4929 <= _1055;
        else
            _4929 <= _432;
    end
    assign _4933 = 9'b001010001;
    assign _4934 = _1062 == _4933;
    assign _4935 = _1059 & _4934;
    assign _4939 = _4935 ? _515 : _4938;
    assign _4941 = _1047 ? _1055 : _4939;
    assign _433 = _4941;
    always @(posedge _1038) begin
        if (_1036)
            _4938 <= _1055;
        else
            _4938 <= _433;
    end
    assign _4942 = 9'b001010000;
    assign _4943 = _1062 == _4942;
    assign _4944 = _1059 & _4943;
    assign _4948 = _4944 ? _515 : _4947;
    assign _4950 = _1047 ? _1055 : _4948;
    assign _434 = _4950;
    always @(posedge _1038) begin
        if (_1036)
            _4947 <= _1055;
        else
            _4947 <= _434;
    end
    assign _4951 = 9'b001001111;
    assign _4952 = _1062 == _4951;
    assign _4953 = _1059 & _4952;
    assign _4957 = _4953 ? _515 : _4956;
    assign _4959 = _1047 ? _1055 : _4957;
    assign _435 = _4959;
    always @(posedge _1038) begin
        if (_1036)
            _4956 <= _1055;
        else
            _4956 <= _435;
    end
    assign _4960 = 9'b001001110;
    assign _4961 = _1062 == _4960;
    assign _4962 = _1059 & _4961;
    assign _4966 = _4962 ? _515 : _4965;
    assign _4968 = _1047 ? _1055 : _4966;
    assign _436 = _4968;
    always @(posedge _1038) begin
        if (_1036)
            _4965 <= _1055;
        else
            _4965 <= _436;
    end
    assign _4969 = 9'b001001101;
    assign _4970 = _1062 == _4969;
    assign _4971 = _1059 & _4970;
    assign _4975 = _4971 ? _515 : _4974;
    assign _4977 = _1047 ? _1055 : _4975;
    assign _437 = _4977;
    always @(posedge _1038) begin
        if (_1036)
            _4974 <= _1055;
        else
            _4974 <= _437;
    end
    assign _4978 = 9'b001001100;
    assign _4979 = _1062 == _4978;
    assign _4980 = _1059 & _4979;
    assign _4984 = _4980 ? _515 : _4983;
    assign _4986 = _1047 ? _1055 : _4984;
    assign _438 = _4986;
    always @(posedge _1038) begin
        if (_1036)
            _4983 <= _1055;
        else
            _4983 <= _438;
    end
    assign _4987 = 9'b001001011;
    assign _4988 = _1062 == _4987;
    assign _4989 = _1059 & _4988;
    assign _4993 = _4989 ? _515 : _4992;
    assign _4995 = _1047 ? _1055 : _4993;
    assign _439 = _4995;
    always @(posedge _1038) begin
        if (_1036)
            _4992 <= _1055;
        else
            _4992 <= _439;
    end
    assign _4996 = 9'b001001010;
    assign _4997 = _1062 == _4996;
    assign _4998 = _1059 & _4997;
    assign _5002 = _4998 ? _515 : _5001;
    assign _5004 = _1047 ? _1055 : _5002;
    assign _440 = _5004;
    always @(posedge _1038) begin
        if (_1036)
            _5001 <= _1055;
        else
            _5001 <= _440;
    end
    assign _5005 = 9'b001001001;
    assign _5006 = _1062 == _5005;
    assign _5007 = _1059 & _5006;
    assign _5011 = _5007 ? _515 : _5010;
    assign _5013 = _1047 ? _1055 : _5011;
    assign _441 = _5013;
    always @(posedge _1038) begin
        if (_1036)
            _5010 <= _1055;
        else
            _5010 <= _441;
    end
    assign _5014 = 9'b001001000;
    assign _5015 = _1062 == _5014;
    assign _5016 = _1059 & _5015;
    assign _5020 = _5016 ? _515 : _5019;
    assign _5022 = _1047 ? _1055 : _5020;
    assign _442 = _5022;
    always @(posedge _1038) begin
        if (_1036)
            _5019 <= _1055;
        else
            _5019 <= _442;
    end
    assign _5023 = 9'b001000111;
    assign _5024 = _1062 == _5023;
    assign _5025 = _1059 & _5024;
    assign _5029 = _5025 ? _515 : _5028;
    assign _5031 = _1047 ? _1055 : _5029;
    assign _443 = _5031;
    always @(posedge _1038) begin
        if (_1036)
            _5028 <= _1055;
        else
            _5028 <= _443;
    end
    assign _5032 = 9'b001000110;
    assign _5033 = _1062 == _5032;
    assign _5034 = _1059 & _5033;
    assign _5038 = _5034 ? _515 : _5037;
    assign _5040 = _1047 ? _1055 : _5038;
    assign _444 = _5040;
    always @(posedge _1038) begin
        if (_1036)
            _5037 <= _1055;
        else
            _5037 <= _444;
    end
    assign _5041 = 9'b001000101;
    assign _5042 = _1062 == _5041;
    assign _5043 = _1059 & _5042;
    assign _5047 = _5043 ? _515 : _5046;
    assign _5049 = _1047 ? _1055 : _5047;
    assign _445 = _5049;
    always @(posedge _1038) begin
        if (_1036)
            _5046 <= _1055;
        else
            _5046 <= _445;
    end
    assign _5050 = 9'b001000100;
    assign _5051 = _1062 == _5050;
    assign _5052 = _1059 & _5051;
    assign _5056 = _5052 ? _515 : _5055;
    assign _5058 = _1047 ? _1055 : _5056;
    assign _446 = _5058;
    always @(posedge _1038) begin
        if (_1036)
            _5055 <= _1055;
        else
            _5055 <= _446;
    end
    assign _5059 = 9'b001000011;
    assign _5060 = _1062 == _5059;
    assign _5061 = _1059 & _5060;
    assign _5065 = _5061 ? _515 : _5064;
    assign _5067 = _1047 ? _1055 : _5065;
    assign _447 = _5067;
    always @(posedge _1038) begin
        if (_1036)
            _5064 <= _1055;
        else
            _5064 <= _447;
    end
    assign _5068 = 9'b001000010;
    assign _5069 = _1062 == _5068;
    assign _5070 = _1059 & _5069;
    assign _5074 = _5070 ? _515 : _5073;
    assign _5076 = _1047 ? _1055 : _5074;
    assign _448 = _5076;
    always @(posedge _1038) begin
        if (_1036)
            _5073 <= _1055;
        else
            _5073 <= _448;
    end
    assign _5077 = 9'b001000001;
    assign _5078 = _1062 == _5077;
    assign _5079 = _1059 & _5078;
    assign _5083 = _5079 ? _515 : _5082;
    assign _5085 = _1047 ? _1055 : _5083;
    assign _449 = _5085;
    always @(posedge _1038) begin
        if (_1036)
            _5082 <= _1055;
        else
            _5082 <= _449;
    end
    assign _5086 = 9'b001000000;
    assign _5087 = _1062 == _5086;
    assign _5088 = _1059 & _5087;
    assign _5092 = _5088 ? _515 : _5091;
    assign _5094 = _1047 ? _1055 : _5092;
    assign _450 = _5094;
    always @(posedge _1038) begin
        if (_1036)
            _5091 <= _1055;
        else
            _5091 <= _450;
    end
    assign _5095 = 9'b000111111;
    assign _5096 = _1062 == _5095;
    assign _5097 = _1059 & _5096;
    assign _5101 = _5097 ? _515 : _5100;
    assign _5103 = _1047 ? _1055 : _5101;
    assign _451 = _5103;
    always @(posedge _1038) begin
        if (_1036)
            _5100 <= _1055;
        else
            _5100 <= _451;
    end
    assign _5104 = 9'b000111110;
    assign _5105 = _1062 == _5104;
    assign _5106 = _1059 & _5105;
    assign _5110 = _5106 ? _515 : _5109;
    assign _5112 = _1047 ? _1055 : _5110;
    assign _452 = _5112;
    always @(posedge _1038) begin
        if (_1036)
            _5109 <= _1055;
        else
            _5109 <= _452;
    end
    assign _5113 = 9'b000111101;
    assign _5114 = _1062 == _5113;
    assign _5115 = _1059 & _5114;
    assign _5119 = _5115 ? _515 : _5118;
    assign _5121 = _1047 ? _1055 : _5119;
    assign _453 = _5121;
    always @(posedge _1038) begin
        if (_1036)
            _5118 <= _1055;
        else
            _5118 <= _453;
    end
    assign _5122 = 9'b000111100;
    assign _5123 = _1062 == _5122;
    assign _5124 = _1059 & _5123;
    assign _5128 = _5124 ? _515 : _5127;
    assign _5130 = _1047 ? _1055 : _5128;
    assign _454 = _5130;
    always @(posedge _1038) begin
        if (_1036)
            _5127 <= _1055;
        else
            _5127 <= _454;
    end
    assign _5131 = 9'b000111011;
    assign _5132 = _1062 == _5131;
    assign _5133 = _1059 & _5132;
    assign _5137 = _5133 ? _515 : _5136;
    assign _5139 = _1047 ? _1055 : _5137;
    assign _455 = _5139;
    always @(posedge _1038) begin
        if (_1036)
            _5136 <= _1055;
        else
            _5136 <= _455;
    end
    assign _5140 = 9'b000111010;
    assign _5141 = _1062 == _5140;
    assign _5142 = _1059 & _5141;
    assign _5146 = _5142 ? _515 : _5145;
    assign _5148 = _1047 ? _1055 : _5146;
    assign _456 = _5148;
    always @(posedge _1038) begin
        if (_1036)
            _5145 <= _1055;
        else
            _5145 <= _456;
    end
    assign _5149 = 9'b000111001;
    assign _5150 = _1062 == _5149;
    assign _5151 = _1059 & _5150;
    assign _5155 = _5151 ? _515 : _5154;
    assign _5157 = _1047 ? _1055 : _5155;
    assign _457 = _5157;
    always @(posedge _1038) begin
        if (_1036)
            _5154 <= _1055;
        else
            _5154 <= _457;
    end
    assign _5158 = 9'b000111000;
    assign _5159 = _1062 == _5158;
    assign _5160 = _1059 & _5159;
    assign _5164 = _5160 ? _515 : _5163;
    assign _5166 = _1047 ? _1055 : _5164;
    assign _458 = _5166;
    always @(posedge _1038) begin
        if (_1036)
            _5163 <= _1055;
        else
            _5163 <= _458;
    end
    assign _5167 = 9'b000110111;
    assign _5168 = _1062 == _5167;
    assign _5169 = _1059 & _5168;
    assign _5173 = _5169 ? _515 : _5172;
    assign _5175 = _1047 ? _1055 : _5173;
    assign _459 = _5175;
    always @(posedge _1038) begin
        if (_1036)
            _5172 <= _1055;
        else
            _5172 <= _459;
    end
    assign _5176 = 9'b000110110;
    assign _5177 = _1062 == _5176;
    assign _5178 = _1059 & _5177;
    assign _5182 = _5178 ? _515 : _5181;
    assign _5184 = _1047 ? _1055 : _5182;
    assign _460 = _5184;
    always @(posedge _1038) begin
        if (_1036)
            _5181 <= _1055;
        else
            _5181 <= _460;
    end
    assign _5185 = 9'b000110101;
    assign _5186 = _1062 == _5185;
    assign _5187 = _1059 & _5186;
    assign _5191 = _5187 ? _515 : _5190;
    assign _5193 = _1047 ? _1055 : _5191;
    assign _461 = _5193;
    always @(posedge _1038) begin
        if (_1036)
            _5190 <= _1055;
        else
            _5190 <= _461;
    end
    assign _5194 = 9'b000110100;
    assign _5195 = _1062 == _5194;
    assign _5196 = _1059 & _5195;
    assign _5200 = _5196 ? _515 : _5199;
    assign _5202 = _1047 ? _1055 : _5200;
    assign _462 = _5202;
    always @(posedge _1038) begin
        if (_1036)
            _5199 <= _1055;
        else
            _5199 <= _462;
    end
    assign _5203 = 9'b000110011;
    assign _5204 = _1062 == _5203;
    assign _5205 = _1059 & _5204;
    assign _5209 = _5205 ? _515 : _5208;
    assign _5211 = _1047 ? _1055 : _5209;
    assign _463 = _5211;
    always @(posedge _1038) begin
        if (_1036)
            _5208 <= _1055;
        else
            _5208 <= _463;
    end
    assign _5212 = 9'b000110010;
    assign _5213 = _1062 == _5212;
    assign _5214 = _1059 & _5213;
    assign _5218 = _5214 ? _515 : _5217;
    assign _5220 = _1047 ? _1055 : _5218;
    assign _464 = _5220;
    always @(posedge _1038) begin
        if (_1036)
            _5217 <= _1055;
        else
            _5217 <= _464;
    end
    assign _5221 = 9'b000110001;
    assign _5222 = _1062 == _5221;
    assign _5223 = _1059 & _5222;
    assign _5227 = _5223 ? _515 : _5226;
    assign _5229 = _1047 ? _1055 : _5227;
    assign _465 = _5229;
    always @(posedge _1038) begin
        if (_1036)
            _5226 <= _1055;
        else
            _5226 <= _465;
    end
    assign _5230 = 9'b000110000;
    assign _5231 = _1062 == _5230;
    assign _5232 = _1059 & _5231;
    assign _5236 = _5232 ? _515 : _5235;
    assign _5238 = _1047 ? _1055 : _5236;
    assign _466 = _5238;
    always @(posedge _1038) begin
        if (_1036)
            _5235 <= _1055;
        else
            _5235 <= _466;
    end
    assign _5239 = 9'b000101111;
    assign _5240 = _1062 == _5239;
    assign _5241 = _1059 & _5240;
    assign _5245 = _5241 ? _515 : _5244;
    assign _5247 = _1047 ? _1055 : _5245;
    assign _467 = _5247;
    always @(posedge _1038) begin
        if (_1036)
            _5244 <= _1055;
        else
            _5244 <= _467;
    end
    assign _5248 = 9'b000101110;
    assign _5249 = _1062 == _5248;
    assign _5250 = _1059 & _5249;
    assign _5254 = _5250 ? _515 : _5253;
    assign _5256 = _1047 ? _1055 : _5254;
    assign _468 = _5256;
    always @(posedge _1038) begin
        if (_1036)
            _5253 <= _1055;
        else
            _5253 <= _468;
    end
    assign _5257 = 9'b000101101;
    assign _5258 = _1062 == _5257;
    assign _5259 = _1059 & _5258;
    assign _5263 = _5259 ? _515 : _5262;
    assign _5265 = _1047 ? _1055 : _5263;
    assign _469 = _5265;
    always @(posedge _1038) begin
        if (_1036)
            _5262 <= _1055;
        else
            _5262 <= _469;
    end
    assign _5266 = 9'b000101100;
    assign _5267 = _1062 == _5266;
    assign _5268 = _1059 & _5267;
    assign _5272 = _5268 ? _515 : _5271;
    assign _5274 = _1047 ? _1055 : _5272;
    assign _470 = _5274;
    always @(posedge _1038) begin
        if (_1036)
            _5271 <= _1055;
        else
            _5271 <= _470;
    end
    assign _5275 = 9'b000101011;
    assign _5276 = _1062 == _5275;
    assign _5277 = _1059 & _5276;
    assign _5281 = _5277 ? _515 : _5280;
    assign _5283 = _1047 ? _1055 : _5281;
    assign _471 = _5283;
    always @(posedge _1038) begin
        if (_1036)
            _5280 <= _1055;
        else
            _5280 <= _471;
    end
    assign _5284 = 9'b000101010;
    assign _5285 = _1062 == _5284;
    assign _5286 = _1059 & _5285;
    assign _5290 = _5286 ? _515 : _5289;
    assign _5292 = _1047 ? _1055 : _5290;
    assign _472 = _5292;
    always @(posedge _1038) begin
        if (_1036)
            _5289 <= _1055;
        else
            _5289 <= _472;
    end
    assign _5293 = 9'b000101001;
    assign _5294 = _1062 == _5293;
    assign _5295 = _1059 & _5294;
    assign _5299 = _5295 ? _515 : _5298;
    assign _5301 = _1047 ? _1055 : _5299;
    assign _473 = _5301;
    always @(posedge _1038) begin
        if (_1036)
            _5298 <= _1055;
        else
            _5298 <= _473;
    end
    assign _5302 = 9'b000101000;
    assign _5303 = _1062 == _5302;
    assign _5304 = _1059 & _5303;
    assign _5308 = _5304 ? _515 : _5307;
    assign _5310 = _1047 ? _1055 : _5308;
    assign _474 = _5310;
    always @(posedge _1038) begin
        if (_1036)
            _5307 <= _1055;
        else
            _5307 <= _474;
    end
    assign _5311 = 9'b000100111;
    assign _5312 = _1062 == _5311;
    assign _5313 = _1059 & _5312;
    assign _5317 = _5313 ? _515 : _5316;
    assign _5319 = _1047 ? _1055 : _5317;
    assign _475 = _5319;
    always @(posedge _1038) begin
        if (_1036)
            _5316 <= _1055;
        else
            _5316 <= _475;
    end
    assign _5320 = 9'b000100110;
    assign _5321 = _1062 == _5320;
    assign _5322 = _1059 & _5321;
    assign _5326 = _5322 ? _515 : _5325;
    assign _5328 = _1047 ? _1055 : _5326;
    assign _476 = _5328;
    always @(posedge _1038) begin
        if (_1036)
            _5325 <= _1055;
        else
            _5325 <= _476;
    end
    assign _5329 = 9'b000100101;
    assign _5330 = _1062 == _5329;
    assign _5331 = _1059 & _5330;
    assign _5335 = _5331 ? _515 : _5334;
    assign _5337 = _1047 ? _1055 : _5335;
    assign _477 = _5337;
    always @(posedge _1038) begin
        if (_1036)
            _5334 <= _1055;
        else
            _5334 <= _477;
    end
    assign _5338 = 9'b000100100;
    assign _5339 = _1062 == _5338;
    assign _5340 = _1059 & _5339;
    assign _5344 = _5340 ? _515 : _5343;
    assign _5346 = _1047 ? _1055 : _5344;
    assign _478 = _5346;
    always @(posedge _1038) begin
        if (_1036)
            _5343 <= _1055;
        else
            _5343 <= _478;
    end
    assign _5347 = 9'b000100011;
    assign _5348 = _1062 == _5347;
    assign _5349 = _1059 & _5348;
    assign _5353 = _5349 ? _515 : _5352;
    assign _5355 = _1047 ? _1055 : _5353;
    assign _479 = _5355;
    always @(posedge _1038) begin
        if (_1036)
            _5352 <= _1055;
        else
            _5352 <= _479;
    end
    assign _5356 = 9'b000100010;
    assign _5357 = _1062 == _5356;
    assign _5358 = _1059 & _5357;
    assign _5362 = _5358 ? _515 : _5361;
    assign _5364 = _1047 ? _1055 : _5362;
    assign _480 = _5364;
    always @(posedge _1038) begin
        if (_1036)
            _5361 <= _1055;
        else
            _5361 <= _480;
    end
    assign _5365 = 9'b000100001;
    assign _5366 = _1062 == _5365;
    assign _5367 = _1059 & _5366;
    assign _5371 = _5367 ? _515 : _5370;
    assign _5373 = _1047 ? _1055 : _5371;
    assign _481 = _5373;
    always @(posedge _1038) begin
        if (_1036)
            _5370 <= _1055;
        else
            _5370 <= _481;
    end
    assign _5374 = 9'b000100000;
    assign _5375 = _1062 == _5374;
    assign _5376 = _1059 & _5375;
    assign _5380 = _5376 ? _515 : _5379;
    assign _5382 = _1047 ? _1055 : _5380;
    assign _482 = _5382;
    always @(posedge _1038) begin
        if (_1036)
            _5379 <= _1055;
        else
            _5379 <= _482;
    end
    assign _5383 = 9'b000011111;
    assign _5384 = _1062 == _5383;
    assign _5385 = _1059 & _5384;
    assign _5389 = _5385 ? _515 : _5388;
    assign _5391 = _1047 ? _1055 : _5389;
    assign _483 = _5391;
    always @(posedge _1038) begin
        if (_1036)
            _5388 <= _1055;
        else
            _5388 <= _483;
    end
    assign _5392 = 9'b000011110;
    assign _5393 = _1062 == _5392;
    assign _5394 = _1059 & _5393;
    assign _5398 = _5394 ? _515 : _5397;
    assign _5400 = _1047 ? _1055 : _5398;
    assign _484 = _5400;
    always @(posedge _1038) begin
        if (_1036)
            _5397 <= _1055;
        else
            _5397 <= _484;
    end
    assign _5401 = 9'b000011101;
    assign _5402 = _1062 == _5401;
    assign _5403 = _1059 & _5402;
    assign _5407 = _5403 ? _515 : _5406;
    assign _5409 = _1047 ? _1055 : _5407;
    assign _485 = _5409;
    always @(posedge _1038) begin
        if (_1036)
            _5406 <= _1055;
        else
            _5406 <= _485;
    end
    assign _5410 = 9'b000011100;
    assign _5411 = _1062 == _5410;
    assign _5412 = _1059 & _5411;
    assign _5416 = _5412 ? _515 : _5415;
    assign _5418 = _1047 ? _1055 : _5416;
    assign _486 = _5418;
    always @(posedge _1038) begin
        if (_1036)
            _5415 <= _1055;
        else
            _5415 <= _486;
    end
    assign _5419 = 9'b000011011;
    assign _5420 = _1062 == _5419;
    assign _5421 = _1059 & _5420;
    assign _5425 = _5421 ? _515 : _5424;
    assign _5427 = _1047 ? _1055 : _5425;
    assign _487 = _5427;
    always @(posedge _1038) begin
        if (_1036)
            _5424 <= _1055;
        else
            _5424 <= _487;
    end
    assign _5428 = 9'b000011010;
    assign _5429 = _1062 == _5428;
    assign _5430 = _1059 & _5429;
    assign _5434 = _5430 ? _515 : _5433;
    assign _5436 = _1047 ? _1055 : _5434;
    assign _488 = _5436;
    always @(posedge _1038) begin
        if (_1036)
            _5433 <= _1055;
        else
            _5433 <= _488;
    end
    assign _5437 = 9'b000011001;
    assign _5438 = _1062 == _5437;
    assign _5439 = _1059 & _5438;
    assign _5443 = _5439 ? _515 : _5442;
    assign _5445 = _1047 ? _1055 : _5443;
    assign _489 = _5445;
    always @(posedge _1038) begin
        if (_1036)
            _5442 <= _1055;
        else
            _5442 <= _489;
    end
    assign _5446 = 9'b000011000;
    assign _5447 = _1062 == _5446;
    assign _5448 = _1059 & _5447;
    assign _5452 = _5448 ? _515 : _5451;
    assign _5454 = _1047 ? _1055 : _5452;
    assign _490 = _5454;
    always @(posedge _1038) begin
        if (_1036)
            _5451 <= _1055;
        else
            _5451 <= _490;
    end
    assign _5455 = 9'b000010111;
    assign _5456 = _1062 == _5455;
    assign _5457 = _1059 & _5456;
    assign _5461 = _5457 ? _515 : _5460;
    assign _5463 = _1047 ? _1055 : _5461;
    assign _491 = _5463;
    always @(posedge _1038) begin
        if (_1036)
            _5460 <= _1055;
        else
            _5460 <= _491;
    end
    assign _5464 = 9'b000010110;
    assign _5465 = _1062 == _5464;
    assign _5466 = _1059 & _5465;
    assign _5470 = _5466 ? _515 : _5469;
    assign _5472 = _1047 ? _1055 : _5470;
    assign _492 = _5472;
    always @(posedge _1038) begin
        if (_1036)
            _5469 <= _1055;
        else
            _5469 <= _492;
    end
    assign _5473 = 9'b000010101;
    assign _5474 = _1062 == _5473;
    assign _5475 = _1059 & _5474;
    assign _5479 = _5475 ? _515 : _5478;
    assign _5481 = _1047 ? _1055 : _5479;
    assign _493 = _5481;
    always @(posedge _1038) begin
        if (_1036)
            _5478 <= _1055;
        else
            _5478 <= _493;
    end
    assign _5482 = 9'b000010100;
    assign _5483 = _1062 == _5482;
    assign _5484 = _1059 & _5483;
    assign _5488 = _5484 ? _515 : _5487;
    assign _5490 = _1047 ? _1055 : _5488;
    assign _494 = _5490;
    always @(posedge _1038) begin
        if (_1036)
            _5487 <= _1055;
        else
            _5487 <= _494;
    end
    assign _5491 = 9'b000010011;
    assign _5492 = _1062 == _5491;
    assign _5493 = _1059 & _5492;
    assign _5497 = _5493 ? _515 : _5496;
    assign _5499 = _1047 ? _1055 : _5497;
    assign _495 = _5499;
    always @(posedge _1038) begin
        if (_1036)
            _5496 <= _1055;
        else
            _5496 <= _495;
    end
    assign _5500 = 9'b000010010;
    assign _5501 = _1062 == _5500;
    assign _5502 = _1059 & _5501;
    assign _5506 = _5502 ? _515 : _5505;
    assign _5508 = _1047 ? _1055 : _5506;
    assign _496 = _5508;
    always @(posedge _1038) begin
        if (_1036)
            _5505 <= _1055;
        else
            _5505 <= _496;
    end
    assign _5509 = 9'b000010001;
    assign _5510 = _1062 == _5509;
    assign _5511 = _1059 & _5510;
    assign _5515 = _5511 ? _515 : _5514;
    assign _5517 = _1047 ? _1055 : _5515;
    assign _497 = _5517;
    always @(posedge _1038) begin
        if (_1036)
            _5514 <= _1055;
        else
            _5514 <= _497;
    end
    assign _5518 = 9'b000010000;
    assign _5519 = _1062 == _5518;
    assign _5520 = _1059 & _5519;
    assign _5524 = _5520 ? _515 : _5523;
    assign _5526 = _1047 ? _1055 : _5524;
    assign _498 = _5526;
    always @(posedge _1038) begin
        if (_1036)
            _5523 <= _1055;
        else
            _5523 <= _498;
    end
    assign _5527 = 9'b000001111;
    assign _5528 = _1062 == _5527;
    assign _5529 = _1059 & _5528;
    assign _5533 = _5529 ? _515 : _5532;
    assign _5535 = _1047 ? _1055 : _5533;
    assign _499 = _5535;
    always @(posedge _1038) begin
        if (_1036)
            _5532 <= _1055;
        else
            _5532 <= _499;
    end
    assign _5536 = 9'b000001110;
    assign _5537 = _1062 == _5536;
    assign _5538 = _1059 & _5537;
    assign _5542 = _5538 ? _515 : _5541;
    assign _5544 = _1047 ? _1055 : _5542;
    assign _500 = _5544;
    always @(posedge _1038) begin
        if (_1036)
            _5541 <= _1055;
        else
            _5541 <= _500;
    end
    assign _5545 = 9'b000001101;
    assign _5546 = _1062 == _5545;
    assign _5547 = _1059 & _5546;
    assign _5551 = _5547 ? _515 : _5550;
    assign _5553 = _1047 ? _1055 : _5551;
    assign _501 = _5553;
    always @(posedge _1038) begin
        if (_1036)
            _5550 <= _1055;
        else
            _5550 <= _501;
    end
    assign _5554 = 9'b000001100;
    assign _5555 = _1062 == _5554;
    assign _5556 = _1059 & _5555;
    assign _5560 = _5556 ? _515 : _5559;
    assign _5562 = _1047 ? _1055 : _5560;
    assign _502 = _5562;
    always @(posedge _1038) begin
        if (_1036)
            _5559 <= _1055;
        else
            _5559 <= _502;
    end
    assign _5563 = 9'b000001011;
    assign _5564 = _1062 == _5563;
    assign _5565 = _1059 & _5564;
    assign _5569 = _5565 ? _515 : _5568;
    assign _5571 = _1047 ? _1055 : _5569;
    assign _503 = _5571;
    always @(posedge _1038) begin
        if (_1036)
            _5568 <= _1055;
        else
            _5568 <= _503;
    end
    assign _5572 = 9'b000001010;
    assign _5573 = _1062 == _5572;
    assign _5574 = _1059 & _5573;
    assign _5578 = _5574 ? _515 : _5577;
    assign _5580 = _1047 ? _1055 : _5578;
    assign _504 = _5580;
    always @(posedge _1038) begin
        if (_1036)
            _5577 <= _1055;
        else
            _5577 <= _504;
    end
    assign _5581 = 9'b000001001;
    assign _5582 = _1062 == _5581;
    assign _5583 = _1059 & _5582;
    assign _5587 = _5583 ? _515 : _5586;
    assign _5589 = _1047 ? _1055 : _5587;
    assign _505 = _5589;
    always @(posedge _1038) begin
        if (_1036)
            _5586 <= _1055;
        else
            _5586 <= _505;
    end
    assign _5590 = 9'b000001000;
    assign _5591 = _1062 == _5590;
    assign _5592 = _1059 & _5591;
    assign _5596 = _5592 ? _515 : _5595;
    assign _5598 = _1047 ? _1055 : _5596;
    assign _506 = _5598;
    always @(posedge _1038) begin
        if (_1036)
            _5595 <= _1055;
        else
            _5595 <= _506;
    end
    assign _5599 = 9'b000000111;
    assign _5600 = _1062 == _5599;
    assign _5601 = _1059 & _5600;
    assign _5605 = _5601 ? _515 : _5604;
    assign _5607 = _1047 ? _1055 : _5605;
    assign _507 = _5607;
    always @(posedge _1038) begin
        if (_1036)
            _5604 <= _1055;
        else
            _5604 <= _507;
    end
    assign _5608 = 9'b000000110;
    assign _5609 = _1062 == _5608;
    assign _5610 = _1059 & _5609;
    assign _5614 = _5610 ? _515 : _5613;
    assign _5616 = _1047 ? _1055 : _5614;
    assign _508 = _5616;
    always @(posedge _1038) begin
        if (_1036)
            _5613 <= _1055;
        else
            _5613 <= _508;
    end
    assign _5617 = 9'b000000101;
    assign _5618 = _1062 == _5617;
    assign _5619 = _1059 & _5618;
    assign _5623 = _5619 ? _515 : _5622;
    assign _5625 = _1047 ? _1055 : _5623;
    assign _509 = _5625;
    always @(posedge _1038) begin
        if (_1036)
            _5622 <= _1055;
        else
            _5622 <= _509;
    end
    assign _5626 = 9'b000000100;
    assign _5627 = _1062 == _5626;
    assign _5628 = _1059 & _5627;
    assign _5632 = _5628 ? _515 : _5631;
    assign _5634 = _1047 ? _1055 : _5632;
    assign _510 = _5634;
    always @(posedge _1038) begin
        if (_1036)
            _5631 <= _1055;
        else
            _5631 <= _510;
    end
    assign _5635 = 9'b000000011;
    assign _5636 = _1062 == _5635;
    assign _5637 = _1059 & _5636;
    assign _5641 = _5637 ? _515 : _5640;
    assign _5643 = _1047 ? _1055 : _5641;
    assign _511 = _5643;
    always @(posedge _1038) begin
        if (_1036)
            _5640 <= _1055;
        else
            _5640 <= _511;
    end
    assign _5644 = 9'b000000010;
    assign _5645 = _1062 == _5644;
    assign _5646 = _1059 & _5645;
    assign _5650 = _5646 ? _515 : _5649;
    assign _5652 = _1047 ? _1055 : _5650;
    assign _512 = _5652;
    always @(posedge _1038) begin
        if (_1036)
            _5649 <= _1055;
        else
            _5649 <= _512;
    end
    assign _5653 = 9'b000000001;
    assign _5654 = _1062 == _5653;
    assign _5655 = _1059 & _5654;
    assign _5659 = _5655 ? _515 : _5658;
    assign _5661 = _1047 ? _1055 : _5659;
    assign _513 = _5661;
    always @(posedge _1038) begin
        if (_1036)
            _5658 <= _1055;
        else
            _5658 <= _513;
    end
    assign _515 = y;
    assign _5662 = 9'b000000000;
    assign _5663 = _1062 == _5662;
    assign _5664 = _1059 & _5663;
    assign _5668 = _5664 ? _515 : _5667;
    assign _5670 = _1047 ? _1055 : _5668;
    assign _516 = _5670;
    always @(posedge _1038) begin
        if (_1036)
            _5667 <= _1055;
        else
            _5667 <= _516;
    end
    always @* begin
        case (_10283)
        0:
            _10304 <= _5667;
        1:
            _10304 <= _5658;
        2:
            _10304 <= _5649;
        3:
            _10304 <= _5640;
        4:
            _10304 <= _5631;
        5:
            _10304 <= _5622;
        6:
            _10304 <= _5613;
        7:
            _10304 <= _5604;
        8:
            _10304 <= _5595;
        9:
            _10304 <= _5586;
        10:
            _10304 <= _5577;
        11:
            _10304 <= _5568;
        12:
            _10304 <= _5559;
        13:
            _10304 <= _5550;
        14:
            _10304 <= _5541;
        15:
            _10304 <= _5532;
        16:
            _10304 <= _5523;
        17:
            _10304 <= _5514;
        18:
            _10304 <= _5505;
        19:
            _10304 <= _5496;
        20:
            _10304 <= _5487;
        21:
            _10304 <= _5478;
        22:
            _10304 <= _5469;
        23:
            _10304 <= _5460;
        24:
            _10304 <= _5451;
        25:
            _10304 <= _5442;
        26:
            _10304 <= _5433;
        27:
            _10304 <= _5424;
        28:
            _10304 <= _5415;
        29:
            _10304 <= _5406;
        30:
            _10304 <= _5397;
        31:
            _10304 <= _5388;
        32:
            _10304 <= _5379;
        33:
            _10304 <= _5370;
        34:
            _10304 <= _5361;
        35:
            _10304 <= _5352;
        36:
            _10304 <= _5343;
        37:
            _10304 <= _5334;
        38:
            _10304 <= _5325;
        39:
            _10304 <= _5316;
        40:
            _10304 <= _5307;
        41:
            _10304 <= _5298;
        42:
            _10304 <= _5289;
        43:
            _10304 <= _5280;
        44:
            _10304 <= _5271;
        45:
            _10304 <= _5262;
        46:
            _10304 <= _5253;
        47:
            _10304 <= _5244;
        48:
            _10304 <= _5235;
        49:
            _10304 <= _5226;
        50:
            _10304 <= _5217;
        51:
            _10304 <= _5208;
        52:
            _10304 <= _5199;
        53:
            _10304 <= _5190;
        54:
            _10304 <= _5181;
        55:
            _10304 <= _5172;
        56:
            _10304 <= _5163;
        57:
            _10304 <= _5154;
        58:
            _10304 <= _5145;
        59:
            _10304 <= _5136;
        60:
            _10304 <= _5127;
        61:
            _10304 <= _5118;
        62:
            _10304 <= _5109;
        63:
            _10304 <= _5100;
        64:
            _10304 <= _5091;
        65:
            _10304 <= _5082;
        66:
            _10304 <= _5073;
        67:
            _10304 <= _5064;
        68:
            _10304 <= _5055;
        69:
            _10304 <= _5046;
        70:
            _10304 <= _5037;
        71:
            _10304 <= _5028;
        72:
            _10304 <= _5019;
        73:
            _10304 <= _5010;
        74:
            _10304 <= _5001;
        75:
            _10304 <= _4992;
        76:
            _10304 <= _4983;
        77:
            _10304 <= _4974;
        78:
            _10304 <= _4965;
        79:
            _10304 <= _4956;
        80:
            _10304 <= _4947;
        81:
            _10304 <= _4938;
        82:
            _10304 <= _4929;
        83:
            _10304 <= _4920;
        84:
            _10304 <= _4911;
        85:
            _10304 <= _4902;
        86:
            _10304 <= _4893;
        87:
            _10304 <= _4884;
        88:
            _10304 <= _4875;
        89:
            _10304 <= _4866;
        90:
            _10304 <= _4857;
        91:
            _10304 <= _4848;
        92:
            _10304 <= _4839;
        93:
            _10304 <= _4830;
        94:
            _10304 <= _4821;
        95:
            _10304 <= _4812;
        96:
            _10304 <= _4803;
        97:
            _10304 <= _4794;
        98:
            _10304 <= _4785;
        99:
            _10304 <= _4776;
        100:
            _10304 <= _4767;
        101:
            _10304 <= _4758;
        102:
            _10304 <= _4749;
        103:
            _10304 <= _4740;
        104:
            _10304 <= _4731;
        105:
            _10304 <= _4722;
        106:
            _10304 <= _4713;
        107:
            _10304 <= _4704;
        108:
            _10304 <= _4695;
        109:
            _10304 <= _4686;
        110:
            _10304 <= _4677;
        111:
            _10304 <= _4668;
        112:
            _10304 <= _4659;
        113:
            _10304 <= _4650;
        114:
            _10304 <= _4641;
        115:
            _10304 <= _4632;
        116:
            _10304 <= _4623;
        117:
            _10304 <= _4614;
        118:
            _10304 <= _4605;
        119:
            _10304 <= _4596;
        120:
            _10304 <= _4587;
        121:
            _10304 <= _4578;
        122:
            _10304 <= _4569;
        123:
            _10304 <= _4560;
        124:
            _10304 <= _4551;
        125:
            _10304 <= _4542;
        126:
            _10304 <= _4533;
        127:
            _10304 <= _4524;
        128:
            _10304 <= _4515;
        129:
            _10304 <= _4506;
        130:
            _10304 <= _4497;
        131:
            _10304 <= _4488;
        132:
            _10304 <= _4479;
        133:
            _10304 <= _4470;
        134:
            _10304 <= _4461;
        135:
            _10304 <= _4452;
        136:
            _10304 <= _4443;
        137:
            _10304 <= _4434;
        138:
            _10304 <= _4425;
        139:
            _10304 <= _4416;
        140:
            _10304 <= _4407;
        141:
            _10304 <= _4398;
        142:
            _10304 <= _4389;
        143:
            _10304 <= _4380;
        144:
            _10304 <= _4371;
        145:
            _10304 <= _4362;
        146:
            _10304 <= _4353;
        147:
            _10304 <= _4344;
        148:
            _10304 <= _4335;
        149:
            _10304 <= _4326;
        150:
            _10304 <= _4317;
        151:
            _10304 <= _4308;
        152:
            _10304 <= _4299;
        153:
            _10304 <= _4290;
        154:
            _10304 <= _4281;
        155:
            _10304 <= _4272;
        156:
            _10304 <= _4263;
        157:
            _10304 <= _4254;
        158:
            _10304 <= _4245;
        159:
            _10304 <= _4236;
        160:
            _10304 <= _4227;
        161:
            _10304 <= _4218;
        162:
            _10304 <= _4209;
        163:
            _10304 <= _4200;
        164:
            _10304 <= _4191;
        165:
            _10304 <= _4182;
        166:
            _10304 <= _4173;
        167:
            _10304 <= _4164;
        168:
            _10304 <= _4155;
        169:
            _10304 <= _4146;
        170:
            _10304 <= _4137;
        171:
            _10304 <= _4128;
        172:
            _10304 <= _4119;
        173:
            _10304 <= _4110;
        174:
            _10304 <= _4101;
        175:
            _10304 <= _4092;
        176:
            _10304 <= _4083;
        177:
            _10304 <= _4074;
        178:
            _10304 <= _4065;
        179:
            _10304 <= _4056;
        180:
            _10304 <= _4047;
        181:
            _10304 <= _4038;
        182:
            _10304 <= _4029;
        183:
            _10304 <= _4020;
        184:
            _10304 <= _4011;
        185:
            _10304 <= _4002;
        186:
            _10304 <= _3993;
        187:
            _10304 <= _3984;
        188:
            _10304 <= _3975;
        189:
            _10304 <= _3966;
        190:
            _10304 <= _3957;
        191:
            _10304 <= _3948;
        192:
            _10304 <= _3939;
        193:
            _10304 <= _3930;
        194:
            _10304 <= _3921;
        195:
            _10304 <= _3912;
        196:
            _10304 <= _3903;
        197:
            _10304 <= _3894;
        198:
            _10304 <= _3885;
        199:
            _10304 <= _3876;
        200:
            _10304 <= _3867;
        201:
            _10304 <= _3858;
        202:
            _10304 <= _3849;
        203:
            _10304 <= _3840;
        204:
            _10304 <= _3831;
        205:
            _10304 <= _3822;
        206:
            _10304 <= _3813;
        207:
            _10304 <= _3804;
        208:
            _10304 <= _3795;
        209:
            _10304 <= _3786;
        210:
            _10304 <= _3777;
        211:
            _10304 <= _3768;
        212:
            _10304 <= _3759;
        213:
            _10304 <= _3750;
        214:
            _10304 <= _3741;
        215:
            _10304 <= _3732;
        216:
            _10304 <= _3723;
        217:
            _10304 <= _3714;
        218:
            _10304 <= _3705;
        219:
            _10304 <= _3696;
        220:
            _10304 <= _3687;
        221:
            _10304 <= _3678;
        222:
            _10304 <= _3669;
        223:
            _10304 <= _3660;
        224:
            _10304 <= _3651;
        225:
            _10304 <= _3642;
        226:
            _10304 <= _3633;
        227:
            _10304 <= _3624;
        228:
            _10304 <= _3615;
        229:
            _10304 <= _3606;
        230:
            _10304 <= _3597;
        231:
            _10304 <= _3588;
        232:
            _10304 <= _3579;
        233:
            _10304 <= _3570;
        234:
            _10304 <= _3561;
        235:
            _10304 <= _3552;
        236:
            _10304 <= _3543;
        237:
            _10304 <= _3534;
        238:
            _10304 <= _3525;
        239:
            _10304 <= _3516;
        240:
            _10304 <= _3507;
        241:
            _10304 <= _3498;
        242:
            _10304 <= _3489;
        243:
            _10304 <= _3480;
        244:
            _10304 <= _3471;
        245:
            _10304 <= _3462;
        246:
            _10304 <= _3453;
        247:
            _10304 <= _3444;
        248:
            _10304 <= _3435;
        249:
            _10304 <= _3426;
        250:
            _10304 <= _3417;
        251:
            _10304 <= _3408;
        252:
            _10304 <= _3399;
        253:
            _10304 <= _3390;
        254:
            _10304 <= _3381;
        255:
            _10304 <= _3372;
        256:
            _10304 <= _3363;
        257:
            _10304 <= _3354;
        258:
            _10304 <= _3345;
        259:
            _10304 <= _3336;
        260:
            _10304 <= _3327;
        261:
            _10304 <= _3318;
        262:
            _10304 <= _3309;
        263:
            _10304 <= _3300;
        264:
            _10304 <= _3291;
        265:
            _10304 <= _3282;
        266:
            _10304 <= _3273;
        267:
            _10304 <= _3264;
        268:
            _10304 <= _3255;
        269:
            _10304 <= _3246;
        270:
            _10304 <= _3237;
        271:
            _10304 <= _3228;
        272:
            _10304 <= _3219;
        273:
            _10304 <= _3210;
        274:
            _10304 <= _3201;
        275:
            _10304 <= _3192;
        276:
            _10304 <= _3183;
        277:
            _10304 <= _3174;
        278:
            _10304 <= _3165;
        279:
            _10304 <= _3156;
        280:
            _10304 <= _3147;
        281:
            _10304 <= _3138;
        282:
            _10304 <= _3129;
        283:
            _10304 <= _3120;
        284:
            _10304 <= _3111;
        285:
            _10304 <= _3102;
        286:
            _10304 <= _3093;
        287:
            _10304 <= _3084;
        288:
            _10304 <= _3075;
        289:
            _10304 <= _3066;
        290:
            _10304 <= _3057;
        291:
            _10304 <= _3048;
        292:
            _10304 <= _3039;
        293:
            _10304 <= _3030;
        294:
            _10304 <= _3021;
        295:
            _10304 <= _3012;
        296:
            _10304 <= _3003;
        297:
            _10304 <= _2994;
        298:
            _10304 <= _2985;
        299:
            _10304 <= _2976;
        300:
            _10304 <= _2967;
        301:
            _10304 <= _2958;
        302:
            _10304 <= _2949;
        303:
            _10304 <= _2940;
        304:
            _10304 <= _2931;
        305:
            _10304 <= _2922;
        306:
            _10304 <= _2913;
        307:
            _10304 <= _2904;
        308:
            _10304 <= _2895;
        309:
            _10304 <= _2886;
        310:
            _10304 <= _2877;
        311:
            _10304 <= _2868;
        312:
            _10304 <= _2859;
        313:
            _10304 <= _2850;
        314:
            _10304 <= _2841;
        315:
            _10304 <= _2832;
        316:
            _10304 <= _2823;
        317:
            _10304 <= _2814;
        318:
            _10304 <= _2805;
        319:
            _10304 <= _2796;
        320:
            _10304 <= _2787;
        321:
            _10304 <= _2778;
        322:
            _10304 <= _2769;
        323:
            _10304 <= _2760;
        324:
            _10304 <= _2751;
        325:
            _10304 <= _2742;
        326:
            _10304 <= _2733;
        327:
            _10304 <= _2724;
        328:
            _10304 <= _2715;
        329:
            _10304 <= _2706;
        330:
            _10304 <= _2697;
        331:
            _10304 <= _2688;
        332:
            _10304 <= _2679;
        333:
            _10304 <= _2670;
        334:
            _10304 <= _2661;
        335:
            _10304 <= _2652;
        336:
            _10304 <= _2643;
        337:
            _10304 <= _2634;
        338:
            _10304 <= _2625;
        339:
            _10304 <= _2616;
        340:
            _10304 <= _2607;
        341:
            _10304 <= _2598;
        342:
            _10304 <= _2589;
        343:
            _10304 <= _2580;
        344:
            _10304 <= _2571;
        345:
            _10304 <= _2562;
        346:
            _10304 <= _2553;
        347:
            _10304 <= _2544;
        348:
            _10304 <= _2535;
        349:
            _10304 <= _2526;
        350:
            _10304 <= _2517;
        351:
            _10304 <= _2508;
        352:
            _10304 <= _2499;
        353:
            _10304 <= _2490;
        354:
            _10304 <= _2481;
        355:
            _10304 <= _2472;
        356:
            _10304 <= _2463;
        357:
            _10304 <= _2454;
        358:
            _10304 <= _2445;
        359:
            _10304 <= _2436;
        360:
            _10304 <= _2427;
        361:
            _10304 <= _2418;
        362:
            _10304 <= _2409;
        363:
            _10304 <= _2400;
        364:
            _10304 <= _2391;
        365:
            _10304 <= _2382;
        366:
            _10304 <= _2373;
        367:
            _10304 <= _2364;
        368:
            _10304 <= _2355;
        369:
            _10304 <= _2346;
        370:
            _10304 <= _2337;
        371:
            _10304 <= _2328;
        372:
            _10304 <= _2319;
        373:
            _10304 <= _2310;
        374:
            _10304 <= _2301;
        375:
            _10304 <= _2292;
        376:
            _10304 <= _2283;
        377:
            _10304 <= _2274;
        378:
            _10304 <= _2265;
        379:
            _10304 <= _2256;
        380:
            _10304 <= _2247;
        381:
            _10304 <= _2238;
        382:
            _10304 <= _2229;
        383:
            _10304 <= _2220;
        384:
            _10304 <= _2211;
        385:
            _10304 <= _2202;
        386:
            _10304 <= _2193;
        387:
            _10304 <= _2184;
        388:
            _10304 <= _2175;
        389:
            _10304 <= _2166;
        390:
            _10304 <= _2157;
        391:
            _10304 <= _2148;
        392:
            _10304 <= _2139;
        393:
            _10304 <= _2130;
        394:
            _10304 <= _2121;
        395:
            _10304 <= _2112;
        396:
            _10304 <= _2103;
        397:
            _10304 <= _2094;
        398:
            _10304 <= _2085;
        399:
            _10304 <= _2076;
        400:
            _10304 <= _2067;
        401:
            _10304 <= _2058;
        402:
            _10304 <= _2049;
        403:
            _10304 <= _2040;
        404:
            _10304 <= _2031;
        405:
            _10304 <= _2022;
        406:
            _10304 <= _2013;
        407:
            _10304 <= _2004;
        408:
            _10304 <= _1995;
        409:
            _10304 <= _1986;
        410:
            _10304 <= _1977;
        411:
            _10304 <= _1968;
        412:
            _10304 <= _1959;
        413:
            _10304 <= _1950;
        414:
            _10304 <= _1941;
        415:
            _10304 <= _1932;
        416:
            _10304 <= _1923;
        417:
            _10304 <= _1914;
        418:
            _10304 <= _1905;
        419:
            _10304 <= _1896;
        420:
            _10304 <= _1887;
        421:
            _10304 <= _1878;
        422:
            _10304 <= _1869;
        423:
            _10304 <= _1860;
        424:
            _10304 <= _1851;
        425:
            _10304 <= _1842;
        426:
            _10304 <= _1833;
        427:
            _10304 <= _1824;
        428:
            _10304 <= _1815;
        429:
            _10304 <= _1806;
        430:
            _10304 <= _1797;
        431:
            _10304 <= _1788;
        432:
            _10304 <= _1779;
        433:
            _10304 <= _1770;
        434:
            _10304 <= _1761;
        435:
            _10304 <= _1752;
        436:
            _10304 <= _1743;
        437:
            _10304 <= _1734;
        438:
            _10304 <= _1725;
        439:
            _10304 <= _1716;
        440:
            _10304 <= _1707;
        441:
            _10304 <= _1698;
        442:
            _10304 <= _1689;
        443:
            _10304 <= _1680;
        444:
            _10304 <= _1671;
        445:
            _10304 <= _1662;
        446:
            _10304 <= _1653;
        447:
            _10304 <= _1644;
        448:
            _10304 <= _1635;
        449:
            _10304 <= _1626;
        450:
            _10304 <= _1617;
        451:
            _10304 <= _1608;
        452:
            _10304 <= _1599;
        453:
            _10304 <= _1590;
        454:
            _10304 <= _1581;
        455:
            _10304 <= _1572;
        456:
            _10304 <= _1563;
        457:
            _10304 <= _1554;
        458:
            _10304 <= _1545;
        459:
            _10304 <= _1536;
        460:
            _10304 <= _1527;
        461:
            _10304 <= _1518;
        462:
            _10304 <= _1509;
        463:
            _10304 <= _1500;
        464:
            _10304 <= _1491;
        465:
            _10304 <= _1482;
        466:
            _10304 <= _1473;
        467:
            _10304 <= _1464;
        468:
            _10304 <= _1455;
        469:
            _10304 <= _1446;
        470:
            _10304 <= _1437;
        471:
            _10304 <= _1428;
        472:
            _10304 <= _1419;
        473:
            _10304 <= _1410;
        474:
            _10304 <= _1401;
        475:
            _10304 <= _1392;
        476:
            _10304 <= _1383;
        477:
            _10304 <= _1374;
        478:
            _10304 <= _1365;
        479:
            _10304 <= _1356;
        480:
            _10304 <= _1347;
        481:
            _10304 <= _1338;
        482:
            _10304 <= _1329;
        483:
            _10304 <= _1320;
        484:
            _10304 <= _1311;
        485:
            _10304 <= _1302;
        486:
            _10304 <= _1293;
        487:
            _10304 <= _1284;
        488:
            _10304 <= _1275;
        489:
            _10304 <= _1266;
        490:
            _10304 <= _1257;
        491:
            _10304 <= _1248;
        492:
            _10304 <= _1239;
        493:
            _10304 <= _1230;
        494:
            _10304 <= _1221;
        495:
            _10304 <= _1212;
        496:
            _10304 <= _1203;
        497:
            _10304 <= _1194;
        498:
            _10304 <= _1185;
        499:
            _10304 <= _1176;
        500:
            _10304 <= _1167;
        501:
            _10304 <= _1158;
        502:
            _10304 <= _1149;
        503:
            _10304 <= _1140;
        504:
            _10304 <= _1131;
        505:
            _10304 <= _1122;
        506:
            _10304 <= _1113;
        507:
            _10304 <= _1104;
        508:
            _10304 <= _1095;
        509:
            _10304 <= _1086;
        510:
            _10304 <= _1077;
        default:
            _10304 <= _1068;
        endcase
    end
    assign _10306 = _10304 < _10305;
    assign _10307 = ~ _10306;
    assign _10310 = _10307 ? _10309 : _10308;
    assign _10312 = _10310 + _10311;
    assign _10300 = _10295 - _10296;
    assign _10299 = _10296 - _10295;
    always @* begin
        case (_10291)
        0:
            _10296 <= _10275;
        1:
            _10296 <= _10266;
        2:
            _10296 <= _10257;
        3:
            _10296 <= _10248;
        4:
            _10296 <= _10239;
        5:
            _10296 <= _10230;
        6:
            _10296 <= _10221;
        7:
            _10296 <= _10212;
        8:
            _10296 <= _10203;
        9:
            _10296 <= _10194;
        10:
            _10296 <= _10185;
        11:
            _10296 <= _10176;
        12:
            _10296 <= _10167;
        13:
            _10296 <= _10158;
        14:
            _10296 <= _10149;
        15:
            _10296 <= _10140;
        16:
            _10296 <= _10131;
        17:
            _10296 <= _10122;
        18:
            _10296 <= _10113;
        19:
            _10296 <= _10104;
        20:
            _10296 <= _10095;
        21:
            _10296 <= _10086;
        22:
            _10296 <= _10077;
        23:
            _10296 <= _10068;
        24:
            _10296 <= _10059;
        25:
            _10296 <= _10050;
        26:
            _10296 <= _10041;
        27:
            _10296 <= _10032;
        28:
            _10296 <= _10023;
        29:
            _10296 <= _10014;
        30:
            _10296 <= _10005;
        31:
            _10296 <= _9996;
        32:
            _10296 <= _9987;
        33:
            _10296 <= _9978;
        34:
            _10296 <= _9969;
        35:
            _10296 <= _9960;
        36:
            _10296 <= _9951;
        37:
            _10296 <= _9942;
        38:
            _10296 <= _9933;
        39:
            _10296 <= _9924;
        40:
            _10296 <= _9915;
        41:
            _10296 <= _9906;
        42:
            _10296 <= _9897;
        43:
            _10296 <= _9888;
        44:
            _10296 <= _9879;
        45:
            _10296 <= _9870;
        46:
            _10296 <= _9861;
        47:
            _10296 <= _9852;
        48:
            _10296 <= _9843;
        49:
            _10296 <= _9834;
        50:
            _10296 <= _9825;
        51:
            _10296 <= _9816;
        52:
            _10296 <= _9807;
        53:
            _10296 <= _9798;
        54:
            _10296 <= _9789;
        55:
            _10296 <= _9780;
        56:
            _10296 <= _9771;
        57:
            _10296 <= _9762;
        58:
            _10296 <= _9753;
        59:
            _10296 <= _9744;
        60:
            _10296 <= _9735;
        61:
            _10296 <= _9726;
        62:
            _10296 <= _9717;
        63:
            _10296 <= _9708;
        64:
            _10296 <= _9699;
        65:
            _10296 <= _9690;
        66:
            _10296 <= _9681;
        67:
            _10296 <= _9672;
        68:
            _10296 <= _9663;
        69:
            _10296 <= _9654;
        70:
            _10296 <= _9645;
        71:
            _10296 <= _9636;
        72:
            _10296 <= _9627;
        73:
            _10296 <= _9618;
        74:
            _10296 <= _9609;
        75:
            _10296 <= _9600;
        76:
            _10296 <= _9591;
        77:
            _10296 <= _9582;
        78:
            _10296 <= _9573;
        79:
            _10296 <= _9564;
        80:
            _10296 <= _9555;
        81:
            _10296 <= _9546;
        82:
            _10296 <= _9537;
        83:
            _10296 <= _9528;
        84:
            _10296 <= _9519;
        85:
            _10296 <= _9510;
        86:
            _10296 <= _9501;
        87:
            _10296 <= _9492;
        88:
            _10296 <= _9483;
        89:
            _10296 <= _9474;
        90:
            _10296 <= _9465;
        91:
            _10296 <= _9456;
        92:
            _10296 <= _9447;
        93:
            _10296 <= _9438;
        94:
            _10296 <= _9429;
        95:
            _10296 <= _9420;
        96:
            _10296 <= _9411;
        97:
            _10296 <= _9402;
        98:
            _10296 <= _9393;
        99:
            _10296 <= _9384;
        100:
            _10296 <= _9375;
        101:
            _10296 <= _9366;
        102:
            _10296 <= _9357;
        103:
            _10296 <= _9348;
        104:
            _10296 <= _9339;
        105:
            _10296 <= _9330;
        106:
            _10296 <= _9321;
        107:
            _10296 <= _9312;
        108:
            _10296 <= _9303;
        109:
            _10296 <= _9294;
        110:
            _10296 <= _9285;
        111:
            _10296 <= _9276;
        112:
            _10296 <= _9267;
        113:
            _10296 <= _9258;
        114:
            _10296 <= _9249;
        115:
            _10296 <= _9240;
        116:
            _10296 <= _9231;
        117:
            _10296 <= _9222;
        118:
            _10296 <= _9213;
        119:
            _10296 <= _9204;
        120:
            _10296 <= _9195;
        121:
            _10296 <= _9186;
        122:
            _10296 <= _9177;
        123:
            _10296 <= _9168;
        124:
            _10296 <= _9159;
        125:
            _10296 <= _9150;
        126:
            _10296 <= _9141;
        127:
            _10296 <= _9132;
        128:
            _10296 <= _9123;
        129:
            _10296 <= _9114;
        130:
            _10296 <= _9105;
        131:
            _10296 <= _9096;
        132:
            _10296 <= _9087;
        133:
            _10296 <= _9078;
        134:
            _10296 <= _9069;
        135:
            _10296 <= _9060;
        136:
            _10296 <= _9051;
        137:
            _10296 <= _9042;
        138:
            _10296 <= _9033;
        139:
            _10296 <= _9024;
        140:
            _10296 <= _9015;
        141:
            _10296 <= _9006;
        142:
            _10296 <= _8997;
        143:
            _10296 <= _8988;
        144:
            _10296 <= _8979;
        145:
            _10296 <= _8970;
        146:
            _10296 <= _8961;
        147:
            _10296 <= _8952;
        148:
            _10296 <= _8943;
        149:
            _10296 <= _8934;
        150:
            _10296 <= _8925;
        151:
            _10296 <= _8916;
        152:
            _10296 <= _8907;
        153:
            _10296 <= _8898;
        154:
            _10296 <= _8889;
        155:
            _10296 <= _8880;
        156:
            _10296 <= _8871;
        157:
            _10296 <= _8862;
        158:
            _10296 <= _8853;
        159:
            _10296 <= _8844;
        160:
            _10296 <= _8835;
        161:
            _10296 <= _8826;
        162:
            _10296 <= _8817;
        163:
            _10296 <= _8808;
        164:
            _10296 <= _8799;
        165:
            _10296 <= _8790;
        166:
            _10296 <= _8781;
        167:
            _10296 <= _8772;
        168:
            _10296 <= _8763;
        169:
            _10296 <= _8754;
        170:
            _10296 <= _8745;
        171:
            _10296 <= _8736;
        172:
            _10296 <= _8727;
        173:
            _10296 <= _8718;
        174:
            _10296 <= _8709;
        175:
            _10296 <= _8700;
        176:
            _10296 <= _8691;
        177:
            _10296 <= _8682;
        178:
            _10296 <= _8673;
        179:
            _10296 <= _8664;
        180:
            _10296 <= _8655;
        181:
            _10296 <= _8646;
        182:
            _10296 <= _8637;
        183:
            _10296 <= _8628;
        184:
            _10296 <= _8619;
        185:
            _10296 <= _8610;
        186:
            _10296 <= _8601;
        187:
            _10296 <= _8592;
        188:
            _10296 <= _8583;
        189:
            _10296 <= _8574;
        190:
            _10296 <= _8565;
        191:
            _10296 <= _8556;
        192:
            _10296 <= _8547;
        193:
            _10296 <= _8538;
        194:
            _10296 <= _8529;
        195:
            _10296 <= _8520;
        196:
            _10296 <= _8511;
        197:
            _10296 <= _8502;
        198:
            _10296 <= _8493;
        199:
            _10296 <= _8484;
        200:
            _10296 <= _8475;
        201:
            _10296 <= _8466;
        202:
            _10296 <= _8457;
        203:
            _10296 <= _8448;
        204:
            _10296 <= _8439;
        205:
            _10296 <= _8430;
        206:
            _10296 <= _8421;
        207:
            _10296 <= _8412;
        208:
            _10296 <= _8403;
        209:
            _10296 <= _8394;
        210:
            _10296 <= _8385;
        211:
            _10296 <= _8376;
        212:
            _10296 <= _8367;
        213:
            _10296 <= _8358;
        214:
            _10296 <= _8349;
        215:
            _10296 <= _8340;
        216:
            _10296 <= _8331;
        217:
            _10296 <= _8322;
        218:
            _10296 <= _8313;
        219:
            _10296 <= _8304;
        220:
            _10296 <= _8295;
        221:
            _10296 <= _8286;
        222:
            _10296 <= _8277;
        223:
            _10296 <= _8268;
        224:
            _10296 <= _8259;
        225:
            _10296 <= _8250;
        226:
            _10296 <= _8241;
        227:
            _10296 <= _8232;
        228:
            _10296 <= _8223;
        229:
            _10296 <= _8214;
        230:
            _10296 <= _8205;
        231:
            _10296 <= _8196;
        232:
            _10296 <= _8187;
        233:
            _10296 <= _8178;
        234:
            _10296 <= _8169;
        235:
            _10296 <= _8160;
        236:
            _10296 <= _8151;
        237:
            _10296 <= _8142;
        238:
            _10296 <= _8133;
        239:
            _10296 <= _8124;
        240:
            _10296 <= _8115;
        241:
            _10296 <= _8106;
        242:
            _10296 <= _8097;
        243:
            _10296 <= _8088;
        244:
            _10296 <= _8079;
        245:
            _10296 <= _8070;
        246:
            _10296 <= _8061;
        247:
            _10296 <= _8052;
        248:
            _10296 <= _8043;
        249:
            _10296 <= _8034;
        250:
            _10296 <= _8025;
        251:
            _10296 <= _8016;
        252:
            _10296 <= _8007;
        253:
            _10296 <= _7998;
        254:
            _10296 <= _7989;
        255:
            _10296 <= _7980;
        256:
            _10296 <= _7971;
        257:
            _10296 <= _7962;
        258:
            _10296 <= _7953;
        259:
            _10296 <= _7944;
        260:
            _10296 <= _7935;
        261:
            _10296 <= _7926;
        262:
            _10296 <= _7917;
        263:
            _10296 <= _7908;
        264:
            _10296 <= _7899;
        265:
            _10296 <= _7890;
        266:
            _10296 <= _7881;
        267:
            _10296 <= _7872;
        268:
            _10296 <= _7863;
        269:
            _10296 <= _7854;
        270:
            _10296 <= _7845;
        271:
            _10296 <= _7836;
        272:
            _10296 <= _7827;
        273:
            _10296 <= _7818;
        274:
            _10296 <= _7809;
        275:
            _10296 <= _7800;
        276:
            _10296 <= _7791;
        277:
            _10296 <= _7782;
        278:
            _10296 <= _7773;
        279:
            _10296 <= _7764;
        280:
            _10296 <= _7755;
        281:
            _10296 <= _7746;
        282:
            _10296 <= _7737;
        283:
            _10296 <= _7728;
        284:
            _10296 <= _7719;
        285:
            _10296 <= _7710;
        286:
            _10296 <= _7701;
        287:
            _10296 <= _7692;
        288:
            _10296 <= _7683;
        289:
            _10296 <= _7674;
        290:
            _10296 <= _7665;
        291:
            _10296 <= _7656;
        292:
            _10296 <= _7647;
        293:
            _10296 <= _7638;
        294:
            _10296 <= _7629;
        295:
            _10296 <= _7620;
        296:
            _10296 <= _7611;
        297:
            _10296 <= _7602;
        298:
            _10296 <= _7593;
        299:
            _10296 <= _7584;
        300:
            _10296 <= _7575;
        301:
            _10296 <= _7566;
        302:
            _10296 <= _7557;
        303:
            _10296 <= _7548;
        304:
            _10296 <= _7539;
        305:
            _10296 <= _7530;
        306:
            _10296 <= _7521;
        307:
            _10296 <= _7512;
        308:
            _10296 <= _7503;
        309:
            _10296 <= _7494;
        310:
            _10296 <= _7485;
        311:
            _10296 <= _7476;
        312:
            _10296 <= _7467;
        313:
            _10296 <= _7458;
        314:
            _10296 <= _7449;
        315:
            _10296 <= _7440;
        316:
            _10296 <= _7431;
        317:
            _10296 <= _7422;
        318:
            _10296 <= _7413;
        319:
            _10296 <= _7404;
        320:
            _10296 <= _7395;
        321:
            _10296 <= _7386;
        322:
            _10296 <= _7377;
        323:
            _10296 <= _7368;
        324:
            _10296 <= _7359;
        325:
            _10296 <= _7350;
        326:
            _10296 <= _7341;
        327:
            _10296 <= _7332;
        328:
            _10296 <= _7323;
        329:
            _10296 <= _7314;
        330:
            _10296 <= _7305;
        331:
            _10296 <= _7296;
        332:
            _10296 <= _7287;
        333:
            _10296 <= _7278;
        334:
            _10296 <= _7269;
        335:
            _10296 <= _7260;
        336:
            _10296 <= _7251;
        337:
            _10296 <= _7242;
        338:
            _10296 <= _7233;
        339:
            _10296 <= _7224;
        340:
            _10296 <= _7215;
        341:
            _10296 <= _7206;
        342:
            _10296 <= _7197;
        343:
            _10296 <= _7188;
        344:
            _10296 <= _7179;
        345:
            _10296 <= _7170;
        346:
            _10296 <= _7161;
        347:
            _10296 <= _7152;
        348:
            _10296 <= _7143;
        349:
            _10296 <= _7134;
        350:
            _10296 <= _7125;
        351:
            _10296 <= _7116;
        352:
            _10296 <= _7107;
        353:
            _10296 <= _7098;
        354:
            _10296 <= _7089;
        355:
            _10296 <= _7080;
        356:
            _10296 <= _7071;
        357:
            _10296 <= _7062;
        358:
            _10296 <= _7053;
        359:
            _10296 <= _7044;
        360:
            _10296 <= _7035;
        361:
            _10296 <= _7026;
        362:
            _10296 <= _7017;
        363:
            _10296 <= _7008;
        364:
            _10296 <= _6999;
        365:
            _10296 <= _6990;
        366:
            _10296 <= _6981;
        367:
            _10296 <= _6972;
        368:
            _10296 <= _6963;
        369:
            _10296 <= _6954;
        370:
            _10296 <= _6945;
        371:
            _10296 <= _6936;
        372:
            _10296 <= _6927;
        373:
            _10296 <= _6918;
        374:
            _10296 <= _6909;
        375:
            _10296 <= _6900;
        376:
            _10296 <= _6891;
        377:
            _10296 <= _6882;
        378:
            _10296 <= _6873;
        379:
            _10296 <= _6864;
        380:
            _10296 <= _6855;
        381:
            _10296 <= _6846;
        382:
            _10296 <= _6837;
        383:
            _10296 <= _6828;
        384:
            _10296 <= _6819;
        385:
            _10296 <= _6810;
        386:
            _10296 <= _6801;
        387:
            _10296 <= _6792;
        388:
            _10296 <= _6783;
        389:
            _10296 <= _6774;
        390:
            _10296 <= _6765;
        391:
            _10296 <= _6756;
        392:
            _10296 <= _6747;
        393:
            _10296 <= _6738;
        394:
            _10296 <= _6729;
        395:
            _10296 <= _6720;
        396:
            _10296 <= _6711;
        397:
            _10296 <= _6702;
        398:
            _10296 <= _6693;
        399:
            _10296 <= _6684;
        400:
            _10296 <= _6675;
        401:
            _10296 <= _6666;
        402:
            _10296 <= _6657;
        403:
            _10296 <= _6648;
        404:
            _10296 <= _6639;
        405:
            _10296 <= _6630;
        406:
            _10296 <= _6621;
        407:
            _10296 <= _6612;
        408:
            _10296 <= _6603;
        409:
            _10296 <= _6594;
        410:
            _10296 <= _6585;
        411:
            _10296 <= _6576;
        412:
            _10296 <= _6567;
        413:
            _10296 <= _6558;
        414:
            _10296 <= _6549;
        415:
            _10296 <= _6540;
        416:
            _10296 <= _6531;
        417:
            _10296 <= _6522;
        418:
            _10296 <= _6513;
        419:
            _10296 <= _6504;
        420:
            _10296 <= _6495;
        421:
            _10296 <= _6486;
        422:
            _10296 <= _6477;
        423:
            _10296 <= _6468;
        424:
            _10296 <= _6459;
        425:
            _10296 <= _6450;
        426:
            _10296 <= _6441;
        427:
            _10296 <= _6432;
        428:
            _10296 <= _6423;
        429:
            _10296 <= _6414;
        430:
            _10296 <= _6405;
        431:
            _10296 <= _6396;
        432:
            _10296 <= _6387;
        433:
            _10296 <= _6378;
        434:
            _10296 <= _6369;
        435:
            _10296 <= _6360;
        436:
            _10296 <= _6351;
        437:
            _10296 <= _6342;
        438:
            _10296 <= _6333;
        439:
            _10296 <= _6324;
        440:
            _10296 <= _6315;
        441:
            _10296 <= _6306;
        442:
            _10296 <= _6297;
        443:
            _10296 <= _6288;
        444:
            _10296 <= _6279;
        445:
            _10296 <= _6270;
        446:
            _10296 <= _6261;
        447:
            _10296 <= _6252;
        448:
            _10296 <= _6243;
        449:
            _10296 <= _6234;
        450:
            _10296 <= _6225;
        451:
            _10296 <= _6216;
        452:
            _10296 <= _6207;
        453:
            _10296 <= _6198;
        454:
            _10296 <= _6189;
        455:
            _10296 <= _6180;
        456:
            _10296 <= _6171;
        457:
            _10296 <= _6162;
        458:
            _10296 <= _6153;
        459:
            _10296 <= _6144;
        460:
            _10296 <= _6135;
        461:
            _10296 <= _6126;
        462:
            _10296 <= _6117;
        463:
            _10296 <= _6108;
        464:
            _10296 <= _6099;
        465:
            _10296 <= _6090;
        466:
            _10296 <= _6081;
        467:
            _10296 <= _6072;
        468:
            _10296 <= _6063;
        469:
            _10296 <= _6054;
        470:
            _10296 <= _6045;
        471:
            _10296 <= _6036;
        472:
            _10296 <= _6027;
        473:
            _10296 <= _6018;
        474:
            _10296 <= _6009;
        475:
            _10296 <= _6000;
        476:
            _10296 <= _5991;
        477:
            _10296 <= _5982;
        478:
            _10296 <= _5973;
        479:
            _10296 <= _5964;
        480:
            _10296 <= _5955;
        481:
            _10296 <= _5946;
        482:
            _10296 <= _5937;
        483:
            _10296 <= _5928;
        484:
            _10296 <= _5919;
        485:
            _10296 <= _5910;
        486:
            _10296 <= _5901;
        487:
            _10296 <= _5892;
        488:
            _10296 <= _5883;
        489:
            _10296 <= _5874;
        490:
            _10296 <= _5865;
        491:
            _10296 <= _5856;
        492:
            _10296 <= _5847;
        493:
            _10296 <= _5838;
        494:
            _10296 <= _5829;
        495:
            _10296 <= _5820;
        496:
            _10296 <= _5811;
        497:
            _10296 <= _5802;
        498:
            _10296 <= _5793;
        499:
            _10296 <= _5784;
        500:
            _10296 <= _5775;
        501:
            _10296 <= _5766;
        502:
            _10296 <= _5757;
        503:
            _10296 <= _5748;
        504:
            _10296 <= _5739;
        505:
            _10296 <= _5730;
        506:
            _10296 <= _5721;
        507:
            _10296 <= _5712;
        508:
            _10296 <= _5703;
        509:
            _10296 <= _5694;
        510:
            _10296 <= _5685;
        default:
            _10296 <= _5676;
        endcase
    end
    assign _5672 = _1062 == _1063;
    assign _5673 = _1059 & _5672;
    assign _5677 = _5673 ? _1029 : _5676;
    assign _5679 = _1047 ? _1055 : _5677;
    assign _517 = _5679;
    always @(posedge _1038) begin
        if (_1036)
            _5676 <= _1055;
        else
            _5676 <= _517;
    end
    assign _5681 = _1062 == _1072;
    assign _5682 = _1059 & _5681;
    assign _5686 = _5682 ? _1029 : _5685;
    assign _5688 = _1047 ? _1055 : _5686;
    assign _518 = _5688;
    always @(posedge _1038) begin
        if (_1036)
            _5685 <= _1055;
        else
            _5685 <= _518;
    end
    assign _5690 = _1062 == _1081;
    assign _5691 = _1059 & _5690;
    assign _5695 = _5691 ? _1029 : _5694;
    assign _5697 = _1047 ? _1055 : _5695;
    assign _519 = _5697;
    always @(posedge _1038) begin
        if (_1036)
            _5694 <= _1055;
        else
            _5694 <= _519;
    end
    assign _5699 = _1062 == _1090;
    assign _5700 = _1059 & _5699;
    assign _5704 = _5700 ? _1029 : _5703;
    assign _5706 = _1047 ? _1055 : _5704;
    assign _520 = _5706;
    always @(posedge _1038) begin
        if (_1036)
            _5703 <= _1055;
        else
            _5703 <= _520;
    end
    assign _5708 = _1062 == _1099;
    assign _5709 = _1059 & _5708;
    assign _5713 = _5709 ? _1029 : _5712;
    assign _5715 = _1047 ? _1055 : _5713;
    assign _521 = _5715;
    always @(posedge _1038) begin
        if (_1036)
            _5712 <= _1055;
        else
            _5712 <= _521;
    end
    assign _5717 = _1062 == _1108;
    assign _5718 = _1059 & _5717;
    assign _5722 = _5718 ? _1029 : _5721;
    assign _5724 = _1047 ? _1055 : _5722;
    assign _522 = _5724;
    always @(posedge _1038) begin
        if (_1036)
            _5721 <= _1055;
        else
            _5721 <= _522;
    end
    assign _5726 = _1062 == _1117;
    assign _5727 = _1059 & _5726;
    assign _5731 = _5727 ? _1029 : _5730;
    assign _5733 = _1047 ? _1055 : _5731;
    assign _523 = _5733;
    always @(posedge _1038) begin
        if (_1036)
            _5730 <= _1055;
        else
            _5730 <= _523;
    end
    assign _5735 = _1062 == _1126;
    assign _5736 = _1059 & _5735;
    assign _5740 = _5736 ? _1029 : _5739;
    assign _5742 = _1047 ? _1055 : _5740;
    assign _524 = _5742;
    always @(posedge _1038) begin
        if (_1036)
            _5739 <= _1055;
        else
            _5739 <= _524;
    end
    assign _5744 = _1062 == _1135;
    assign _5745 = _1059 & _5744;
    assign _5749 = _5745 ? _1029 : _5748;
    assign _5751 = _1047 ? _1055 : _5749;
    assign _525 = _5751;
    always @(posedge _1038) begin
        if (_1036)
            _5748 <= _1055;
        else
            _5748 <= _525;
    end
    assign _5753 = _1062 == _1144;
    assign _5754 = _1059 & _5753;
    assign _5758 = _5754 ? _1029 : _5757;
    assign _5760 = _1047 ? _1055 : _5758;
    assign _526 = _5760;
    always @(posedge _1038) begin
        if (_1036)
            _5757 <= _1055;
        else
            _5757 <= _526;
    end
    assign _5762 = _1062 == _1153;
    assign _5763 = _1059 & _5762;
    assign _5767 = _5763 ? _1029 : _5766;
    assign _5769 = _1047 ? _1055 : _5767;
    assign _527 = _5769;
    always @(posedge _1038) begin
        if (_1036)
            _5766 <= _1055;
        else
            _5766 <= _527;
    end
    assign _5771 = _1062 == _1162;
    assign _5772 = _1059 & _5771;
    assign _5776 = _5772 ? _1029 : _5775;
    assign _5778 = _1047 ? _1055 : _5776;
    assign _528 = _5778;
    always @(posedge _1038) begin
        if (_1036)
            _5775 <= _1055;
        else
            _5775 <= _528;
    end
    assign _5780 = _1062 == _1171;
    assign _5781 = _1059 & _5780;
    assign _5785 = _5781 ? _1029 : _5784;
    assign _5787 = _1047 ? _1055 : _5785;
    assign _529 = _5787;
    always @(posedge _1038) begin
        if (_1036)
            _5784 <= _1055;
        else
            _5784 <= _529;
    end
    assign _5789 = _1062 == _1180;
    assign _5790 = _1059 & _5789;
    assign _5794 = _5790 ? _1029 : _5793;
    assign _5796 = _1047 ? _1055 : _5794;
    assign _530 = _5796;
    always @(posedge _1038) begin
        if (_1036)
            _5793 <= _1055;
        else
            _5793 <= _530;
    end
    assign _5798 = _1062 == _1189;
    assign _5799 = _1059 & _5798;
    assign _5803 = _5799 ? _1029 : _5802;
    assign _5805 = _1047 ? _1055 : _5803;
    assign _531 = _5805;
    always @(posedge _1038) begin
        if (_1036)
            _5802 <= _1055;
        else
            _5802 <= _531;
    end
    assign _5807 = _1062 == _1198;
    assign _5808 = _1059 & _5807;
    assign _5812 = _5808 ? _1029 : _5811;
    assign _5814 = _1047 ? _1055 : _5812;
    assign _532 = _5814;
    always @(posedge _1038) begin
        if (_1036)
            _5811 <= _1055;
        else
            _5811 <= _532;
    end
    assign _5816 = _1062 == _1207;
    assign _5817 = _1059 & _5816;
    assign _5821 = _5817 ? _1029 : _5820;
    assign _5823 = _1047 ? _1055 : _5821;
    assign _533 = _5823;
    always @(posedge _1038) begin
        if (_1036)
            _5820 <= _1055;
        else
            _5820 <= _533;
    end
    assign _5825 = _1062 == _1216;
    assign _5826 = _1059 & _5825;
    assign _5830 = _5826 ? _1029 : _5829;
    assign _5832 = _1047 ? _1055 : _5830;
    assign _534 = _5832;
    always @(posedge _1038) begin
        if (_1036)
            _5829 <= _1055;
        else
            _5829 <= _534;
    end
    assign _5834 = _1062 == _1225;
    assign _5835 = _1059 & _5834;
    assign _5839 = _5835 ? _1029 : _5838;
    assign _5841 = _1047 ? _1055 : _5839;
    assign _535 = _5841;
    always @(posedge _1038) begin
        if (_1036)
            _5838 <= _1055;
        else
            _5838 <= _535;
    end
    assign _5843 = _1062 == _1234;
    assign _5844 = _1059 & _5843;
    assign _5848 = _5844 ? _1029 : _5847;
    assign _5850 = _1047 ? _1055 : _5848;
    assign _536 = _5850;
    always @(posedge _1038) begin
        if (_1036)
            _5847 <= _1055;
        else
            _5847 <= _536;
    end
    assign _5852 = _1062 == _1243;
    assign _5853 = _1059 & _5852;
    assign _5857 = _5853 ? _1029 : _5856;
    assign _5859 = _1047 ? _1055 : _5857;
    assign _537 = _5859;
    always @(posedge _1038) begin
        if (_1036)
            _5856 <= _1055;
        else
            _5856 <= _537;
    end
    assign _5861 = _1062 == _1252;
    assign _5862 = _1059 & _5861;
    assign _5866 = _5862 ? _1029 : _5865;
    assign _5868 = _1047 ? _1055 : _5866;
    assign _538 = _5868;
    always @(posedge _1038) begin
        if (_1036)
            _5865 <= _1055;
        else
            _5865 <= _538;
    end
    assign _5870 = _1062 == _1261;
    assign _5871 = _1059 & _5870;
    assign _5875 = _5871 ? _1029 : _5874;
    assign _5877 = _1047 ? _1055 : _5875;
    assign _539 = _5877;
    always @(posedge _1038) begin
        if (_1036)
            _5874 <= _1055;
        else
            _5874 <= _539;
    end
    assign _5879 = _1062 == _1270;
    assign _5880 = _1059 & _5879;
    assign _5884 = _5880 ? _1029 : _5883;
    assign _5886 = _1047 ? _1055 : _5884;
    assign _540 = _5886;
    always @(posedge _1038) begin
        if (_1036)
            _5883 <= _1055;
        else
            _5883 <= _540;
    end
    assign _5888 = _1062 == _1279;
    assign _5889 = _1059 & _5888;
    assign _5893 = _5889 ? _1029 : _5892;
    assign _5895 = _1047 ? _1055 : _5893;
    assign _541 = _5895;
    always @(posedge _1038) begin
        if (_1036)
            _5892 <= _1055;
        else
            _5892 <= _541;
    end
    assign _5897 = _1062 == _1288;
    assign _5898 = _1059 & _5897;
    assign _5902 = _5898 ? _1029 : _5901;
    assign _5904 = _1047 ? _1055 : _5902;
    assign _542 = _5904;
    always @(posedge _1038) begin
        if (_1036)
            _5901 <= _1055;
        else
            _5901 <= _542;
    end
    assign _5906 = _1062 == _1297;
    assign _5907 = _1059 & _5906;
    assign _5911 = _5907 ? _1029 : _5910;
    assign _5913 = _1047 ? _1055 : _5911;
    assign _543 = _5913;
    always @(posedge _1038) begin
        if (_1036)
            _5910 <= _1055;
        else
            _5910 <= _543;
    end
    assign _5915 = _1062 == _1306;
    assign _5916 = _1059 & _5915;
    assign _5920 = _5916 ? _1029 : _5919;
    assign _5922 = _1047 ? _1055 : _5920;
    assign _544 = _5922;
    always @(posedge _1038) begin
        if (_1036)
            _5919 <= _1055;
        else
            _5919 <= _544;
    end
    assign _5924 = _1062 == _1315;
    assign _5925 = _1059 & _5924;
    assign _5929 = _5925 ? _1029 : _5928;
    assign _5931 = _1047 ? _1055 : _5929;
    assign _545 = _5931;
    always @(posedge _1038) begin
        if (_1036)
            _5928 <= _1055;
        else
            _5928 <= _545;
    end
    assign _5933 = _1062 == _1324;
    assign _5934 = _1059 & _5933;
    assign _5938 = _5934 ? _1029 : _5937;
    assign _5940 = _1047 ? _1055 : _5938;
    assign _546 = _5940;
    always @(posedge _1038) begin
        if (_1036)
            _5937 <= _1055;
        else
            _5937 <= _546;
    end
    assign _5942 = _1062 == _1333;
    assign _5943 = _1059 & _5942;
    assign _5947 = _5943 ? _1029 : _5946;
    assign _5949 = _1047 ? _1055 : _5947;
    assign _547 = _5949;
    always @(posedge _1038) begin
        if (_1036)
            _5946 <= _1055;
        else
            _5946 <= _547;
    end
    assign _5951 = _1062 == _1342;
    assign _5952 = _1059 & _5951;
    assign _5956 = _5952 ? _1029 : _5955;
    assign _5958 = _1047 ? _1055 : _5956;
    assign _548 = _5958;
    always @(posedge _1038) begin
        if (_1036)
            _5955 <= _1055;
        else
            _5955 <= _548;
    end
    assign _5960 = _1062 == _1351;
    assign _5961 = _1059 & _5960;
    assign _5965 = _5961 ? _1029 : _5964;
    assign _5967 = _1047 ? _1055 : _5965;
    assign _549 = _5967;
    always @(posedge _1038) begin
        if (_1036)
            _5964 <= _1055;
        else
            _5964 <= _549;
    end
    assign _5969 = _1062 == _1360;
    assign _5970 = _1059 & _5969;
    assign _5974 = _5970 ? _1029 : _5973;
    assign _5976 = _1047 ? _1055 : _5974;
    assign _550 = _5976;
    always @(posedge _1038) begin
        if (_1036)
            _5973 <= _1055;
        else
            _5973 <= _550;
    end
    assign _5978 = _1062 == _1369;
    assign _5979 = _1059 & _5978;
    assign _5983 = _5979 ? _1029 : _5982;
    assign _5985 = _1047 ? _1055 : _5983;
    assign _551 = _5985;
    always @(posedge _1038) begin
        if (_1036)
            _5982 <= _1055;
        else
            _5982 <= _551;
    end
    assign _5987 = _1062 == _1378;
    assign _5988 = _1059 & _5987;
    assign _5992 = _5988 ? _1029 : _5991;
    assign _5994 = _1047 ? _1055 : _5992;
    assign _552 = _5994;
    always @(posedge _1038) begin
        if (_1036)
            _5991 <= _1055;
        else
            _5991 <= _552;
    end
    assign _5996 = _1062 == _1387;
    assign _5997 = _1059 & _5996;
    assign _6001 = _5997 ? _1029 : _6000;
    assign _6003 = _1047 ? _1055 : _6001;
    assign _553 = _6003;
    always @(posedge _1038) begin
        if (_1036)
            _6000 <= _1055;
        else
            _6000 <= _553;
    end
    assign _6005 = _1062 == _1396;
    assign _6006 = _1059 & _6005;
    assign _6010 = _6006 ? _1029 : _6009;
    assign _6012 = _1047 ? _1055 : _6010;
    assign _554 = _6012;
    always @(posedge _1038) begin
        if (_1036)
            _6009 <= _1055;
        else
            _6009 <= _554;
    end
    assign _6014 = _1062 == _1405;
    assign _6015 = _1059 & _6014;
    assign _6019 = _6015 ? _1029 : _6018;
    assign _6021 = _1047 ? _1055 : _6019;
    assign _555 = _6021;
    always @(posedge _1038) begin
        if (_1036)
            _6018 <= _1055;
        else
            _6018 <= _555;
    end
    assign _6023 = _1062 == _1414;
    assign _6024 = _1059 & _6023;
    assign _6028 = _6024 ? _1029 : _6027;
    assign _6030 = _1047 ? _1055 : _6028;
    assign _556 = _6030;
    always @(posedge _1038) begin
        if (_1036)
            _6027 <= _1055;
        else
            _6027 <= _556;
    end
    assign _6032 = _1062 == _1423;
    assign _6033 = _1059 & _6032;
    assign _6037 = _6033 ? _1029 : _6036;
    assign _6039 = _1047 ? _1055 : _6037;
    assign _557 = _6039;
    always @(posedge _1038) begin
        if (_1036)
            _6036 <= _1055;
        else
            _6036 <= _557;
    end
    assign _6041 = _1062 == _1432;
    assign _6042 = _1059 & _6041;
    assign _6046 = _6042 ? _1029 : _6045;
    assign _6048 = _1047 ? _1055 : _6046;
    assign _558 = _6048;
    always @(posedge _1038) begin
        if (_1036)
            _6045 <= _1055;
        else
            _6045 <= _558;
    end
    assign _6050 = _1062 == _1441;
    assign _6051 = _1059 & _6050;
    assign _6055 = _6051 ? _1029 : _6054;
    assign _6057 = _1047 ? _1055 : _6055;
    assign _559 = _6057;
    always @(posedge _1038) begin
        if (_1036)
            _6054 <= _1055;
        else
            _6054 <= _559;
    end
    assign _6059 = _1062 == _1450;
    assign _6060 = _1059 & _6059;
    assign _6064 = _6060 ? _1029 : _6063;
    assign _6066 = _1047 ? _1055 : _6064;
    assign _560 = _6066;
    always @(posedge _1038) begin
        if (_1036)
            _6063 <= _1055;
        else
            _6063 <= _560;
    end
    assign _6068 = _1062 == _1459;
    assign _6069 = _1059 & _6068;
    assign _6073 = _6069 ? _1029 : _6072;
    assign _6075 = _1047 ? _1055 : _6073;
    assign _561 = _6075;
    always @(posedge _1038) begin
        if (_1036)
            _6072 <= _1055;
        else
            _6072 <= _561;
    end
    assign _6077 = _1062 == _1468;
    assign _6078 = _1059 & _6077;
    assign _6082 = _6078 ? _1029 : _6081;
    assign _6084 = _1047 ? _1055 : _6082;
    assign _562 = _6084;
    always @(posedge _1038) begin
        if (_1036)
            _6081 <= _1055;
        else
            _6081 <= _562;
    end
    assign _6086 = _1062 == _1477;
    assign _6087 = _1059 & _6086;
    assign _6091 = _6087 ? _1029 : _6090;
    assign _6093 = _1047 ? _1055 : _6091;
    assign _563 = _6093;
    always @(posedge _1038) begin
        if (_1036)
            _6090 <= _1055;
        else
            _6090 <= _563;
    end
    assign _6095 = _1062 == _1486;
    assign _6096 = _1059 & _6095;
    assign _6100 = _6096 ? _1029 : _6099;
    assign _6102 = _1047 ? _1055 : _6100;
    assign _564 = _6102;
    always @(posedge _1038) begin
        if (_1036)
            _6099 <= _1055;
        else
            _6099 <= _564;
    end
    assign _6104 = _1062 == _1495;
    assign _6105 = _1059 & _6104;
    assign _6109 = _6105 ? _1029 : _6108;
    assign _6111 = _1047 ? _1055 : _6109;
    assign _565 = _6111;
    always @(posedge _1038) begin
        if (_1036)
            _6108 <= _1055;
        else
            _6108 <= _565;
    end
    assign _6113 = _1062 == _1504;
    assign _6114 = _1059 & _6113;
    assign _6118 = _6114 ? _1029 : _6117;
    assign _6120 = _1047 ? _1055 : _6118;
    assign _566 = _6120;
    always @(posedge _1038) begin
        if (_1036)
            _6117 <= _1055;
        else
            _6117 <= _566;
    end
    assign _6122 = _1062 == _1513;
    assign _6123 = _1059 & _6122;
    assign _6127 = _6123 ? _1029 : _6126;
    assign _6129 = _1047 ? _1055 : _6127;
    assign _567 = _6129;
    always @(posedge _1038) begin
        if (_1036)
            _6126 <= _1055;
        else
            _6126 <= _567;
    end
    assign _6131 = _1062 == _1522;
    assign _6132 = _1059 & _6131;
    assign _6136 = _6132 ? _1029 : _6135;
    assign _6138 = _1047 ? _1055 : _6136;
    assign _568 = _6138;
    always @(posedge _1038) begin
        if (_1036)
            _6135 <= _1055;
        else
            _6135 <= _568;
    end
    assign _6140 = _1062 == _1531;
    assign _6141 = _1059 & _6140;
    assign _6145 = _6141 ? _1029 : _6144;
    assign _6147 = _1047 ? _1055 : _6145;
    assign _569 = _6147;
    always @(posedge _1038) begin
        if (_1036)
            _6144 <= _1055;
        else
            _6144 <= _569;
    end
    assign _6149 = _1062 == _1540;
    assign _6150 = _1059 & _6149;
    assign _6154 = _6150 ? _1029 : _6153;
    assign _6156 = _1047 ? _1055 : _6154;
    assign _570 = _6156;
    always @(posedge _1038) begin
        if (_1036)
            _6153 <= _1055;
        else
            _6153 <= _570;
    end
    assign _6158 = _1062 == _1549;
    assign _6159 = _1059 & _6158;
    assign _6163 = _6159 ? _1029 : _6162;
    assign _6165 = _1047 ? _1055 : _6163;
    assign _571 = _6165;
    always @(posedge _1038) begin
        if (_1036)
            _6162 <= _1055;
        else
            _6162 <= _571;
    end
    assign _6167 = _1062 == _1558;
    assign _6168 = _1059 & _6167;
    assign _6172 = _6168 ? _1029 : _6171;
    assign _6174 = _1047 ? _1055 : _6172;
    assign _572 = _6174;
    always @(posedge _1038) begin
        if (_1036)
            _6171 <= _1055;
        else
            _6171 <= _572;
    end
    assign _6176 = _1062 == _1567;
    assign _6177 = _1059 & _6176;
    assign _6181 = _6177 ? _1029 : _6180;
    assign _6183 = _1047 ? _1055 : _6181;
    assign _573 = _6183;
    always @(posedge _1038) begin
        if (_1036)
            _6180 <= _1055;
        else
            _6180 <= _573;
    end
    assign _6185 = _1062 == _1576;
    assign _6186 = _1059 & _6185;
    assign _6190 = _6186 ? _1029 : _6189;
    assign _6192 = _1047 ? _1055 : _6190;
    assign _574 = _6192;
    always @(posedge _1038) begin
        if (_1036)
            _6189 <= _1055;
        else
            _6189 <= _574;
    end
    assign _6194 = _1062 == _1585;
    assign _6195 = _1059 & _6194;
    assign _6199 = _6195 ? _1029 : _6198;
    assign _6201 = _1047 ? _1055 : _6199;
    assign _575 = _6201;
    always @(posedge _1038) begin
        if (_1036)
            _6198 <= _1055;
        else
            _6198 <= _575;
    end
    assign _6203 = _1062 == _1594;
    assign _6204 = _1059 & _6203;
    assign _6208 = _6204 ? _1029 : _6207;
    assign _6210 = _1047 ? _1055 : _6208;
    assign _576 = _6210;
    always @(posedge _1038) begin
        if (_1036)
            _6207 <= _1055;
        else
            _6207 <= _576;
    end
    assign _6212 = _1062 == _1603;
    assign _6213 = _1059 & _6212;
    assign _6217 = _6213 ? _1029 : _6216;
    assign _6219 = _1047 ? _1055 : _6217;
    assign _577 = _6219;
    always @(posedge _1038) begin
        if (_1036)
            _6216 <= _1055;
        else
            _6216 <= _577;
    end
    assign _6221 = _1062 == _1612;
    assign _6222 = _1059 & _6221;
    assign _6226 = _6222 ? _1029 : _6225;
    assign _6228 = _1047 ? _1055 : _6226;
    assign _578 = _6228;
    always @(posedge _1038) begin
        if (_1036)
            _6225 <= _1055;
        else
            _6225 <= _578;
    end
    assign _6230 = _1062 == _1621;
    assign _6231 = _1059 & _6230;
    assign _6235 = _6231 ? _1029 : _6234;
    assign _6237 = _1047 ? _1055 : _6235;
    assign _579 = _6237;
    always @(posedge _1038) begin
        if (_1036)
            _6234 <= _1055;
        else
            _6234 <= _579;
    end
    assign _6239 = _1062 == _1630;
    assign _6240 = _1059 & _6239;
    assign _6244 = _6240 ? _1029 : _6243;
    assign _6246 = _1047 ? _1055 : _6244;
    assign _580 = _6246;
    always @(posedge _1038) begin
        if (_1036)
            _6243 <= _1055;
        else
            _6243 <= _580;
    end
    assign _6248 = _1062 == _1639;
    assign _6249 = _1059 & _6248;
    assign _6253 = _6249 ? _1029 : _6252;
    assign _6255 = _1047 ? _1055 : _6253;
    assign _581 = _6255;
    always @(posedge _1038) begin
        if (_1036)
            _6252 <= _1055;
        else
            _6252 <= _581;
    end
    assign _6257 = _1062 == _1648;
    assign _6258 = _1059 & _6257;
    assign _6262 = _6258 ? _1029 : _6261;
    assign _6264 = _1047 ? _1055 : _6262;
    assign _582 = _6264;
    always @(posedge _1038) begin
        if (_1036)
            _6261 <= _1055;
        else
            _6261 <= _582;
    end
    assign _6266 = _1062 == _1657;
    assign _6267 = _1059 & _6266;
    assign _6271 = _6267 ? _1029 : _6270;
    assign _6273 = _1047 ? _1055 : _6271;
    assign _583 = _6273;
    always @(posedge _1038) begin
        if (_1036)
            _6270 <= _1055;
        else
            _6270 <= _583;
    end
    assign _6275 = _1062 == _1666;
    assign _6276 = _1059 & _6275;
    assign _6280 = _6276 ? _1029 : _6279;
    assign _6282 = _1047 ? _1055 : _6280;
    assign _584 = _6282;
    always @(posedge _1038) begin
        if (_1036)
            _6279 <= _1055;
        else
            _6279 <= _584;
    end
    assign _6284 = _1062 == _1675;
    assign _6285 = _1059 & _6284;
    assign _6289 = _6285 ? _1029 : _6288;
    assign _6291 = _1047 ? _1055 : _6289;
    assign _585 = _6291;
    always @(posedge _1038) begin
        if (_1036)
            _6288 <= _1055;
        else
            _6288 <= _585;
    end
    assign _6293 = _1062 == _1684;
    assign _6294 = _1059 & _6293;
    assign _6298 = _6294 ? _1029 : _6297;
    assign _6300 = _1047 ? _1055 : _6298;
    assign _586 = _6300;
    always @(posedge _1038) begin
        if (_1036)
            _6297 <= _1055;
        else
            _6297 <= _586;
    end
    assign _6302 = _1062 == _1693;
    assign _6303 = _1059 & _6302;
    assign _6307 = _6303 ? _1029 : _6306;
    assign _6309 = _1047 ? _1055 : _6307;
    assign _587 = _6309;
    always @(posedge _1038) begin
        if (_1036)
            _6306 <= _1055;
        else
            _6306 <= _587;
    end
    assign _6311 = _1062 == _1702;
    assign _6312 = _1059 & _6311;
    assign _6316 = _6312 ? _1029 : _6315;
    assign _6318 = _1047 ? _1055 : _6316;
    assign _588 = _6318;
    always @(posedge _1038) begin
        if (_1036)
            _6315 <= _1055;
        else
            _6315 <= _588;
    end
    assign _6320 = _1062 == _1711;
    assign _6321 = _1059 & _6320;
    assign _6325 = _6321 ? _1029 : _6324;
    assign _6327 = _1047 ? _1055 : _6325;
    assign _589 = _6327;
    always @(posedge _1038) begin
        if (_1036)
            _6324 <= _1055;
        else
            _6324 <= _589;
    end
    assign _6329 = _1062 == _1720;
    assign _6330 = _1059 & _6329;
    assign _6334 = _6330 ? _1029 : _6333;
    assign _6336 = _1047 ? _1055 : _6334;
    assign _590 = _6336;
    always @(posedge _1038) begin
        if (_1036)
            _6333 <= _1055;
        else
            _6333 <= _590;
    end
    assign _6338 = _1062 == _1729;
    assign _6339 = _1059 & _6338;
    assign _6343 = _6339 ? _1029 : _6342;
    assign _6345 = _1047 ? _1055 : _6343;
    assign _591 = _6345;
    always @(posedge _1038) begin
        if (_1036)
            _6342 <= _1055;
        else
            _6342 <= _591;
    end
    assign _6347 = _1062 == _1738;
    assign _6348 = _1059 & _6347;
    assign _6352 = _6348 ? _1029 : _6351;
    assign _6354 = _1047 ? _1055 : _6352;
    assign _592 = _6354;
    always @(posedge _1038) begin
        if (_1036)
            _6351 <= _1055;
        else
            _6351 <= _592;
    end
    assign _6356 = _1062 == _1747;
    assign _6357 = _1059 & _6356;
    assign _6361 = _6357 ? _1029 : _6360;
    assign _6363 = _1047 ? _1055 : _6361;
    assign _593 = _6363;
    always @(posedge _1038) begin
        if (_1036)
            _6360 <= _1055;
        else
            _6360 <= _593;
    end
    assign _6365 = _1062 == _1756;
    assign _6366 = _1059 & _6365;
    assign _6370 = _6366 ? _1029 : _6369;
    assign _6372 = _1047 ? _1055 : _6370;
    assign _594 = _6372;
    always @(posedge _1038) begin
        if (_1036)
            _6369 <= _1055;
        else
            _6369 <= _594;
    end
    assign _6374 = _1062 == _1765;
    assign _6375 = _1059 & _6374;
    assign _6379 = _6375 ? _1029 : _6378;
    assign _6381 = _1047 ? _1055 : _6379;
    assign _595 = _6381;
    always @(posedge _1038) begin
        if (_1036)
            _6378 <= _1055;
        else
            _6378 <= _595;
    end
    assign _6383 = _1062 == _1774;
    assign _6384 = _1059 & _6383;
    assign _6388 = _6384 ? _1029 : _6387;
    assign _6390 = _1047 ? _1055 : _6388;
    assign _596 = _6390;
    always @(posedge _1038) begin
        if (_1036)
            _6387 <= _1055;
        else
            _6387 <= _596;
    end
    assign _6392 = _1062 == _1783;
    assign _6393 = _1059 & _6392;
    assign _6397 = _6393 ? _1029 : _6396;
    assign _6399 = _1047 ? _1055 : _6397;
    assign _597 = _6399;
    always @(posedge _1038) begin
        if (_1036)
            _6396 <= _1055;
        else
            _6396 <= _597;
    end
    assign _6401 = _1062 == _1792;
    assign _6402 = _1059 & _6401;
    assign _6406 = _6402 ? _1029 : _6405;
    assign _6408 = _1047 ? _1055 : _6406;
    assign _598 = _6408;
    always @(posedge _1038) begin
        if (_1036)
            _6405 <= _1055;
        else
            _6405 <= _598;
    end
    assign _6410 = _1062 == _1801;
    assign _6411 = _1059 & _6410;
    assign _6415 = _6411 ? _1029 : _6414;
    assign _6417 = _1047 ? _1055 : _6415;
    assign _599 = _6417;
    always @(posedge _1038) begin
        if (_1036)
            _6414 <= _1055;
        else
            _6414 <= _599;
    end
    assign _6419 = _1062 == _1810;
    assign _6420 = _1059 & _6419;
    assign _6424 = _6420 ? _1029 : _6423;
    assign _6426 = _1047 ? _1055 : _6424;
    assign _600 = _6426;
    always @(posedge _1038) begin
        if (_1036)
            _6423 <= _1055;
        else
            _6423 <= _600;
    end
    assign _6428 = _1062 == _1819;
    assign _6429 = _1059 & _6428;
    assign _6433 = _6429 ? _1029 : _6432;
    assign _6435 = _1047 ? _1055 : _6433;
    assign _601 = _6435;
    always @(posedge _1038) begin
        if (_1036)
            _6432 <= _1055;
        else
            _6432 <= _601;
    end
    assign _6437 = _1062 == _1828;
    assign _6438 = _1059 & _6437;
    assign _6442 = _6438 ? _1029 : _6441;
    assign _6444 = _1047 ? _1055 : _6442;
    assign _602 = _6444;
    always @(posedge _1038) begin
        if (_1036)
            _6441 <= _1055;
        else
            _6441 <= _602;
    end
    assign _6446 = _1062 == _1837;
    assign _6447 = _1059 & _6446;
    assign _6451 = _6447 ? _1029 : _6450;
    assign _6453 = _1047 ? _1055 : _6451;
    assign _603 = _6453;
    always @(posedge _1038) begin
        if (_1036)
            _6450 <= _1055;
        else
            _6450 <= _603;
    end
    assign _6455 = _1062 == _1846;
    assign _6456 = _1059 & _6455;
    assign _6460 = _6456 ? _1029 : _6459;
    assign _6462 = _1047 ? _1055 : _6460;
    assign _604 = _6462;
    always @(posedge _1038) begin
        if (_1036)
            _6459 <= _1055;
        else
            _6459 <= _604;
    end
    assign _6464 = _1062 == _1855;
    assign _6465 = _1059 & _6464;
    assign _6469 = _6465 ? _1029 : _6468;
    assign _6471 = _1047 ? _1055 : _6469;
    assign _605 = _6471;
    always @(posedge _1038) begin
        if (_1036)
            _6468 <= _1055;
        else
            _6468 <= _605;
    end
    assign _6473 = _1062 == _1864;
    assign _6474 = _1059 & _6473;
    assign _6478 = _6474 ? _1029 : _6477;
    assign _6480 = _1047 ? _1055 : _6478;
    assign _606 = _6480;
    always @(posedge _1038) begin
        if (_1036)
            _6477 <= _1055;
        else
            _6477 <= _606;
    end
    assign _6482 = _1062 == _1873;
    assign _6483 = _1059 & _6482;
    assign _6487 = _6483 ? _1029 : _6486;
    assign _6489 = _1047 ? _1055 : _6487;
    assign _607 = _6489;
    always @(posedge _1038) begin
        if (_1036)
            _6486 <= _1055;
        else
            _6486 <= _607;
    end
    assign _6491 = _1062 == _1882;
    assign _6492 = _1059 & _6491;
    assign _6496 = _6492 ? _1029 : _6495;
    assign _6498 = _1047 ? _1055 : _6496;
    assign _608 = _6498;
    always @(posedge _1038) begin
        if (_1036)
            _6495 <= _1055;
        else
            _6495 <= _608;
    end
    assign _6500 = _1062 == _1891;
    assign _6501 = _1059 & _6500;
    assign _6505 = _6501 ? _1029 : _6504;
    assign _6507 = _1047 ? _1055 : _6505;
    assign _609 = _6507;
    always @(posedge _1038) begin
        if (_1036)
            _6504 <= _1055;
        else
            _6504 <= _609;
    end
    assign _6509 = _1062 == _1900;
    assign _6510 = _1059 & _6509;
    assign _6514 = _6510 ? _1029 : _6513;
    assign _6516 = _1047 ? _1055 : _6514;
    assign _610 = _6516;
    always @(posedge _1038) begin
        if (_1036)
            _6513 <= _1055;
        else
            _6513 <= _610;
    end
    assign _6518 = _1062 == _1909;
    assign _6519 = _1059 & _6518;
    assign _6523 = _6519 ? _1029 : _6522;
    assign _6525 = _1047 ? _1055 : _6523;
    assign _611 = _6525;
    always @(posedge _1038) begin
        if (_1036)
            _6522 <= _1055;
        else
            _6522 <= _611;
    end
    assign _6527 = _1062 == _1918;
    assign _6528 = _1059 & _6527;
    assign _6532 = _6528 ? _1029 : _6531;
    assign _6534 = _1047 ? _1055 : _6532;
    assign _612 = _6534;
    always @(posedge _1038) begin
        if (_1036)
            _6531 <= _1055;
        else
            _6531 <= _612;
    end
    assign _6536 = _1062 == _1927;
    assign _6537 = _1059 & _6536;
    assign _6541 = _6537 ? _1029 : _6540;
    assign _6543 = _1047 ? _1055 : _6541;
    assign _613 = _6543;
    always @(posedge _1038) begin
        if (_1036)
            _6540 <= _1055;
        else
            _6540 <= _613;
    end
    assign _6545 = _1062 == _1936;
    assign _6546 = _1059 & _6545;
    assign _6550 = _6546 ? _1029 : _6549;
    assign _6552 = _1047 ? _1055 : _6550;
    assign _614 = _6552;
    always @(posedge _1038) begin
        if (_1036)
            _6549 <= _1055;
        else
            _6549 <= _614;
    end
    assign _6554 = _1062 == _1945;
    assign _6555 = _1059 & _6554;
    assign _6559 = _6555 ? _1029 : _6558;
    assign _6561 = _1047 ? _1055 : _6559;
    assign _615 = _6561;
    always @(posedge _1038) begin
        if (_1036)
            _6558 <= _1055;
        else
            _6558 <= _615;
    end
    assign _6563 = _1062 == _1954;
    assign _6564 = _1059 & _6563;
    assign _6568 = _6564 ? _1029 : _6567;
    assign _6570 = _1047 ? _1055 : _6568;
    assign _616 = _6570;
    always @(posedge _1038) begin
        if (_1036)
            _6567 <= _1055;
        else
            _6567 <= _616;
    end
    assign _6572 = _1062 == _1963;
    assign _6573 = _1059 & _6572;
    assign _6577 = _6573 ? _1029 : _6576;
    assign _6579 = _1047 ? _1055 : _6577;
    assign _617 = _6579;
    always @(posedge _1038) begin
        if (_1036)
            _6576 <= _1055;
        else
            _6576 <= _617;
    end
    assign _6581 = _1062 == _1972;
    assign _6582 = _1059 & _6581;
    assign _6586 = _6582 ? _1029 : _6585;
    assign _6588 = _1047 ? _1055 : _6586;
    assign _618 = _6588;
    always @(posedge _1038) begin
        if (_1036)
            _6585 <= _1055;
        else
            _6585 <= _618;
    end
    assign _6590 = _1062 == _1981;
    assign _6591 = _1059 & _6590;
    assign _6595 = _6591 ? _1029 : _6594;
    assign _6597 = _1047 ? _1055 : _6595;
    assign _619 = _6597;
    always @(posedge _1038) begin
        if (_1036)
            _6594 <= _1055;
        else
            _6594 <= _619;
    end
    assign _6599 = _1062 == _1990;
    assign _6600 = _1059 & _6599;
    assign _6604 = _6600 ? _1029 : _6603;
    assign _6606 = _1047 ? _1055 : _6604;
    assign _620 = _6606;
    always @(posedge _1038) begin
        if (_1036)
            _6603 <= _1055;
        else
            _6603 <= _620;
    end
    assign _6608 = _1062 == _1999;
    assign _6609 = _1059 & _6608;
    assign _6613 = _6609 ? _1029 : _6612;
    assign _6615 = _1047 ? _1055 : _6613;
    assign _621 = _6615;
    always @(posedge _1038) begin
        if (_1036)
            _6612 <= _1055;
        else
            _6612 <= _621;
    end
    assign _6617 = _1062 == _2008;
    assign _6618 = _1059 & _6617;
    assign _6622 = _6618 ? _1029 : _6621;
    assign _6624 = _1047 ? _1055 : _6622;
    assign _622 = _6624;
    always @(posedge _1038) begin
        if (_1036)
            _6621 <= _1055;
        else
            _6621 <= _622;
    end
    assign _6626 = _1062 == _2017;
    assign _6627 = _1059 & _6626;
    assign _6631 = _6627 ? _1029 : _6630;
    assign _6633 = _1047 ? _1055 : _6631;
    assign _623 = _6633;
    always @(posedge _1038) begin
        if (_1036)
            _6630 <= _1055;
        else
            _6630 <= _623;
    end
    assign _6635 = _1062 == _2026;
    assign _6636 = _1059 & _6635;
    assign _6640 = _6636 ? _1029 : _6639;
    assign _6642 = _1047 ? _1055 : _6640;
    assign _624 = _6642;
    always @(posedge _1038) begin
        if (_1036)
            _6639 <= _1055;
        else
            _6639 <= _624;
    end
    assign _6644 = _1062 == _2035;
    assign _6645 = _1059 & _6644;
    assign _6649 = _6645 ? _1029 : _6648;
    assign _6651 = _1047 ? _1055 : _6649;
    assign _625 = _6651;
    always @(posedge _1038) begin
        if (_1036)
            _6648 <= _1055;
        else
            _6648 <= _625;
    end
    assign _6653 = _1062 == _2044;
    assign _6654 = _1059 & _6653;
    assign _6658 = _6654 ? _1029 : _6657;
    assign _6660 = _1047 ? _1055 : _6658;
    assign _626 = _6660;
    always @(posedge _1038) begin
        if (_1036)
            _6657 <= _1055;
        else
            _6657 <= _626;
    end
    assign _6662 = _1062 == _2053;
    assign _6663 = _1059 & _6662;
    assign _6667 = _6663 ? _1029 : _6666;
    assign _6669 = _1047 ? _1055 : _6667;
    assign _627 = _6669;
    always @(posedge _1038) begin
        if (_1036)
            _6666 <= _1055;
        else
            _6666 <= _627;
    end
    assign _6671 = _1062 == _2062;
    assign _6672 = _1059 & _6671;
    assign _6676 = _6672 ? _1029 : _6675;
    assign _6678 = _1047 ? _1055 : _6676;
    assign _628 = _6678;
    always @(posedge _1038) begin
        if (_1036)
            _6675 <= _1055;
        else
            _6675 <= _628;
    end
    assign _6680 = _1062 == _2071;
    assign _6681 = _1059 & _6680;
    assign _6685 = _6681 ? _1029 : _6684;
    assign _6687 = _1047 ? _1055 : _6685;
    assign _629 = _6687;
    always @(posedge _1038) begin
        if (_1036)
            _6684 <= _1055;
        else
            _6684 <= _629;
    end
    assign _6689 = _1062 == _2080;
    assign _6690 = _1059 & _6689;
    assign _6694 = _6690 ? _1029 : _6693;
    assign _6696 = _1047 ? _1055 : _6694;
    assign _630 = _6696;
    always @(posedge _1038) begin
        if (_1036)
            _6693 <= _1055;
        else
            _6693 <= _630;
    end
    assign _6698 = _1062 == _2089;
    assign _6699 = _1059 & _6698;
    assign _6703 = _6699 ? _1029 : _6702;
    assign _6705 = _1047 ? _1055 : _6703;
    assign _631 = _6705;
    always @(posedge _1038) begin
        if (_1036)
            _6702 <= _1055;
        else
            _6702 <= _631;
    end
    assign _6707 = _1062 == _2098;
    assign _6708 = _1059 & _6707;
    assign _6712 = _6708 ? _1029 : _6711;
    assign _6714 = _1047 ? _1055 : _6712;
    assign _632 = _6714;
    always @(posedge _1038) begin
        if (_1036)
            _6711 <= _1055;
        else
            _6711 <= _632;
    end
    assign _6716 = _1062 == _2107;
    assign _6717 = _1059 & _6716;
    assign _6721 = _6717 ? _1029 : _6720;
    assign _6723 = _1047 ? _1055 : _6721;
    assign _633 = _6723;
    always @(posedge _1038) begin
        if (_1036)
            _6720 <= _1055;
        else
            _6720 <= _633;
    end
    assign _6725 = _1062 == _2116;
    assign _6726 = _1059 & _6725;
    assign _6730 = _6726 ? _1029 : _6729;
    assign _6732 = _1047 ? _1055 : _6730;
    assign _634 = _6732;
    always @(posedge _1038) begin
        if (_1036)
            _6729 <= _1055;
        else
            _6729 <= _634;
    end
    assign _6734 = _1062 == _2125;
    assign _6735 = _1059 & _6734;
    assign _6739 = _6735 ? _1029 : _6738;
    assign _6741 = _1047 ? _1055 : _6739;
    assign _635 = _6741;
    always @(posedge _1038) begin
        if (_1036)
            _6738 <= _1055;
        else
            _6738 <= _635;
    end
    assign _6743 = _1062 == _2134;
    assign _6744 = _1059 & _6743;
    assign _6748 = _6744 ? _1029 : _6747;
    assign _6750 = _1047 ? _1055 : _6748;
    assign _636 = _6750;
    always @(posedge _1038) begin
        if (_1036)
            _6747 <= _1055;
        else
            _6747 <= _636;
    end
    assign _6752 = _1062 == _2143;
    assign _6753 = _1059 & _6752;
    assign _6757 = _6753 ? _1029 : _6756;
    assign _6759 = _1047 ? _1055 : _6757;
    assign _637 = _6759;
    always @(posedge _1038) begin
        if (_1036)
            _6756 <= _1055;
        else
            _6756 <= _637;
    end
    assign _6761 = _1062 == _2152;
    assign _6762 = _1059 & _6761;
    assign _6766 = _6762 ? _1029 : _6765;
    assign _6768 = _1047 ? _1055 : _6766;
    assign _638 = _6768;
    always @(posedge _1038) begin
        if (_1036)
            _6765 <= _1055;
        else
            _6765 <= _638;
    end
    assign _6770 = _1062 == _2161;
    assign _6771 = _1059 & _6770;
    assign _6775 = _6771 ? _1029 : _6774;
    assign _6777 = _1047 ? _1055 : _6775;
    assign _639 = _6777;
    always @(posedge _1038) begin
        if (_1036)
            _6774 <= _1055;
        else
            _6774 <= _639;
    end
    assign _6779 = _1062 == _2170;
    assign _6780 = _1059 & _6779;
    assign _6784 = _6780 ? _1029 : _6783;
    assign _6786 = _1047 ? _1055 : _6784;
    assign _640 = _6786;
    always @(posedge _1038) begin
        if (_1036)
            _6783 <= _1055;
        else
            _6783 <= _640;
    end
    assign _6788 = _1062 == _2179;
    assign _6789 = _1059 & _6788;
    assign _6793 = _6789 ? _1029 : _6792;
    assign _6795 = _1047 ? _1055 : _6793;
    assign _641 = _6795;
    always @(posedge _1038) begin
        if (_1036)
            _6792 <= _1055;
        else
            _6792 <= _641;
    end
    assign _6797 = _1062 == _2188;
    assign _6798 = _1059 & _6797;
    assign _6802 = _6798 ? _1029 : _6801;
    assign _6804 = _1047 ? _1055 : _6802;
    assign _642 = _6804;
    always @(posedge _1038) begin
        if (_1036)
            _6801 <= _1055;
        else
            _6801 <= _642;
    end
    assign _6806 = _1062 == _2197;
    assign _6807 = _1059 & _6806;
    assign _6811 = _6807 ? _1029 : _6810;
    assign _6813 = _1047 ? _1055 : _6811;
    assign _643 = _6813;
    always @(posedge _1038) begin
        if (_1036)
            _6810 <= _1055;
        else
            _6810 <= _643;
    end
    assign _6815 = _1062 == _2206;
    assign _6816 = _1059 & _6815;
    assign _6820 = _6816 ? _1029 : _6819;
    assign _6822 = _1047 ? _1055 : _6820;
    assign _644 = _6822;
    always @(posedge _1038) begin
        if (_1036)
            _6819 <= _1055;
        else
            _6819 <= _644;
    end
    assign _6824 = _1062 == _2215;
    assign _6825 = _1059 & _6824;
    assign _6829 = _6825 ? _1029 : _6828;
    assign _6831 = _1047 ? _1055 : _6829;
    assign _645 = _6831;
    always @(posedge _1038) begin
        if (_1036)
            _6828 <= _1055;
        else
            _6828 <= _645;
    end
    assign _6833 = _1062 == _2224;
    assign _6834 = _1059 & _6833;
    assign _6838 = _6834 ? _1029 : _6837;
    assign _6840 = _1047 ? _1055 : _6838;
    assign _646 = _6840;
    always @(posedge _1038) begin
        if (_1036)
            _6837 <= _1055;
        else
            _6837 <= _646;
    end
    assign _6842 = _1062 == _2233;
    assign _6843 = _1059 & _6842;
    assign _6847 = _6843 ? _1029 : _6846;
    assign _6849 = _1047 ? _1055 : _6847;
    assign _647 = _6849;
    always @(posedge _1038) begin
        if (_1036)
            _6846 <= _1055;
        else
            _6846 <= _647;
    end
    assign _6851 = _1062 == _2242;
    assign _6852 = _1059 & _6851;
    assign _6856 = _6852 ? _1029 : _6855;
    assign _6858 = _1047 ? _1055 : _6856;
    assign _648 = _6858;
    always @(posedge _1038) begin
        if (_1036)
            _6855 <= _1055;
        else
            _6855 <= _648;
    end
    assign _6860 = _1062 == _2251;
    assign _6861 = _1059 & _6860;
    assign _6865 = _6861 ? _1029 : _6864;
    assign _6867 = _1047 ? _1055 : _6865;
    assign _649 = _6867;
    always @(posedge _1038) begin
        if (_1036)
            _6864 <= _1055;
        else
            _6864 <= _649;
    end
    assign _6869 = _1062 == _2260;
    assign _6870 = _1059 & _6869;
    assign _6874 = _6870 ? _1029 : _6873;
    assign _6876 = _1047 ? _1055 : _6874;
    assign _650 = _6876;
    always @(posedge _1038) begin
        if (_1036)
            _6873 <= _1055;
        else
            _6873 <= _650;
    end
    assign _6878 = _1062 == _2269;
    assign _6879 = _1059 & _6878;
    assign _6883 = _6879 ? _1029 : _6882;
    assign _6885 = _1047 ? _1055 : _6883;
    assign _651 = _6885;
    always @(posedge _1038) begin
        if (_1036)
            _6882 <= _1055;
        else
            _6882 <= _651;
    end
    assign _6887 = _1062 == _2278;
    assign _6888 = _1059 & _6887;
    assign _6892 = _6888 ? _1029 : _6891;
    assign _6894 = _1047 ? _1055 : _6892;
    assign _652 = _6894;
    always @(posedge _1038) begin
        if (_1036)
            _6891 <= _1055;
        else
            _6891 <= _652;
    end
    assign _6896 = _1062 == _2287;
    assign _6897 = _1059 & _6896;
    assign _6901 = _6897 ? _1029 : _6900;
    assign _6903 = _1047 ? _1055 : _6901;
    assign _653 = _6903;
    always @(posedge _1038) begin
        if (_1036)
            _6900 <= _1055;
        else
            _6900 <= _653;
    end
    assign _6905 = _1062 == _2296;
    assign _6906 = _1059 & _6905;
    assign _6910 = _6906 ? _1029 : _6909;
    assign _6912 = _1047 ? _1055 : _6910;
    assign _654 = _6912;
    always @(posedge _1038) begin
        if (_1036)
            _6909 <= _1055;
        else
            _6909 <= _654;
    end
    assign _6914 = _1062 == _2305;
    assign _6915 = _1059 & _6914;
    assign _6919 = _6915 ? _1029 : _6918;
    assign _6921 = _1047 ? _1055 : _6919;
    assign _655 = _6921;
    always @(posedge _1038) begin
        if (_1036)
            _6918 <= _1055;
        else
            _6918 <= _655;
    end
    assign _6923 = _1062 == _2314;
    assign _6924 = _1059 & _6923;
    assign _6928 = _6924 ? _1029 : _6927;
    assign _6930 = _1047 ? _1055 : _6928;
    assign _656 = _6930;
    always @(posedge _1038) begin
        if (_1036)
            _6927 <= _1055;
        else
            _6927 <= _656;
    end
    assign _6932 = _1062 == _2323;
    assign _6933 = _1059 & _6932;
    assign _6937 = _6933 ? _1029 : _6936;
    assign _6939 = _1047 ? _1055 : _6937;
    assign _657 = _6939;
    always @(posedge _1038) begin
        if (_1036)
            _6936 <= _1055;
        else
            _6936 <= _657;
    end
    assign _6941 = _1062 == _2332;
    assign _6942 = _1059 & _6941;
    assign _6946 = _6942 ? _1029 : _6945;
    assign _6948 = _1047 ? _1055 : _6946;
    assign _658 = _6948;
    always @(posedge _1038) begin
        if (_1036)
            _6945 <= _1055;
        else
            _6945 <= _658;
    end
    assign _6950 = _1062 == _2341;
    assign _6951 = _1059 & _6950;
    assign _6955 = _6951 ? _1029 : _6954;
    assign _6957 = _1047 ? _1055 : _6955;
    assign _659 = _6957;
    always @(posedge _1038) begin
        if (_1036)
            _6954 <= _1055;
        else
            _6954 <= _659;
    end
    assign _6959 = _1062 == _2350;
    assign _6960 = _1059 & _6959;
    assign _6964 = _6960 ? _1029 : _6963;
    assign _6966 = _1047 ? _1055 : _6964;
    assign _660 = _6966;
    always @(posedge _1038) begin
        if (_1036)
            _6963 <= _1055;
        else
            _6963 <= _660;
    end
    assign _6968 = _1062 == _2359;
    assign _6969 = _1059 & _6968;
    assign _6973 = _6969 ? _1029 : _6972;
    assign _6975 = _1047 ? _1055 : _6973;
    assign _661 = _6975;
    always @(posedge _1038) begin
        if (_1036)
            _6972 <= _1055;
        else
            _6972 <= _661;
    end
    assign _6977 = _1062 == _2368;
    assign _6978 = _1059 & _6977;
    assign _6982 = _6978 ? _1029 : _6981;
    assign _6984 = _1047 ? _1055 : _6982;
    assign _662 = _6984;
    always @(posedge _1038) begin
        if (_1036)
            _6981 <= _1055;
        else
            _6981 <= _662;
    end
    assign _6986 = _1062 == _2377;
    assign _6987 = _1059 & _6986;
    assign _6991 = _6987 ? _1029 : _6990;
    assign _6993 = _1047 ? _1055 : _6991;
    assign _663 = _6993;
    always @(posedge _1038) begin
        if (_1036)
            _6990 <= _1055;
        else
            _6990 <= _663;
    end
    assign _6995 = _1062 == _2386;
    assign _6996 = _1059 & _6995;
    assign _7000 = _6996 ? _1029 : _6999;
    assign _7002 = _1047 ? _1055 : _7000;
    assign _664 = _7002;
    always @(posedge _1038) begin
        if (_1036)
            _6999 <= _1055;
        else
            _6999 <= _664;
    end
    assign _7004 = _1062 == _2395;
    assign _7005 = _1059 & _7004;
    assign _7009 = _7005 ? _1029 : _7008;
    assign _7011 = _1047 ? _1055 : _7009;
    assign _665 = _7011;
    always @(posedge _1038) begin
        if (_1036)
            _7008 <= _1055;
        else
            _7008 <= _665;
    end
    assign _7013 = _1062 == _2404;
    assign _7014 = _1059 & _7013;
    assign _7018 = _7014 ? _1029 : _7017;
    assign _7020 = _1047 ? _1055 : _7018;
    assign _666 = _7020;
    always @(posedge _1038) begin
        if (_1036)
            _7017 <= _1055;
        else
            _7017 <= _666;
    end
    assign _7022 = _1062 == _2413;
    assign _7023 = _1059 & _7022;
    assign _7027 = _7023 ? _1029 : _7026;
    assign _7029 = _1047 ? _1055 : _7027;
    assign _667 = _7029;
    always @(posedge _1038) begin
        if (_1036)
            _7026 <= _1055;
        else
            _7026 <= _667;
    end
    assign _7031 = _1062 == _2422;
    assign _7032 = _1059 & _7031;
    assign _7036 = _7032 ? _1029 : _7035;
    assign _7038 = _1047 ? _1055 : _7036;
    assign _668 = _7038;
    always @(posedge _1038) begin
        if (_1036)
            _7035 <= _1055;
        else
            _7035 <= _668;
    end
    assign _7040 = _1062 == _2431;
    assign _7041 = _1059 & _7040;
    assign _7045 = _7041 ? _1029 : _7044;
    assign _7047 = _1047 ? _1055 : _7045;
    assign _669 = _7047;
    always @(posedge _1038) begin
        if (_1036)
            _7044 <= _1055;
        else
            _7044 <= _669;
    end
    assign _7049 = _1062 == _2440;
    assign _7050 = _1059 & _7049;
    assign _7054 = _7050 ? _1029 : _7053;
    assign _7056 = _1047 ? _1055 : _7054;
    assign _670 = _7056;
    always @(posedge _1038) begin
        if (_1036)
            _7053 <= _1055;
        else
            _7053 <= _670;
    end
    assign _7058 = _1062 == _2449;
    assign _7059 = _1059 & _7058;
    assign _7063 = _7059 ? _1029 : _7062;
    assign _7065 = _1047 ? _1055 : _7063;
    assign _671 = _7065;
    always @(posedge _1038) begin
        if (_1036)
            _7062 <= _1055;
        else
            _7062 <= _671;
    end
    assign _7067 = _1062 == _2458;
    assign _7068 = _1059 & _7067;
    assign _7072 = _7068 ? _1029 : _7071;
    assign _7074 = _1047 ? _1055 : _7072;
    assign _672 = _7074;
    always @(posedge _1038) begin
        if (_1036)
            _7071 <= _1055;
        else
            _7071 <= _672;
    end
    assign _7076 = _1062 == _2467;
    assign _7077 = _1059 & _7076;
    assign _7081 = _7077 ? _1029 : _7080;
    assign _7083 = _1047 ? _1055 : _7081;
    assign _673 = _7083;
    always @(posedge _1038) begin
        if (_1036)
            _7080 <= _1055;
        else
            _7080 <= _673;
    end
    assign _7085 = _1062 == _2476;
    assign _7086 = _1059 & _7085;
    assign _7090 = _7086 ? _1029 : _7089;
    assign _7092 = _1047 ? _1055 : _7090;
    assign _674 = _7092;
    always @(posedge _1038) begin
        if (_1036)
            _7089 <= _1055;
        else
            _7089 <= _674;
    end
    assign _7094 = _1062 == _2485;
    assign _7095 = _1059 & _7094;
    assign _7099 = _7095 ? _1029 : _7098;
    assign _7101 = _1047 ? _1055 : _7099;
    assign _675 = _7101;
    always @(posedge _1038) begin
        if (_1036)
            _7098 <= _1055;
        else
            _7098 <= _675;
    end
    assign _7103 = _1062 == _2494;
    assign _7104 = _1059 & _7103;
    assign _7108 = _7104 ? _1029 : _7107;
    assign _7110 = _1047 ? _1055 : _7108;
    assign _676 = _7110;
    always @(posedge _1038) begin
        if (_1036)
            _7107 <= _1055;
        else
            _7107 <= _676;
    end
    assign _7112 = _1062 == _2503;
    assign _7113 = _1059 & _7112;
    assign _7117 = _7113 ? _1029 : _7116;
    assign _7119 = _1047 ? _1055 : _7117;
    assign _677 = _7119;
    always @(posedge _1038) begin
        if (_1036)
            _7116 <= _1055;
        else
            _7116 <= _677;
    end
    assign _7121 = _1062 == _2512;
    assign _7122 = _1059 & _7121;
    assign _7126 = _7122 ? _1029 : _7125;
    assign _7128 = _1047 ? _1055 : _7126;
    assign _678 = _7128;
    always @(posedge _1038) begin
        if (_1036)
            _7125 <= _1055;
        else
            _7125 <= _678;
    end
    assign _7130 = _1062 == _2521;
    assign _7131 = _1059 & _7130;
    assign _7135 = _7131 ? _1029 : _7134;
    assign _7137 = _1047 ? _1055 : _7135;
    assign _679 = _7137;
    always @(posedge _1038) begin
        if (_1036)
            _7134 <= _1055;
        else
            _7134 <= _679;
    end
    assign _7139 = _1062 == _2530;
    assign _7140 = _1059 & _7139;
    assign _7144 = _7140 ? _1029 : _7143;
    assign _7146 = _1047 ? _1055 : _7144;
    assign _680 = _7146;
    always @(posedge _1038) begin
        if (_1036)
            _7143 <= _1055;
        else
            _7143 <= _680;
    end
    assign _7148 = _1062 == _2539;
    assign _7149 = _1059 & _7148;
    assign _7153 = _7149 ? _1029 : _7152;
    assign _7155 = _1047 ? _1055 : _7153;
    assign _681 = _7155;
    always @(posedge _1038) begin
        if (_1036)
            _7152 <= _1055;
        else
            _7152 <= _681;
    end
    assign _7157 = _1062 == _2548;
    assign _7158 = _1059 & _7157;
    assign _7162 = _7158 ? _1029 : _7161;
    assign _7164 = _1047 ? _1055 : _7162;
    assign _682 = _7164;
    always @(posedge _1038) begin
        if (_1036)
            _7161 <= _1055;
        else
            _7161 <= _682;
    end
    assign _7166 = _1062 == _2557;
    assign _7167 = _1059 & _7166;
    assign _7171 = _7167 ? _1029 : _7170;
    assign _7173 = _1047 ? _1055 : _7171;
    assign _683 = _7173;
    always @(posedge _1038) begin
        if (_1036)
            _7170 <= _1055;
        else
            _7170 <= _683;
    end
    assign _7175 = _1062 == _2566;
    assign _7176 = _1059 & _7175;
    assign _7180 = _7176 ? _1029 : _7179;
    assign _7182 = _1047 ? _1055 : _7180;
    assign _684 = _7182;
    always @(posedge _1038) begin
        if (_1036)
            _7179 <= _1055;
        else
            _7179 <= _684;
    end
    assign _7184 = _1062 == _2575;
    assign _7185 = _1059 & _7184;
    assign _7189 = _7185 ? _1029 : _7188;
    assign _7191 = _1047 ? _1055 : _7189;
    assign _685 = _7191;
    always @(posedge _1038) begin
        if (_1036)
            _7188 <= _1055;
        else
            _7188 <= _685;
    end
    assign _7193 = _1062 == _2584;
    assign _7194 = _1059 & _7193;
    assign _7198 = _7194 ? _1029 : _7197;
    assign _7200 = _1047 ? _1055 : _7198;
    assign _686 = _7200;
    always @(posedge _1038) begin
        if (_1036)
            _7197 <= _1055;
        else
            _7197 <= _686;
    end
    assign _7202 = _1062 == _2593;
    assign _7203 = _1059 & _7202;
    assign _7207 = _7203 ? _1029 : _7206;
    assign _7209 = _1047 ? _1055 : _7207;
    assign _687 = _7209;
    always @(posedge _1038) begin
        if (_1036)
            _7206 <= _1055;
        else
            _7206 <= _687;
    end
    assign _7211 = _1062 == _2602;
    assign _7212 = _1059 & _7211;
    assign _7216 = _7212 ? _1029 : _7215;
    assign _7218 = _1047 ? _1055 : _7216;
    assign _688 = _7218;
    always @(posedge _1038) begin
        if (_1036)
            _7215 <= _1055;
        else
            _7215 <= _688;
    end
    assign _7220 = _1062 == _2611;
    assign _7221 = _1059 & _7220;
    assign _7225 = _7221 ? _1029 : _7224;
    assign _7227 = _1047 ? _1055 : _7225;
    assign _689 = _7227;
    always @(posedge _1038) begin
        if (_1036)
            _7224 <= _1055;
        else
            _7224 <= _689;
    end
    assign _7229 = _1062 == _2620;
    assign _7230 = _1059 & _7229;
    assign _7234 = _7230 ? _1029 : _7233;
    assign _7236 = _1047 ? _1055 : _7234;
    assign _690 = _7236;
    always @(posedge _1038) begin
        if (_1036)
            _7233 <= _1055;
        else
            _7233 <= _690;
    end
    assign _7238 = _1062 == _2629;
    assign _7239 = _1059 & _7238;
    assign _7243 = _7239 ? _1029 : _7242;
    assign _7245 = _1047 ? _1055 : _7243;
    assign _691 = _7245;
    always @(posedge _1038) begin
        if (_1036)
            _7242 <= _1055;
        else
            _7242 <= _691;
    end
    assign _7247 = _1062 == _2638;
    assign _7248 = _1059 & _7247;
    assign _7252 = _7248 ? _1029 : _7251;
    assign _7254 = _1047 ? _1055 : _7252;
    assign _692 = _7254;
    always @(posedge _1038) begin
        if (_1036)
            _7251 <= _1055;
        else
            _7251 <= _692;
    end
    assign _7256 = _1062 == _2647;
    assign _7257 = _1059 & _7256;
    assign _7261 = _7257 ? _1029 : _7260;
    assign _7263 = _1047 ? _1055 : _7261;
    assign _693 = _7263;
    always @(posedge _1038) begin
        if (_1036)
            _7260 <= _1055;
        else
            _7260 <= _693;
    end
    assign _7265 = _1062 == _2656;
    assign _7266 = _1059 & _7265;
    assign _7270 = _7266 ? _1029 : _7269;
    assign _7272 = _1047 ? _1055 : _7270;
    assign _694 = _7272;
    always @(posedge _1038) begin
        if (_1036)
            _7269 <= _1055;
        else
            _7269 <= _694;
    end
    assign _7274 = _1062 == _2665;
    assign _7275 = _1059 & _7274;
    assign _7279 = _7275 ? _1029 : _7278;
    assign _7281 = _1047 ? _1055 : _7279;
    assign _695 = _7281;
    always @(posedge _1038) begin
        if (_1036)
            _7278 <= _1055;
        else
            _7278 <= _695;
    end
    assign _7283 = _1062 == _2674;
    assign _7284 = _1059 & _7283;
    assign _7288 = _7284 ? _1029 : _7287;
    assign _7290 = _1047 ? _1055 : _7288;
    assign _696 = _7290;
    always @(posedge _1038) begin
        if (_1036)
            _7287 <= _1055;
        else
            _7287 <= _696;
    end
    assign _7292 = _1062 == _2683;
    assign _7293 = _1059 & _7292;
    assign _7297 = _7293 ? _1029 : _7296;
    assign _7299 = _1047 ? _1055 : _7297;
    assign _697 = _7299;
    always @(posedge _1038) begin
        if (_1036)
            _7296 <= _1055;
        else
            _7296 <= _697;
    end
    assign _7301 = _1062 == _2692;
    assign _7302 = _1059 & _7301;
    assign _7306 = _7302 ? _1029 : _7305;
    assign _7308 = _1047 ? _1055 : _7306;
    assign _698 = _7308;
    always @(posedge _1038) begin
        if (_1036)
            _7305 <= _1055;
        else
            _7305 <= _698;
    end
    assign _7310 = _1062 == _2701;
    assign _7311 = _1059 & _7310;
    assign _7315 = _7311 ? _1029 : _7314;
    assign _7317 = _1047 ? _1055 : _7315;
    assign _699 = _7317;
    always @(posedge _1038) begin
        if (_1036)
            _7314 <= _1055;
        else
            _7314 <= _699;
    end
    assign _7319 = _1062 == _2710;
    assign _7320 = _1059 & _7319;
    assign _7324 = _7320 ? _1029 : _7323;
    assign _7326 = _1047 ? _1055 : _7324;
    assign _700 = _7326;
    always @(posedge _1038) begin
        if (_1036)
            _7323 <= _1055;
        else
            _7323 <= _700;
    end
    assign _7328 = _1062 == _2719;
    assign _7329 = _1059 & _7328;
    assign _7333 = _7329 ? _1029 : _7332;
    assign _7335 = _1047 ? _1055 : _7333;
    assign _701 = _7335;
    always @(posedge _1038) begin
        if (_1036)
            _7332 <= _1055;
        else
            _7332 <= _701;
    end
    assign _7337 = _1062 == _2728;
    assign _7338 = _1059 & _7337;
    assign _7342 = _7338 ? _1029 : _7341;
    assign _7344 = _1047 ? _1055 : _7342;
    assign _702 = _7344;
    always @(posedge _1038) begin
        if (_1036)
            _7341 <= _1055;
        else
            _7341 <= _702;
    end
    assign _7346 = _1062 == _2737;
    assign _7347 = _1059 & _7346;
    assign _7351 = _7347 ? _1029 : _7350;
    assign _7353 = _1047 ? _1055 : _7351;
    assign _703 = _7353;
    always @(posedge _1038) begin
        if (_1036)
            _7350 <= _1055;
        else
            _7350 <= _703;
    end
    assign _7355 = _1062 == _2746;
    assign _7356 = _1059 & _7355;
    assign _7360 = _7356 ? _1029 : _7359;
    assign _7362 = _1047 ? _1055 : _7360;
    assign _704 = _7362;
    always @(posedge _1038) begin
        if (_1036)
            _7359 <= _1055;
        else
            _7359 <= _704;
    end
    assign _7364 = _1062 == _2755;
    assign _7365 = _1059 & _7364;
    assign _7369 = _7365 ? _1029 : _7368;
    assign _7371 = _1047 ? _1055 : _7369;
    assign _705 = _7371;
    always @(posedge _1038) begin
        if (_1036)
            _7368 <= _1055;
        else
            _7368 <= _705;
    end
    assign _7373 = _1062 == _2764;
    assign _7374 = _1059 & _7373;
    assign _7378 = _7374 ? _1029 : _7377;
    assign _7380 = _1047 ? _1055 : _7378;
    assign _706 = _7380;
    always @(posedge _1038) begin
        if (_1036)
            _7377 <= _1055;
        else
            _7377 <= _706;
    end
    assign _7382 = _1062 == _2773;
    assign _7383 = _1059 & _7382;
    assign _7387 = _7383 ? _1029 : _7386;
    assign _7389 = _1047 ? _1055 : _7387;
    assign _707 = _7389;
    always @(posedge _1038) begin
        if (_1036)
            _7386 <= _1055;
        else
            _7386 <= _707;
    end
    assign _7391 = _1062 == _2782;
    assign _7392 = _1059 & _7391;
    assign _7396 = _7392 ? _1029 : _7395;
    assign _7398 = _1047 ? _1055 : _7396;
    assign _708 = _7398;
    always @(posedge _1038) begin
        if (_1036)
            _7395 <= _1055;
        else
            _7395 <= _708;
    end
    assign _7400 = _1062 == _2791;
    assign _7401 = _1059 & _7400;
    assign _7405 = _7401 ? _1029 : _7404;
    assign _7407 = _1047 ? _1055 : _7405;
    assign _709 = _7407;
    always @(posedge _1038) begin
        if (_1036)
            _7404 <= _1055;
        else
            _7404 <= _709;
    end
    assign _7409 = _1062 == _2800;
    assign _7410 = _1059 & _7409;
    assign _7414 = _7410 ? _1029 : _7413;
    assign _7416 = _1047 ? _1055 : _7414;
    assign _710 = _7416;
    always @(posedge _1038) begin
        if (_1036)
            _7413 <= _1055;
        else
            _7413 <= _710;
    end
    assign _7418 = _1062 == _2809;
    assign _7419 = _1059 & _7418;
    assign _7423 = _7419 ? _1029 : _7422;
    assign _7425 = _1047 ? _1055 : _7423;
    assign _711 = _7425;
    always @(posedge _1038) begin
        if (_1036)
            _7422 <= _1055;
        else
            _7422 <= _711;
    end
    assign _7427 = _1062 == _2818;
    assign _7428 = _1059 & _7427;
    assign _7432 = _7428 ? _1029 : _7431;
    assign _7434 = _1047 ? _1055 : _7432;
    assign _712 = _7434;
    always @(posedge _1038) begin
        if (_1036)
            _7431 <= _1055;
        else
            _7431 <= _712;
    end
    assign _7436 = _1062 == _2827;
    assign _7437 = _1059 & _7436;
    assign _7441 = _7437 ? _1029 : _7440;
    assign _7443 = _1047 ? _1055 : _7441;
    assign _713 = _7443;
    always @(posedge _1038) begin
        if (_1036)
            _7440 <= _1055;
        else
            _7440 <= _713;
    end
    assign _7445 = _1062 == _2836;
    assign _7446 = _1059 & _7445;
    assign _7450 = _7446 ? _1029 : _7449;
    assign _7452 = _1047 ? _1055 : _7450;
    assign _714 = _7452;
    always @(posedge _1038) begin
        if (_1036)
            _7449 <= _1055;
        else
            _7449 <= _714;
    end
    assign _7454 = _1062 == _2845;
    assign _7455 = _1059 & _7454;
    assign _7459 = _7455 ? _1029 : _7458;
    assign _7461 = _1047 ? _1055 : _7459;
    assign _715 = _7461;
    always @(posedge _1038) begin
        if (_1036)
            _7458 <= _1055;
        else
            _7458 <= _715;
    end
    assign _7463 = _1062 == _2854;
    assign _7464 = _1059 & _7463;
    assign _7468 = _7464 ? _1029 : _7467;
    assign _7470 = _1047 ? _1055 : _7468;
    assign _716 = _7470;
    always @(posedge _1038) begin
        if (_1036)
            _7467 <= _1055;
        else
            _7467 <= _716;
    end
    assign _7472 = _1062 == _2863;
    assign _7473 = _1059 & _7472;
    assign _7477 = _7473 ? _1029 : _7476;
    assign _7479 = _1047 ? _1055 : _7477;
    assign _717 = _7479;
    always @(posedge _1038) begin
        if (_1036)
            _7476 <= _1055;
        else
            _7476 <= _717;
    end
    assign _7481 = _1062 == _2872;
    assign _7482 = _1059 & _7481;
    assign _7486 = _7482 ? _1029 : _7485;
    assign _7488 = _1047 ? _1055 : _7486;
    assign _718 = _7488;
    always @(posedge _1038) begin
        if (_1036)
            _7485 <= _1055;
        else
            _7485 <= _718;
    end
    assign _7490 = _1062 == _2881;
    assign _7491 = _1059 & _7490;
    assign _7495 = _7491 ? _1029 : _7494;
    assign _7497 = _1047 ? _1055 : _7495;
    assign _719 = _7497;
    always @(posedge _1038) begin
        if (_1036)
            _7494 <= _1055;
        else
            _7494 <= _719;
    end
    assign _7499 = _1062 == _2890;
    assign _7500 = _1059 & _7499;
    assign _7504 = _7500 ? _1029 : _7503;
    assign _7506 = _1047 ? _1055 : _7504;
    assign _720 = _7506;
    always @(posedge _1038) begin
        if (_1036)
            _7503 <= _1055;
        else
            _7503 <= _720;
    end
    assign _7508 = _1062 == _2899;
    assign _7509 = _1059 & _7508;
    assign _7513 = _7509 ? _1029 : _7512;
    assign _7515 = _1047 ? _1055 : _7513;
    assign _721 = _7515;
    always @(posedge _1038) begin
        if (_1036)
            _7512 <= _1055;
        else
            _7512 <= _721;
    end
    assign _7517 = _1062 == _2908;
    assign _7518 = _1059 & _7517;
    assign _7522 = _7518 ? _1029 : _7521;
    assign _7524 = _1047 ? _1055 : _7522;
    assign _722 = _7524;
    always @(posedge _1038) begin
        if (_1036)
            _7521 <= _1055;
        else
            _7521 <= _722;
    end
    assign _7526 = _1062 == _2917;
    assign _7527 = _1059 & _7526;
    assign _7531 = _7527 ? _1029 : _7530;
    assign _7533 = _1047 ? _1055 : _7531;
    assign _723 = _7533;
    always @(posedge _1038) begin
        if (_1036)
            _7530 <= _1055;
        else
            _7530 <= _723;
    end
    assign _7535 = _1062 == _2926;
    assign _7536 = _1059 & _7535;
    assign _7540 = _7536 ? _1029 : _7539;
    assign _7542 = _1047 ? _1055 : _7540;
    assign _724 = _7542;
    always @(posedge _1038) begin
        if (_1036)
            _7539 <= _1055;
        else
            _7539 <= _724;
    end
    assign _7544 = _1062 == _2935;
    assign _7545 = _1059 & _7544;
    assign _7549 = _7545 ? _1029 : _7548;
    assign _7551 = _1047 ? _1055 : _7549;
    assign _725 = _7551;
    always @(posedge _1038) begin
        if (_1036)
            _7548 <= _1055;
        else
            _7548 <= _725;
    end
    assign _7553 = _1062 == _2944;
    assign _7554 = _1059 & _7553;
    assign _7558 = _7554 ? _1029 : _7557;
    assign _7560 = _1047 ? _1055 : _7558;
    assign _726 = _7560;
    always @(posedge _1038) begin
        if (_1036)
            _7557 <= _1055;
        else
            _7557 <= _726;
    end
    assign _7562 = _1062 == _2953;
    assign _7563 = _1059 & _7562;
    assign _7567 = _7563 ? _1029 : _7566;
    assign _7569 = _1047 ? _1055 : _7567;
    assign _727 = _7569;
    always @(posedge _1038) begin
        if (_1036)
            _7566 <= _1055;
        else
            _7566 <= _727;
    end
    assign _7571 = _1062 == _2962;
    assign _7572 = _1059 & _7571;
    assign _7576 = _7572 ? _1029 : _7575;
    assign _7578 = _1047 ? _1055 : _7576;
    assign _728 = _7578;
    always @(posedge _1038) begin
        if (_1036)
            _7575 <= _1055;
        else
            _7575 <= _728;
    end
    assign _7580 = _1062 == _2971;
    assign _7581 = _1059 & _7580;
    assign _7585 = _7581 ? _1029 : _7584;
    assign _7587 = _1047 ? _1055 : _7585;
    assign _729 = _7587;
    always @(posedge _1038) begin
        if (_1036)
            _7584 <= _1055;
        else
            _7584 <= _729;
    end
    assign _7589 = _1062 == _2980;
    assign _7590 = _1059 & _7589;
    assign _7594 = _7590 ? _1029 : _7593;
    assign _7596 = _1047 ? _1055 : _7594;
    assign _730 = _7596;
    always @(posedge _1038) begin
        if (_1036)
            _7593 <= _1055;
        else
            _7593 <= _730;
    end
    assign _7598 = _1062 == _2989;
    assign _7599 = _1059 & _7598;
    assign _7603 = _7599 ? _1029 : _7602;
    assign _7605 = _1047 ? _1055 : _7603;
    assign _731 = _7605;
    always @(posedge _1038) begin
        if (_1036)
            _7602 <= _1055;
        else
            _7602 <= _731;
    end
    assign _7607 = _1062 == _2998;
    assign _7608 = _1059 & _7607;
    assign _7612 = _7608 ? _1029 : _7611;
    assign _7614 = _1047 ? _1055 : _7612;
    assign _732 = _7614;
    always @(posedge _1038) begin
        if (_1036)
            _7611 <= _1055;
        else
            _7611 <= _732;
    end
    assign _7616 = _1062 == _3007;
    assign _7617 = _1059 & _7616;
    assign _7621 = _7617 ? _1029 : _7620;
    assign _7623 = _1047 ? _1055 : _7621;
    assign _733 = _7623;
    always @(posedge _1038) begin
        if (_1036)
            _7620 <= _1055;
        else
            _7620 <= _733;
    end
    assign _7625 = _1062 == _3016;
    assign _7626 = _1059 & _7625;
    assign _7630 = _7626 ? _1029 : _7629;
    assign _7632 = _1047 ? _1055 : _7630;
    assign _734 = _7632;
    always @(posedge _1038) begin
        if (_1036)
            _7629 <= _1055;
        else
            _7629 <= _734;
    end
    assign _7634 = _1062 == _3025;
    assign _7635 = _1059 & _7634;
    assign _7639 = _7635 ? _1029 : _7638;
    assign _7641 = _1047 ? _1055 : _7639;
    assign _735 = _7641;
    always @(posedge _1038) begin
        if (_1036)
            _7638 <= _1055;
        else
            _7638 <= _735;
    end
    assign _7643 = _1062 == _3034;
    assign _7644 = _1059 & _7643;
    assign _7648 = _7644 ? _1029 : _7647;
    assign _7650 = _1047 ? _1055 : _7648;
    assign _736 = _7650;
    always @(posedge _1038) begin
        if (_1036)
            _7647 <= _1055;
        else
            _7647 <= _736;
    end
    assign _7652 = _1062 == _3043;
    assign _7653 = _1059 & _7652;
    assign _7657 = _7653 ? _1029 : _7656;
    assign _7659 = _1047 ? _1055 : _7657;
    assign _737 = _7659;
    always @(posedge _1038) begin
        if (_1036)
            _7656 <= _1055;
        else
            _7656 <= _737;
    end
    assign _7661 = _1062 == _3052;
    assign _7662 = _1059 & _7661;
    assign _7666 = _7662 ? _1029 : _7665;
    assign _7668 = _1047 ? _1055 : _7666;
    assign _738 = _7668;
    always @(posedge _1038) begin
        if (_1036)
            _7665 <= _1055;
        else
            _7665 <= _738;
    end
    assign _7670 = _1062 == _3061;
    assign _7671 = _1059 & _7670;
    assign _7675 = _7671 ? _1029 : _7674;
    assign _7677 = _1047 ? _1055 : _7675;
    assign _739 = _7677;
    always @(posedge _1038) begin
        if (_1036)
            _7674 <= _1055;
        else
            _7674 <= _739;
    end
    assign _7679 = _1062 == _3070;
    assign _7680 = _1059 & _7679;
    assign _7684 = _7680 ? _1029 : _7683;
    assign _7686 = _1047 ? _1055 : _7684;
    assign _740 = _7686;
    always @(posedge _1038) begin
        if (_1036)
            _7683 <= _1055;
        else
            _7683 <= _740;
    end
    assign _7688 = _1062 == _3079;
    assign _7689 = _1059 & _7688;
    assign _7693 = _7689 ? _1029 : _7692;
    assign _7695 = _1047 ? _1055 : _7693;
    assign _741 = _7695;
    always @(posedge _1038) begin
        if (_1036)
            _7692 <= _1055;
        else
            _7692 <= _741;
    end
    assign _7697 = _1062 == _3088;
    assign _7698 = _1059 & _7697;
    assign _7702 = _7698 ? _1029 : _7701;
    assign _7704 = _1047 ? _1055 : _7702;
    assign _742 = _7704;
    always @(posedge _1038) begin
        if (_1036)
            _7701 <= _1055;
        else
            _7701 <= _742;
    end
    assign _7706 = _1062 == _3097;
    assign _7707 = _1059 & _7706;
    assign _7711 = _7707 ? _1029 : _7710;
    assign _7713 = _1047 ? _1055 : _7711;
    assign _743 = _7713;
    always @(posedge _1038) begin
        if (_1036)
            _7710 <= _1055;
        else
            _7710 <= _743;
    end
    assign _7715 = _1062 == _3106;
    assign _7716 = _1059 & _7715;
    assign _7720 = _7716 ? _1029 : _7719;
    assign _7722 = _1047 ? _1055 : _7720;
    assign _744 = _7722;
    always @(posedge _1038) begin
        if (_1036)
            _7719 <= _1055;
        else
            _7719 <= _744;
    end
    assign _7724 = _1062 == _3115;
    assign _7725 = _1059 & _7724;
    assign _7729 = _7725 ? _1029 : _7728;
    assign _7731 = _1047 ? _1055 : _7729;
    assign _745 = _7731;
    always @(posedge _1038) begin
        if (_1036)
            _7728 <= _1055;
        else
            _7728 <= _745;
    end
    assign _7733 = _1062 == _3124;
    assign _7734 = _1059 & _7733;
    assign _7738 = _7734 ? _1029 : _7737;
    assign _7740 = _1047 ? _1055 : _7738;
    assign _746 = _7740;
    always @(posedge _1038) begin
        if (_1036)
            _7737 <= _1055;
        else
            _7737 <= _746;
    end
    assign _7742 = _1062 == _3133;
    assign _7743 = _1059 & _7742;
    assign _7747 = _7743 ? _1029 : _7746;
    assign _7749 = _1047 ? _1055 : _7747;
    assign _747 = _7749;
    always @(posedge _1038) begin
        if (_1036)
            _7746 <= _1055;
        else
            _7746 <= _747;
    end
    assign _7751 = _1062 == _3142;
    assign _7752 = _1059 & _7751;
    assign _7756 = _7752 ? _1029 : _7755;
    assign _7758 = _1047 ? _1055 : _7756;
    assign _748 = _7758;
    always @(posedge _1038) begin
        if (_1036)
            _7755 <= _1055;
        else
            _7755 <= _748;
    end
    assign _7760 = _1062 == _3151;
    assign _7761 = _1059 & _7760;
    assign _7765 = _7761 ? _1029 : _7764;
    assign _7767 = _1047 ? _1055 : _7765;
    assign _749 = _7767;
    always @(posedge _1038) begin
        if (_1036)
            _7764 <= _1055;
        else
            _7764 <= _749;
    end
    assign _7769 = _1062 == _3160;
    assign _7770 = _1059 & _7769;
    assign _7774 = _7770 ? _1029 : _7773;
    assign _7776 = _1047 ? _1055 : _7774;
    assign _750 = _7776;
    always @(posedge _1038) begin
        if (_1036)
            _7773 <= _1055;
        else
            _7773 <= _750;
    end
    assign _7778 = _1062 == _3169;
    assign _7779 = _1059 & _7778;
    assign _7783 = _7779 ? _1029 : _7782;
    assign _7785 = _1047 ? _1055 : _7783;
    assign _751 = _7785;
    always @(posedge _1038) begin
        if (_1036)
            _7782 <= _1055;
        else
            _7782 <= _751;
    end
    assign _7787 = _1062 == _3178;
    assign _7788 = _1059 & _7787;
    assign _7792 = _7788 ? _1029 : _7791;
    assign _7794 = _1047 ? _1055 : _7792;
    assign _752 = _7794;
    always @(posedge _1038) begin
        if (_1036)
            _7791 <= _1055;
        else
            _7791 <= _752;
    end
    assign _7796 = _1062 == _3187;
    assign _7797 = _1059 & _7796;
    assign _7801 = _7797 ? _1029 : _7800;
    assign _7803 = _1047 ? _1055 : _7801;
    assign _753 = _7803;
    always @(posedge _1038) begin
        if (_1036)
            _7800 <= _1055;
        else
            _7800 <= _753;
    end
    assign _7805 = _1062 == _3196;
    assign _7806 = _1059 & _7805;
    assign _7810 = _7806 ? _1029 : _7809;
    assign _7812 = _1047 ? _1055 : _7810;
    assign _754 = _7812;
    always @(posedge _1038) begin
        if (_1036)
            _7809 <= _1055;
        else
            _7809 <= _754;
    end
    assign _7814 = _1062 == _3205;
    assign _7815 = _1059 & _7814;
    assign _7819 = _7815 ? _1029 : _7818;
    assign _7821 = _1047 ? _1055 : _7819;
    assign _755 = _7821;
    always @(posedge _1038) begin
        if (_1036)
            _7818 <= _1055;
        else
            _7818 <= _755;
    end
    assign _7823 = _1062 == _3214;
    assign _7824 = _1059 & _7823;
    assign _7828 = _7824 ? _1029 : _7827;
    assign _7830 = _1047 ? _1055 : _7828;
    assign _756 = _7830;
    always @(posedge _1038) begin
        if (_1036)
            _7827 <= _1055;
        else
            _7827 <= _756;
    end
    assign _7832 = _1062 == _3223;
    assign _7833 = _1059 & _7832;
    assign _7837 = _7833 ? _1029 : _7836;
    assign _7839 = _1047 ? _1055 : _7837;
    assign _757 = _7839;
    always @(posedge _1038) begin
        if (_1036)
            _7836 <= _1055;
        else
            _7836 <= _757;
    end
    assign _7841 = _1062 == _3232;
    assign _7842 = _1059 & _7841;
    assign _7846 = _7842 ? _1029 : _7845;
    assign _7848 = _1047 ? _1055 : _7846;
    assign _758 = _7848;
    always @(posedge _1038) begin
        if (_1036)
            _7845 <= _1055;
        else
            _7845 <= _758;
    end
    assign _7850 = _1062 == _3241;
    assign _7851 = _1059 & _7850;
    assign _7855 = _7851 ? _1029 : _7854;
    assign _7857 = _1047 ? _1055 : _7855;
    assign _759 = _7857;
    always @(posedge _1038) begin
        if (_1036)
            _7854 <= _1055;
        else
            _7854 <= _759;
    end
    assign _7859 = _1062 == _3250;
    assign _7860 = _1059 & _7859;
    assign _7864 = _7860 ? _1029 : _7863;
    assign _7866 = _1047 ? _1055 : _7864;
    assign _760 = _7866;
    always @(posedge _1038) begin
        if (_1036)
            _7863 <= _1055;
        else
            _7863 <= _760;
    end
    assign _7868 = _1062 == _3259;
    assign _7869 = _1059 & _7868;
    assign _7873 = _7869 ? _1029 : _7872;
    assign _7875 = _1047 ? _1055 : _7873;
    assign _761 = _7875;
    always @(posedge _1038) begin
        if (_1036)
            _7872 <= _1055;
        else
            _7872 <= _761;
    end
    assign _7877 = _1062 == _3268;
    assign _7878 = _1059 & _7877;
    assign _7882 = _7878 ? _1029 : _7881;
    assign _7884 = _1047 ? _1055 : _7882;
    assign _762 = _7884;
    always @(posedge _1038) begin
        if (_1036)
            _7881 <= _1055;
        else
            _7881 <= _762;
    end
    assign _7886 = _1062 == _3277;
    assign _7887 = _1059 & _7886;
    assign _7891 = _7887 ? _1029 : _7890;
    assign _7893 = _1047 ? _1055 : _7891;
    assign _763 = _7893;
    always @(posedge _1038) begin
        if (_1036)
            _7890 <= _1055;
        else
            _7890 <= _763;
    end
    assign _7895 = _1062 == _3286;
    assign _7896 = _1059 & _7895;
    assign _7900 = _7896 ? _1029 : _7899;
    assign _7902 = _1047 ? _1055 : _7900;
    assign _764 = _7902;
    always @(posedge _1038) begin
        if (_1036)
            _7899 <= _1055;
        else
            _7899 <= _764;
    end
    assign _7904 = _1062 == _3295;
    assign _7905 = _1059 & _7904;
    assign _7909 = _7905 ? _1029 : _7908;
    assign _7911 = _1047 ? _1055 : _7909;
    assign _765 = _7911;
    always @(posedge _1038) begin
        if (_1036)
            _7908 <= _1055;
        else
            _7908 <= _765;
    end
    assign _7913 = _1062 == _3304;
    assign _7914 = _1059 & _7913;
    assign _7918 = _7914 ? _1029 : _7917;
    assign _7920 = _1047 ? _1055 : _7918;
    assign _766 = _7920;
    always @(posedge _1038) begin
        if (_1036)
            _7917 <= _1055;
        else
            _7917 <= _766;
    end
    assign _7922 = _1062 == _3313;
    assign _7923 = _1059 & _7922;
    assign _7927 = _7923 ? _1029 : _7926;
    assign _7929 = _1047 ? _1055 : _7927;
    assign _767 = _7929;
    always @(posedge _1038) begin
        if (_1036)
            _7926 <= _1055;
        else
            _7926 <= _767;
    end
    assign _7931 = _1062 == _3322;
    assign _7932 = _1059 & _7931;
    assign _7936 = _7932 ? _1029 : _7935;
    assign _7938 = _1047 ? _1055 : _7936;
    assign _768 = _7938;
    always @(posedge _1038) begin
        if (_1036)
            _7935 <= _1055;
        else
            _7935 <= _768;
    end
    assign _7940 = _1062 == _3331;
    assign _7941 = _1059 & _7940;
    assign _7945 = _7941 ? _1029 : _7944;
    assign _7947 = _1047 ? _1055 : _7945;
    assign _769 = _7947;
    always @(posedge _1038) begin
        if (_1036)
            _7944 <= _1055;
        else
            _7944 <= _769;
    end
    assign _7949 = _1062 == _3340;
    assign _7950 = _1059 & _7949;
    assign _7954 = _7950 ? _1029 : _7953;
    assign _7956 = _1047 ? _1055 : _7954;
    assign _770 = _7956;
    always @(posedge _1038) begin
        if (_1036)
            _7953 <= _1055;
        else
            _7953 <= _770;
    end
    assign _7958 = _1062 == _3349;
    assign _7959 = _1059 & _7958;
    assign _7963 = _7959 ? _1029 : _7962;
    assign _7965 = _1047 ? _1055 : _7963;
    assign _771 = _7965;
    always @(posedge _1038) begin
        if (_1036)
            _7962 <= _1055;
        else
            _7962 <= _771;
    end
    assign _7967 = _1062 == _3358;
    assign _7968 = _1059 & _7967;
    assign _7972 = _7968 ? _1029 : _7971;
    assign _7974 = _1047 ? _1055 : _7972;
    assign _772 = _7974;
    always @(posedge _1038) begin
        if (_1036)
            _7971 <= _1055;
        else
            _7971 <= _772;
    end
    assign _7976 = _1062 == _3367;
    assign _7977 = _1059 & _7976;
    assign _7981 = _7977 ? _1029 : _7980;
    assign _7983 = _1047 ? _1055 : _7981;
    assign _773 = _7983;
    always @(posedge _1038) begin
        if (_1036)
            _7980 <= _1055;
        else
            _7980 <= _773;
    end
    assign _7985 = _1062 == _3376;
    assign _7986 = _1059 & _7985;
    assign _7990 = _7986 ? _1029 : _7989;
    assign _7992 = _1047 ? _1055 : _7990;
    assign _774 = _7992;
    always @(posedge _1038) begin
        if (_1036)
            _7989 <= _1055;
        else
            _7989 <= _774;
    end
    assign _7994 = _1062 == _3385;
    assign _7995 = _1059 & _7994;
    assign _7999 = _7995 ? _1029 : _7998;
    assign _8001 = _1047 ? _1055 : _7999;
    assign _775 = _8001;
    always @(posedge _1038) begin
        if (_1036)
            _7998 <= _1055;
        else
            _7998 <= _775;
    end
    assign _8003 = _1062 == _3394;
    assign _8004 = _1059 & _8003;
    assign _8008 = _8004 ? _1029 : _8007;
    assign _8010 = _1047 ? _1055 : _8008;
    assign _776 = _8010;
    always @(posedge _1038) begin
        if (_1036)
            _8007 <= _1055;
        else
            _8007 <= _776;
    end
    assign _8012 = _1062 == _3403;
    assign _8013 = _1059 & _8012;
    assign _8017 = _8013 ? _1029 : _8016;
    assign _8019 = _1047 ? _1055 : _8017;
    assign _777 = _8019;
    always @(posedge _1038) begin
        if (_1036)
            _8016 <= _1055;
        else
            _8016 <= _777;
    end
    assign _8021 = _1062 == _3412;
    assign _8022 = _1059 & _8021;
    assign _8026 = _8022 ? _1029 : _8025;
    assign _8028 = _1047 ? _1055 : _8026;
    assign _778 = _8028;
    always @(posedge _1038) begin
        if (_1036)
            _8025 <= _1055;
        else
            _8025 <= _778;
    end
    assign _8030 = _1062 == _3421;
    assign _8031 = _1059 & _8030;
    assign _8035 = _8031 ? _1029 : _8034;
    assign _8037 = _1047 ? _1055 : _8035;
    assign _779 = _8037;
    always @(posedge _1038) begin
        if (_1036)
            _8034 <= _1055;
        else
            _8034 <= _779;
    end
    assign _8039 = _1062 == _3430;
    assign _8040 = _1059 & _8039;
    assign _8044 = _8040 ? _1029 : _8043;
    assign _8046 = _1047 ? _1055 : _8044;
    assign _780 = _8046;
    always @(posedge _1038) begin
        if (_1036)
            _8043 <= _1055;
        else
            _8043 <= _780;
    end
    assign _8048 = _1062 == _3439;
    assign _8049 = _1059 & _8048;
    assign _8053 = _8049 ? _1029 : _8052;
    assign _8055 = _1047 ? _1055 : _8053;
    assign _781 = _8055;
    always @(posedge _1038) begin
        if (_1036)
            _8052 <= _1055;
        else
            _8052 <= _781;
    end
    assign _8057 = _1062 == _3448;
    assign _8058 = _1059 & _8057;
    assign _8062 = _8058 ? _1029 : _8061;
    assign _8064 = _1047 ? _1055 : _8062;
    assign _782 = _8064;
    always @(posedge _1038) begin
        if (_1036)
            _8061 <= _1055;
        else
            _8061 <= _782;
    end
    assign _8066 = _1062 == _3457;
    assign _8067 = _1059 & _8066;
    assign _8071 = _8067 ? _1029 : _8070;
    assign _8073 = _1047 ? _1055 : _8071;
    assign _783 = _8073;
    always @(posedge _1038) begin
        if (_1036)
            _8070 <= _1055;
        else
            _8070 <= _783;
    end
    assign _8075 = _1062 == _3466;
    assign _8076 = _1059 & _8075;
    assign _8080 = _8076 ? _1029 : _8079;
    assign _8082 = _1047 ? _1055 : _8080;
    assign _784 = _8082;
    always @(posedge _1038) begin
        if (_1036)
            _8079 <= _1055;
        else
            _8079 <= _784;
    end
    assign _8084 = _1062 == _3475;
    assign _8085 = _1059 & _8084;
    assign _8089 = _8085 ? _1029 : _8088;
    assign _8091 = _1047 ? _1055 : _8089;
    assign _785 = _8091;
    always @(posedge _1038) begin
        if (_1036)
            _8088 <= _1055;
        else
            _8088 <= _785;
    end
    assign _8093 = _1062 == _3484;
    assign _8094 = _1059 & _8093;
    assign _8098 = _8094 ? _1029 : _8097;
    assign _8100 = _1047 ? _1055 : _8098;
    assign _786 = _8100;
    always @(posedge _1038) begin
        if (_1036)
            _8097 <= _1055;
        else
            _8097 <= _786;
    end
    assign _8102 = _1062 == _3493;
    assign _8103 = _1059 & _8102;
    assign _8107 = _8103 ? _1029 : _8106;
    assign _8109 = _1047 ? _1055 : _8107;
    assign _787 = _8109;
    always @(posedge _1038) begin
        if (_1036)
            _8106 <= _1055;
        else
            _8106 <= _787;
    end
    assign _8111 = _1062 == _3502;
    assign _8112 = _1059 & _8111;
    assign _8116 = _8112 ? _1029 : _8115;
    assign _8118 = _1047 ? _1055 : _8116;
    assign _788 = _8118;
    always @(posedge _1038) begin
        if (_1036)
            _8115 <= _1055;
        else
            _8115 <= _788;
    end
    assign _8120 = _1062 == _3511;
    assign _8121 = _1059 & _8120;
    assign _8125 = _8121 ? _1029 : _8124;
    assign _8127 = _1047 ? _1055 : _8125;
    assign _789 = _8127;
    always @(posedge _1038) begin
        if (_1036)
            _8124 <= _1055;
        else
            _8124 <= _789;
    end
    assign _8129 = _1062 == _3520;
    assign _8130 = _1059 & _8129;
    assign _8134 = _8130 ? _1029 : _8133;
    assign _8136 = _1047 ? _1055 : _8134;
    assign _790 = _8136;
    always @(posedge _1038) begin
        if (_1036)
            _8133 <= _1055;
        else
            _8133 <= _790;
    end
    assign _8138 = _1062 == _3529;
    assign _8139 = _1059 & _8138;
    assign _8143 = _8139 ? _1029 : _8142;
    assign _8145 = _1047 ? _1055 : _8143;
    assign _791 = _8145;
    always @(posedge _1038) begin
        if (_1036)
            _8142 <= _1055;
        else
            _8142 <= _791;
    end
    assign _8147 = _1062 == _3538;
    assign _8148 = _1059 & _8147;
    assign _8152 = _8148 ? _1029 : _8151;
    assign _8154 = _1047 ? _1055 : _8152;
    assign _792 = _8154;
    always @(posedge _1038) begin
        if (_1036)
            _8151 <= _1055;
        else
            _8151 <= _792;
    end
    assign _8156 = _1062 == _3547;
    assign _8157 = _1059 & _8156;
    assign _8161 = _8157 ? _1029 : _8160;
    assign _8163 = _1047 ? _1055 : _8161;
    assign _793 = _8163;
    always @(posedge _1038) begin
        if (_1036)
            _8160 <= _1055;
        else
            _8160 <= _793;
    end
    assign _8165 = _1062 == _3556;
    assign _8166 = _1059 & _8165;
    assign _8170 = _8166 ? _1029 : _8169;
    assign _8172 = _1047 ? _1055 : _8170;
    assign _794 = _8172;
    always @(posedge _1038) begin
        if (_1036)
            _8169 <= _1055;
        else
            _8169 <= _794;
    end
    assign _8174 = _1062 == _3565;
    assign _8175 = _1059 & _8174;
    assign _8179 = _8175 ? _1029 : _8178;
    assign _8181 = _1047 ? _1055 : _8179;
    assign _795 = _8181;
    always @(posedge _1038) begin
        if (_1036)
            _8178 <= _1055;
        else
            _8178 <= _795;
    end
    assign _8183 = _1062 == _3574;
    assign _8184 = _1059 & _8183;
    assign _8188 = _8184 ? _1029 : _8187;
    assign _8190 = _1047 ? _1055 : _8188;
    assign _796 = _8190;
    always @(posedge _1038) begin
        if (_1036)
            _8187 <= _1055;
        else
            _8187 <= _796;
    end
    assign _8192 = _1062 == _3583;
    assign _8193 = _1059 & _8192;
    assign _8197 = _8193 ? _1029 : _8196;
    assign _8199 = _1047 ? _1055 : _8197;
    assign _797 = _8199;
    always @(posedge _1038) begin
        if (_1036)
            _8196 <= _1055;
        else
            _8196 <= _797;
    end
    assign _8201 = _1062 == _3592;
    assign _8202 = _1059 & _8201;
    assign _8206 = _8202 ? _1029 : _8205;
    assign _8208 = _1047 ? _1055 : _8206;
    assign _798 = _8208;
    always @(posedge _1038) begin
        if (_1036)
            _8205 <= _1055;
        else
            _8205 <= _798;
    end
    assign _8210 = _1062 == _3601;
    assign _8211 = _1059 & _8210;
    assign _8215 = _8211 ? _1029 : _8214;
    assign _8217 = _1047 ? _1055 : _8215;
    assign _799 = _8217;
    always @(posedge _1038) begin
        if (_1036)
            _8214 <= _1055;
        else
            _8214 <= _799;
    end
    assign _8219 = _1062 == _3610;
    assign _8220 = _1059 & _8219;
    assign _8224 = _8220 ? _1029 : _8223;
    assign _8226 = _1047 ? _1055 : _8224;
    assign _800 = _8226;
    always @(posedge _1038) begin
        if (_1036)
            _8223 <= _1055;
        else
            _8223 <= _800;
    end
    assign _8228 = _1062 == _3619;
    assign _8229 = _1059 & _8228;
    assign _8233 = _8229 ? _1029 : _8232;
    assign _8235 = _1047 ? _1055 : _8233;
    assign _801 = _8235;
    always @(posedge _1038) begin
        if (_1036)
            _8232 <= _1055;
        else
            _8232 <= _801;
    end
    assign _8237 = _1062 == _3628;
    assign _8238 = _1059 & _8237;
    assign _8242 = _8238 ? _1029 : _8241;
    assign _8244 = _1047 ? _1055 : _8242;
    assign _802 = _8244;
    always @(posedge _1038) begin
        if (_1036)
            _8241 <= _1055;
        else
            _8241 <= _802;
    end
    assign _8246 = _1062 == _3637;
    assign _8247 = _1059 & _8246;
    assign _8251 = _8247 ? _1029 : _8250;
    assign _8253 = _1047 ? _1055 : _8251;
    assign _803 = _8253;
    always @(posedge _1038) begin
        if (_1036)
            _8250 <= _1055;
        else
            _8250 <= _803;
    end
    assign _8255 = _1062 == _3646;
    assign _8256 = _1059 & _8255;
    assign _8260 = _8256 ? _1029 : _8259;
    assign _8262 = _1047 ? _1055 : _8260;
    assign _804 = _8262;
    always @(posedge _1038) begin
        if (_1036)
            _8259 <= _1055;
        else
            _8259 <= _804;
    end
    assign _8264 = _1062 == _3655;
    assign _8265 = _1059 & _8264;
    assign _8269 = _8265 ? _1029 : _8268;
    assign _8271 = _1047 ? _1055 : _8269;
    assign _805 = _8271;
    always @(posedge _1038) begin
        if (_1036)
            _8268 <= _1055;
        else
            _8268 <= _805;
    end
    assign _8273 = _1062 == _3664;
    assign _8274 = _1059 & _8273;
    assign _8278 = _8274 ? _1029 : _8277;
    assign _8280 = _1047 ? _1055 : _8278;
    assign _806 = _8280;
    always @(posedge _1038) begin
        if (_1036)
            _8277 <= _1055;
        else
            _8277 <= _806;
    end
    assign _8282 = _1062 == _3673;
    assign _8283 = _1059 & _8282;
    assign _8287 = _8283 ? _1029 : _8286;
    assign _8289 = _1047 ? _1055 : _8287;
    assign _807 = _8289;
    always @(posedge _1038) begin
        if (_1036)
            _8286 <= _1055;
        else
            _8286 <= _807;
    end
    assign _8291 = _1062 == _3682;
    assign _8292 = _1059 & _8291;
    assign _8296 = _8292 ? _1029 : _8295;
    assign _8298 = _1047 ? _1055 : _8296;
    assign _808 = _8298;
    always @(posedge _1038) begin
        if (_1036)
            _8295 <= _1055;
        else
            _8295 <= _808;
    end
    assign _8300 = _1062 == _3691;
    assign _8301 = _1059 & _8300;
    assign _8305 = _8301 ? _1029 : _8304;
    assign _8307 = _1047 ? _1055 : _8305;
    assign _809 = _8307;
    always @(posedge _1038) begin
        if (_1036)
            _8304 <= _1055;
        else
            _8304 <= _809;
    end
    assign _8309 = _1062 == _3700;
    assign _8310 = _1059 & _8309;
    assign _8314 = _8310 ? _1029 : _8313;
    assign _8316 = _1047 ? _1055 : _8314;
    assign _810 = _8316;
    always @(posedge _1038) begin
        if (_1036)
            _8313 <= _1055;
        else
            _8313 <= _810;
    end
    assign _8318 = _1062 == _3709;
    assign _8319 = _1059 & _8318;
    assign _8323 = _8319 ? _1029 : _8322;
    assign _8325 = _1047 ? _1055 : _8323;
    assign _811 = _8325;
    always @(posedge _1038) begin
        if (_1036)
            _8322 <= _1055;
        else
            _8322 <= _811;
    end
    assign _8327 = _1062 == _3718;
    assign _8328 = _1059 & _8327;
    assign _8332 = _8328 ? _1029 : _8331;
    assign _8334 = _1047 ? _1055 : _8332;
    assign _812 = _8334;
    always @(posedge _1038) begin
        if (_1036)
            _8331 <= _1055;
        else
            _8331 <= _812;
    end
    assign _8336 = _1062 == _3727;
    assign _8337 = _1059 & _8336;
    assign _8341 = _8337 ? _1029 : _8340;
    assign _8343 = _1047 ? _1055 : _8341;
    assign _813 = _8343;
    always @(posedge _1038) begin
        if (_1036)
            _8340 <= _1055;
        else
            _8340 <= _813;
    end
    assign _8345 = _1062 == _3736;
    assign _8346 = _1059 & _8345;
    assign _8350 = _8346 ? _1029 : _8349;
    assign _8352 = _1047 ? _1055 : _8350;
    assign _814 = _8352;
    always @(posedge _1038) begin
        if (_1036)
            _8349 <= _1055;
        else
            _8349 <= _814;
    end
    assign _8354 = _1062 == _3745;
    assign _8355 = _1059 & _8354;
    assign _8359 = _8355 ? _1029 : _8358;
    assign _8361 = _1047 ? _1055 : _8359;
    assign _815 = _8361;
    always @(posedge _1038) begin
        if (_1036)
            _8358 <= _1055;
        else
            _8358 <= _815;
    end
    assign _8363 = _1062 == _3754;
    assign _8364 = _1059 & _8363;
    assign _8368 = _8364 ? _1029 : _8367;
    assign _8370 = _1047 ? _1055 : _8368;
    assign _816 = _8370;
    always @(posedge _1038) begin
        if (_1036)
            _8367 <= _1055;
        else
            _8367 <= _816;
    end
    assign _8372 = _1062 == _3763;
    assign _8373 = _1059 & _8372;
    assign _8377 = _8373 ? _1029 : _8376;
    assign _8379 = _1047 ? _1055 : _8377;
    assign _817 = _8379;
    always @(posedge _1038) begin
        if (_1036)
            _8376 <= _1055;
        else
            _8376 <= _817;
    end
    assign _8381 = _1062 == _3772;
    assign _8382 = _1059 & _8381;
    assign _8386 = _8382 ? _1029 : _8385;
    assign _8388 = _1047 ? _1055 : _8386;
    assign _818 = _8388;
    always @(posedge _1038) begin
        if (_1036)
            _8385 <= _1055;
        else
            _8385 <= _818;
    end
    assign _8390 = _1062 == _3781;
    assign _8391 = _1059 & _8390;
    assign _8395 = _8391 ? _1029 : _8394;
    assign _8397 = _1047 ? _1055 : _8395;
    assign _819 = _8397;
    always @(posedge _1038) begin
        if (_1036)
            _8394 <= _1055;
        else
            _8394 <= _819;
    end
    assign _8399 = _1062 == _3790;
    assign _8400 = _1059 & _8399;
    assign _8404 = _8400 ? _1029 : _8403;
    assign _8406 = _1047 ? _1055 : _8404;
    assign _820 = _8406;
    always @(posedge _1038) begin
        if (_1036)
            _8403 <= _1055;
        else
            _8403 <= _820;
    end
    assign _8408 = _1062 == _3799;
    assign _8409 = _1059 & _8408;
    assign _8413 = _8409 ? _1029 : _8412;
    assign _8415 = _1047 ? _1055 : _8413;
    assign _821 = _8415;
    always @(posedge _1038) begin
        if (_1036)
            _8412 <= _1055;
        else
            _8412 <= _821;
    end
    assign _8417 = _1062 == _3808;
    assign _8418 = _1059 & _8417;
    assign _8422 = _8418 ? _1029 : _8421;
    assign _8424 = _1047 ? _1055 : _8422;
    assign _822 = _8424;
    always @(posedge _1038) begin
        if (_1036)
            _8421 <= _1055;
        else
            _8421 <= _822;
    end
    assign _8426 = _1062 == _3817;
    assign _8427 = _1059 & _8426;
    assign _8431 = _8427 ? _1029 : _8430;
    assign _8433 = _1047 ? _1055 : _8431;
    assign _823 = _8433;
    always @(posedge _1038) begin
        if (_1036)
            _8430 <= _1055;
        else
            _8430 <= _823;
    end
    assign _8435 = _1062 == _3826;
    assign _8436 = _1059 & _8435;
    assign _8440 = _8436 ? _1029 : _8439;
    assign _8442 = _1047 ? _1055 : _8440;
    assign _824 = _8442;
    always @(posedge _1038) begin
        if (_1036)
            _8439 <= _1055;
        else
            _8439 <= _824;
    end
    assign _8444 = _1062 == _3835;
    assign _8445 = _1059 & _8444;
    assign _8449 = _8445 ? _1029 : _8448;
    assign _8451 = _1047 ? _1055 : _8449;
    assign _825 = _8451;
    always @(posedge _1038) begin
        if (_1036)
            _8448 <= _1055;
        else
            _8448 <= _825;
    end
    assign _8453 = _1062 == _3844;
    assign _8454 = _1059 & _8453;
    assign _8458 = _8454 ? _1029 : _8457;
    assign _8460 = _1047 ? _1055 : _8458;
    assign _826 = _8460;
    always @(posedge _1038) begin
        if (_1036)
            _8457 <= _1055;
        else
            _8457 <= _826;
    end
    assign _8462 = _1062 == _3853;
    assign _8463 = _1059 & _8462;
    assign _8467 = _8463 ? _1029 : _8466;
    assign _8469 = _1047 ? _1055 : _8467;
    assign _827 = _8469;
    always @(posedge _1038) begin
        if (_1036)
            _8466 <= _1055;
        else
            _8466 <= _827;
    end
    assign _8471 = _1062 == _3862;
    assign _8472 = _1059 & _8471;
    assign _8476 = _8472 ? _1029 : _8475;
    assign _8478 = _1047 ? _1055 : _8476;
    assign _828 = _8478;
    always @(posedge _1038) begin
        if (_1036)
            _8475 <= _1055;
        else
            _8475 <= _828;
    end
    assign _8480 = _1062 == _3871;
    assign _8481 = _1059 & _8480;
    assign _8485 = _8481 ? _1029 : _8484;
    assign _8487 = _1047 ? _1055 : _8485;
    assign _829 = _8487;
    always @(posedge _1038) begin
        if (_1036)
            _8484 <= _1055;
        else
            _8484 <= _829;
    end
    assign _8489 = _1062 == _3880;
    assign _8490 = _1059 & _8489;
    assign _8494 = _8490 ? _1029 : _8493;
    assign _8496 = _1047 ? _1055 : _8494;
    assign _830 = _8496;
    always @(posedge _1038) begin
        if (_1036)
            _8493 <= _1055;
        else
            _8493 <= _830;
    end
    assign _8498 = _1062 == _3889;
    assign _8499 = _1059 & _8498;
    assign _8503 = _8499 ? _1029 : _8502;
    assign _8505 = _1047 ? _1055 : _8503;
    assign _831 = _8505;
    always @(posedge _1038) begin
        if (_1036)
            _8502 <= _1055;
        else
            _8502 <= _831;
    end
    assign _8507 = _1062 == _3898;
    assign _8508 = _1059 & _8507;
    assign _8512 = _8508 ? _1029 : _8511;
    assign _8514 = _1047 ? _1055 : _8512;
    assign _832 = _8514;
    always @(posedge _1038) begin
        if (_1036)
            _8511 <= _1055;
        else
            _8511 <= _832;
    end
    assign _8516 = _1062 == _3907;
    assign _8517 = _1059 & _8516;
    assign _8521 = _8517 ? _1029 : _8520;
    assign _8523 = _1047 ? _1055 : _8521;
    assign _833 = _8523;
    always @(posedge _1038) begin
        if (_1036)
            _8520 <= _1055;
        else
            _8520 <= _833;
    end
    assign _8525 = _1062 == _3916;
    assign _8526 = _1059 & _8525;
    assign _8530 = _8526 ? _1029 : _8529;
    assign _8532 = _1047 ? _1055 : _8530;
    assign _834 = _8532;
    always @(posedge _1038) begin
        if (_1036)
            _8529 <= _1055;
        else
            _8529 <= _834;
    end
    assign _8534 = _1062 == _3925;
    assign _8535 = _1059 & _8534;
    assign _8539 = _8535 ? _1029 : _8538;
    assign _8541 = _1047 ? _1055 : _8539;
    assign _835 = _8541;
    always @(posedge _1038) begin
        if (_1036)
            _8538 <= _1055;
        else
            _8538 <= _835;
    end
    assign _8543 = _1062 == _3934;
    assign _8544 = _1059 & _8543;
    assign _8548 = _8544 ? _1029 : _8547;
    assign _8550 = _1047 ? _1055 : _8548;
    assign _836 = _8550;
    always @(posedge _1038) begin
        if (_1036)
            _8547 <= _1055;
        else
            _8547 <= _836;
    end
    assign _8552 = _1062 == _3943;
    assign _8553 = _1059 & _8552;
    assign _8557 = _8553 ? _1029 : _8556;
    assign _8559 = _1047 ? _1055 : _8557;
    assign _837 = _8559;
    always @(posedge _1038) begin
        if (_1036)
            _8556 <= _1055;
        else
            _8556 <= _837;
    end
    assign _8561 = _1062 == _3952;
    assign _8562 = _1059 & _8561;
    assign _8566 = _8562 ? _1029 : _8565;
    assign _8568 = _1047 ? _1055 : _8566;
    assign _838 = _8568;
    always @(posedge _1038) begin
        if (_1036)
            _8565 <= _1055;
        else
            _8565 <= _838;
    end
    assign _8570 = _1062 == _3961;
    assign _8571 = _1059 & _8570;
    assign _8575 = _8571 ? _1029 : _8574;
    assign _8577 = _1047 ? _1055 : _8575;
    assign _839 = _8577;
    always @(posedge _1038) begin
        if (_1036)
            _8574 <= _1055;
        else
            _8574 <= _839;
    end
    assign _8579 = _1062 == _3970;
    assign _8580 = _1059 & _8579;
    assign _8584 = _8580 ? _1029 : _8583;
    assign _8586 = _1047 ? _1055 : _8584;
    assign _840 = _8586;
    always @(posedge _1038) begin
        if (_1036)
            _8583 <= _1055;
        else
            _8583 <= _840;
    end
    assign _8588 = _1062 == _3979;
    assign _8589 = _1059 & _8588;
    assign _8593 = _8589 ? _1029 : _8592;
    assign _8595 = _1047 ? _1055 : _8593;
    assign _841 = _8595;
    always @(posedge _1038) begin
        if (_1036)
            _8592 <= _1055;
        else
            _8592 <= _841;
    end
    assign _8597 = _1062 == _3988;
    assign _8598 = _1059 & _8597;
    assign _8602 = _8598 ? _1029 : _8601;
    assign _8604 = _1047 ? _1055 : _8602;
    assign _842 = _8604;
    always @(posedge _1038) begin
        if (_1036)
            _8601 <= _1055;
        else
            _8601 <= _842;
    end
    assign _8606 = _1062 == _3997;
    assign _8607 = _1059 & _8606;
    assign _8611 = _8607 ? _1029 : _8610;
    assign _8613 = _1047 ? _1055 : _8611;
    assign _843 = _8613;
    always @(posedge _1038) begin
        if (_1036)
            _8610 <= _1055;
        else
            _8610 <= _843;
    end
    assign _8615 = _1062 == _4006;
    assign _8616 = _1059 & _8615;
    assign _8620 = _8616 ? _1029 : _8619;
    assign _8622 = _1047 ? _1055 : _8620;
    assign _844 = _8622;
    always @(posedge _1038) begin
        if (_1036)
            _8619 <= _1055;
        else
            _8619 <= _844;
    end
    assign _8624 = _1062 == _4015;
    assign _8625 = _1059 & _8624;
    assign _8629 = _8625 ? _1029 : _8628;
    assign _8631 = _1047 ? _1055 : _8629;
    assign _845 = _8631;
    always @(posedge _1038) begin
        if (_1036)
            _8628 <= _1055;
        else
            _8628 <= _845;
    end
    assign _8633 = _1062 == _4024;
    assign _8634 = _1059 & _8633;
    assign _8638 = _8634 ? _1029 : _8637;
    assign _8640 = _1047 ? _1055 : _8638;
    assign _846 = _8640;
    always @(posedge _1038) begin
        if (_1036)
            _8637 <= _1055;
        else
            _8637 <= _846;
    end
    assign _8642 = _1062 == _4033;
    assign _8643 = _1059 & _8642;
    assign _8647 = _8643 ? _1029 : _8646;
    assign _8649 = _1047 ? _1055 : _8647;
    assign _847 = _8649;
    always @(posedge _1038) begin
        if (_1036)
            _8646 <= _1055;
        else
            _8646 <= _847;
    end
    assign _8651 = _1062 == _4042;
    assign _8652 = _1059 & _8651;
    assign _8656 = _8652 ? _1029 : _8655;
    assign _8658 = _1047 ? _1055 : _8656;
    assign _848 = _8658;
    always @(posedge _1038) begin
        if (_1036)
            _8655 <= _1055;
        else
            _8655 <= _848;
    end
    assign _8660 = _1062 == _4051;
    assign _8661 = _1059 & _8660;
    assign _8665 = _8661 ? _1029 : _8664;
    assign _8667 = _1047 ? _1055 : _8665;
    assign _849 = _8667;
    always @(posedge _1038) begin
        if (_1036)
            _8664 <= _1055;
        else
            _8664 <= _849;
    end
    assign _8669 = _1062 == _4060;
    assign _8670 = _1059 & _8669;
    assign _8674 = _8670 ? _1029 : _8673;
    assign _8676 = _1047 ? _1055 : _8674;
    assign _850 = _8676;
    always @(posedge _1038) begin
        if (_1036)
            _8673 <= _1055;
        else
            _8673 <= _850;
    end
    assign _8678 = _1062 == _4069;
    assign _8679 = _1059 & _8678;
    assign _8683 = _8679 ? _1029 : _8682;
    assign _8685 = _1047 ? _1055 : _8683;
    assign _851 = _8685;
    always @(posedge _1038) begin
        if (_1036)
            _8682 <= _1055;
        else
            _8682 <= _851;
    end
    assign _8687 = _1062 == _4078;
    assign _8688 = _1059 & _8687;
    assign _8692 = _8688 ? _1029 : _8691;
    assign _8694 = _1047 ? _1055 : _8692;
    assign _852 = _8694;
    always @(posedge _1038) begin
        if (_1036)
            _8691 <= _1055;
        else
            _8691 <= _852;
    end
    assign _8696 = _1062 == _4087;
    assign _8697 = _1059 & _8696;
    assign _8701 = _8697 ? _1029 : _8700;
    assign _8703 = _1047 ? _1055 : _8701;
    assign _853 = _8703;
    always @(posedge _1038) begin
        if (_1036)
            _8700 <= _1055;
        else
            _8700 <= _853;
    end
    assign _8705 = _1062 == _4096;
    assign _8706 = _1059 & _8705;
    assign _8710 = _8706 ? _1029 : _8709;
    assign _8712 = _1047 ? _1055 : _8710;
    assign _854 = _8712;
    always @(posedge _1038) begin
        if (_1036)
            _8709 <= _1055;
        else
            _8709 <= _854;
    end
    assign _8714 = _1062 == _4105;
    assign _8715 = _1059 & _8714;
    assign _8719 = _8715 ? _1029 : _8718;
    assign _8721 = _1047 ? _1055 : _8719;
    assign _855 = _8721;
    always @(posedge _1038) begin
        if (_1036)
            _8718 <= _1055;
        else
            _8718 <= _855;
    end
    assign _8723 = _1062 == _4114;
    assign _8724 = _1059 & _8723;
    assign _8728 = _8724 ? _1029 : _8727;
    assign _8730 = _1047 ? _1055 : _8728;
    assign _856 = _8730;
    always @(posedge _1038) begin
        if (_1036)
            _8727 <= _1055;
        else
            _8727 <= _856;
    end
    assign _8732 = _1062 == _4123;
    assign _8733 = _1059 & _8732;
    assign _8737 = _8733 ? _1029 : _8736;
    assign _8739 = _1047 ? _1055 : _8737;
    assign _857 = _8739;
    always @(posedge _1038) begin
        if (_1036)
            _8736 <= _1055;
        else
            _8736 <= _857;
    end
    assign _8741 = _1062 == _4132;
    assign _8742 = _1059 & _8741;
    assign _8746 = _8742 ? _1029 : _8745;
    assign _8748 = _1047 ? _1055 : _8746;
    assign _858 = _8748;
    always @(posedge _1038) begin
        if (_1036)
            _8745 <= _1055;
        else
            _8745 <= _858;
    end
    assign _8750 = _1062 == _4141;
    assign _8751 = _1059 & _8750;
    assign _8755 = _8751 ? _1029 : _8754;
    assign _8757 = _1047 ? _1055 : _8755;
    assign _859 = _8757;
    always @(posedge _1038) begin
        if (_1036)
            _8754 <= _1055;
        else
            _8754 <= _859;
    end
    assign _8759 = _1062 == _4150;
    assign _8760 = _1059 & _8759;
    assign _8764 = _8760 ? _1029 : _8763;
    assign _8766 = _1047 ? _1055 : _8764;
    assign _860 = _8766;
    always @(posedge _1038) begin
        if (_1036)
            _8763 <= _1055;
        else
            _8763 <= _860;
    end
    assign _8768 = _1062 == _4159;
    assign _8769 = _1059 & _8768;
    assign _8773 = _8769 ? _1029 : _8772;
    assign _8775 = _1047 ? _1055 : _8773;
    assign _861 = _8775;
    always @(posedge _1038) begin
        if (_1036)
            _8772 <= _1055;
        else
            _8772 <= _861;
    end
    assign _8777 = _1062 == _4168;
    assign _8778 = _1059 & _8777;
    assign _8782 = _8778 ? _1029 : _8781;
    assign _8784 = _1047 ? _1055 : _8782;
    assign _862 = _8784;
    always @(posedge _1038) begin
        if (_1036)
            _8781 <= _1055;
        else
            _8781 <= _862;
    end
    assign _8786 = _1062 == _4177;
    assign _8787 = _1059 & _8786;
    assign _8791 = _8787 ? _1029 : _8790;
    assign _8793 = _1047 ? _1055 : _8791;
    assign _863 = _8793;
    always @(posedge _1038) begin
        if (_1036)
            _8790 <= _1055;
        else
            _8790 <= _863;
    end
    assign _8795 = _1062 == _4186;
    assign _8796 = _1059 & _8795;
    assign _8800 = _8796 ? _1029 : _8799;
    assign _8802 = _1047 ? _1055 : _8800;
    assign _864 = _8802;
    always @(posedge _1038) begin
        if (_1036)
            _8799 <= _1055;
        else
            _8799 <= _864;
    end
    assign _8804 = _1062 == _4195;
    assign _8805 = _1059 & _8804;
    assign _8809 = _8805 ? _1029 : _8808;
    assign _8811 = _1047 ? _1055 : _8809;
    assign _865 = _8811;
    always @(posedge _1038) begin
        if (_1036)
            _8808 <= _1055;
        else
            _8808 <= _865;
    end
    assign _8813 = _1062 == _4204;
    assign _8814 = _1059 & _8813;
    assign _8818 = _8814 ? _1029 : _8817;
    assign _8820 = _1047 ? _1055 : _8818;
    assign _866 = _8820;
    always @(posedge _1038) begin
        if (_1036)
            _8817 <= _1055;
        else
            _8817 <= _866;
    end
    assign _8822 = _1062 == _4213;
    assign _8823 = _1059 & _8822;
    assign _8827 = _8823 ? _1029 : _8826;
    assign _8829 = _1047 ? _1055 : _8827;
    assign _867 = _8829;
    always @(posedge _1038) begin
        if (_1036)
            _8826 <= _1055;
        else
            _8826 <= _867;
    end
    assign _8831 = _1062 == _4222;
    assign _8832 = _1059 & _8831;
    assign _8836 = _8832 ? _1029 : _8835;
    assign _8838 = _1047 ? _1055 : _8836;
    assign _868 = _8838;
    always @(posedge _1038) begin
        if (_1036)
            _8835 <= _1055;
        else
            _8835 <= _868;
    end
    assign _8840 = _1062 == _4231;
    assign _8841 = _1059 & _8840;
    assign _8845 = _8841 ? _1029 : _8844;
    assign _8847 = _1047 ? _1055 : _8845;
    assign _869 = _8847;
    always @(posedge _1038) begin
        if (_1036)
            _8844 <= _1055;
        else
            _8844 <= _869;
    end
    assign _8849 = _1062 == _4240;
    assign _8850 = _1059 & _8849;
    assign _8854 = _8850 ? _1029 : _8853;
    assign _8856 = _1047 ? _1055 : _8854;
    assign _870 = _8856;
    always @(posedge _1038) begin
        if (_1036)
            _8853 <= _1055;
        else
            _8853 <= _870;
    end
    assign _8858 = _1062 == _4249;
    assign _8859 = _1059 & _8858;
    assign _8863 = _8859 ? _1029 : _8862;
    assign _8865 = _1047 ? _1055 : _8863;
    assign _871 = _8865;
    always @(posedge _1038) begin
        if (_1036)
            _8862 <= _1055;
        else
            _8862 <= _871;
    end
    assign _8867 = _1062 == _4258;
    assign _8868 = _1059 & _8867;
    assign _8872 = _8868 ? _1029 : _8871;
    assign _8874 = _1047 ? _1055 : _8872;
    assign _872 = _8874;
    always @(posedge _1038) begin
        if (_1036)
            _8871 <= _1055;
        else
            _8871 <= _872;
    end
    assign _8876 = _1062 == _4267;
    assign _8877 = _1059 & _8876;
    assign _8881 = _8877 ? _1029 : _8880;
    assign _8883 = _1047 ? _1055 : _8881;
    assign _873 = _8883;
    always @(posedge _1038) begin
        if (_1036)
            _8880 <= _1055;
        else
            _8880 <= _873;
    end
    assign _8885 = _1062 == _4276;
    assign _8886 = _1059 & _8885;
    assign _8890 = _8886 ? _1029 : _8889;
    assign _8892 = _1047 ? _1055 : _8890;
    assign _874 = _8892;
    always @(posedge _1038) begin
        if (_1036)
            _8889 <= _1055;
        else
            _8889 <= _874;
    end
    assign _8894 = _1062 == _4285;
    assign _8895 = _1059 & _8894;
    assign _8899 = _8895 ? _1029 : _8898;
    assign _8901 = _1047 ? _1055 : _8899;
    assign _875 = _8901;
    always @(posedge _1038) begin
        if (_1036)
            _8898 <= _1055;
        else
            _8898 <= _875;
    end
    assign _8903 = _1062 == _4294;
    assign _8904 = _1059 & _8903;
    assign _8908 = _8904 ? _1029 : _8907;
    assign _8910 = _1047 ? _1055 : _8908;
    assign _876 = _8910;
    always @(posedge _1038) begin
        if (_1036)
            _8907 <= _1055;
        else
            _8907 <= _876;
    end
    assign _8912 = _1062 == _4303;
    assign _8913 = _1059 & _8912;
    assign _8917 = _8913 ? _1029 : _8916;
    assign _8919 = _1047 ? _1055 : _8917;
    assign _877 = _8919;
    always @(posedge _1038) begin
        if (_1036)
            _8916 <= _1055;
        else
            _8916 <= _877;
    end
    assign _8921 = _1062 == _4312;
    assign _8922 = _1059 & _8921;
    assign _8926 = _8922 ? _1029 : _8925;
    assign _8928 = _1047 ? _1055 : _8926;
    assign _878 = _8928;
    always @(posedge _1038) begin
        if (_1036)
            _8925 <= _1055;
        else
            _8925 <= _878;
    end
    assign _8930 = _1062 == _4321;
    assign _8931 = _1059 & _8930;
    assign _8935 = _8931 ? _1029 : _8934;
    assign _8937 = _1047 ? _1055 : _8935;
    assign _879 = _8937;
    always @(posedge _1038) begin
        if (_1036)
            _8934 <= _1055;
        else
            _8934 <= _879;
    end
    assign _8939 = _1062 == _4330;
    assign _8940 = _1059 & _8939;
    assign _8944 = _8940 ? _1029 : _8943;
    assign _8946 = _1047 ? _1055 : _8944;
    assign _880 = _8946;
    always @(posedge _1038) begin
        if (_1036)
            _8943 <= _1055;
        else
            _8943 <= _880;
    end
    assign _8948 = _1062 == _4339;
    assign _8949 = _1059 & _8948;
    assign _8953 = _8949 ? _1029 : _8952;
    assign _8955 = _1047 ? _1055 : _8953;
    assign _881 = _8955;
    always @(posedge _1038) begin
        if (_1036)
            _8952 <= _1055;
        else
            _8952 <= _881;
    end
    assign _8957 = _1062 == _4348;
    assign _8958 = _1059 & _8957;
    assign _8962 = _8958 ? _1029 : _8961;
    assign _8964 = _1047 ? _1055 : _8962;
    assign _882 = _8964;
    always @(posedge _1038) begin
        if (_1036)
            _8961 <= _1055;
        else
            _8961 <= _882;
    end
    assign _8966 = _1062 == _4357;
    assign _8967 = _1059 & _8966;
    assign _8971 = _8967 ? _1029 : _8970;
    assign _8973 = _1047 ? _1055 : _8971;
    assign _883 = _8973;
    always @(posedge _1038) begin
        if (_1036)
            _8970 <= _1055;
        else
            _8970 <= _883;
    end
    assign _8975 = _1062 == _4366;
    assign _8976 = _1059 & _8975;
    assign _8980 = _8976 ? _1029 : _8979;
    assign _8982 = _1047 ? _1055 : _8980;
    assign _884 = _8982;
    always @(posedge _1038) begin
        if (_1036)
            _8979 <= _1055;
        else
            _8979 <= _884;
    end
    assign _8984 = _1062 == _4375;
    assign _8985 = _1059 & _8984;
    assign _8989 = _8985 ? _1029 : _8988;
    assign _8991 = _1047 ? _1055 : _8989;
    assign _885 = _8991;
    always @(posedge _1038) begin
        if (_1036)
            _8988 <= _1055;
        else
            _8988 <= _885;
    end
    assign _8993 = _1062 == _4384;
    assign _8994 = _1059 & _8993;
    assign _8998 = _8994 ? _1029 : _8997;
    assign _9000 = _1047 ? _1055 : _8998;
    assign _886 = _9000;
    always @(posedge _1038) begin
        if (_1036)
            _8997 <= _1055;
        else
            _8997 <= _886;
    end
    assign _9002 = _1062 == _4393;
    assign _9003 = _1059 & _9002;
    assign _9007 = _9003 ? _1029 : _9006;
    assign _9009 = _1047 ? _1055 : _9007;
    assign _887 = _9009;
    always @(posedge _1038) begin
        if (_1036)
            _9006 <= _1055;
        else
            _9006 <= _887;
    end
    assign _9011 = _1062 == _4402;
    assign _9012 = _1059 & _9011;
    assign _9016 = _9012 ? _1029 : _9015;
    assign _9018 = _1047 ? _1055 : _9016;
    assign _888 = _9018;
    always @(posedge _1038) begin
        if (_1036)
            _9015 <= _1055;
        else
            _9015 <= _888;
    end
    assign _9020 = _1062 == _4411;
    assign _9021 = _1059 & _9020;
    assign _9025 = _9021 ? _1029 : _9024;
    assign _9027 = _1047 ? _1055 : _9025;
    assign _889 = _9027;
    always @(posedge _1038) begin
        if (_1036)
            _9024 <= _1055;
        else
            _9024 <= _889;
    end
    assign _9029 = _1062 == _4420;
    assign _9030 = _1059 & _9029;
    assign _9034 = _9030 ? _1029 : _9033;
    assign _9036 = _1047 ? _1055 : _9034;
    assign _890 = _9036;
    always @(posedge _1038) begin
        if (_1036)
            _9033 <= _1055;
        else
            _9033 <= _890;
    end
    assign _9038 = _1062 == _4429;
    assign _9039 = _1059 & _9038;
    assign _9043 = _9039 ? _1029 : _9042;
    assign _9045 = _1047 ? _1055 : _9043;
    assign _891 = _9045;
    always @(posedge _1038) begin
        if (_1036)
            _9042 <= _1055;
        else
            _9042 <= _891;
    end
    assign _9047 = _1062 == _4438;
    assign _9048 = _1059 & _9047;
    assign _9052 = _9048 ? _1029 : _9051;
    assign _9054 = _1047 ? _1055 : _9052;
    assign _892 = _9054;
    always @(posedge _1038) begin
        if (_1036)
            _9051 <= _1055;
        else
            _9051 <= _892;
    end
    assign _9056 = _1062 == _4447;
    assign _9057 = _1059 & _9056;
    assign _9061 = _9057 ? _1029 : _9060;
    assign _9063 = _1047 ? _1055 : _9061;
    assign _893 = _9063;
    always @(posedge _1038) begin
        if (_1036)
            _9060 <= _1055;
        else
            _9060 <= _893;
    end
    assign _9065 = _1062 == _4456;
    assign _9066 = _1059 & _9065;
    assign _9070 = _9066 ? _1029 : _9069;
    assign _9072 = _1047 ? _1055 : _9070;
    assign _894 = _9072;
    always @(posedge _1038) begin
        if (_1036)
            _9069 <= _1055;
        else
            _9069 <= _894;
    end
    assign _9074 = _1062 == _4465;
    assign _9075 = _1059 & _9074;
    assign _9079 = _9075 ? _1029 : _9078;
    assign _9081 = _1047 ? _1055 : _9079;
    assign _895 = _9081;
    always @(posedge _1038) begin
        if (_1036)
            _9078 <= _1055;
        else
            _9078 <= _895;
    end
    assign _9083 = _1062 == _4474;
    assign _9084 = _1059 & _9083;
    assign _9088 = _9084 ? _1029 : _9087;
    assign _9090 = _1047 ? _1055 : _9088;
    assign _896 = _9090;
    always @(posedge _1038) begin
        if (_1036)
            _9087 <= _1055;
        else
            _9087 <= _896;
    end
    assign _9092 = _1062 == _4483;
    assign _9093 = _1059 & _9092;
    assign _9097 = _9093 ? _1029 : _9096;
    assign _9099 = _1047 ? _1055 : _9097;
    assign _897 = _9099;
    always @(posedge _1038) begin
        if (_1036)
            _9096 <= _1055;
        else
            _9096 <= _897;
    end
    assign _9101 = _1062 == _4492;
    assign _9102 = _1059 & _9101;
    assign _9106 = _9102 ? _1029 : _9105;
    assign _9108 = _1047 ? _1055 : _9106;
    assign _898 = _9108;
    always @(posedge _1038) begin
        if (_1036)
            _9105 <= _1055;
        else
            _9105 <= _898;
    end
    assign _9110 = _1062 == _4501;
    assign _9111 = _1059 & _9110;
    assign _9115 = _9111 ? _1029 : _9114;
    assign _9117 = _1047 ? _1055 : _9115;
    assign _899 = _9117;
    always @(posedge _1038) begin
        if (_1036)
            _9114 <= _1055;
        else
            _9114 <= _899;
    end
    assign _9119 = _1062 == _4510;
    assign _9120 = _1059 & _9119;
    assign _9124 = _9120 ? _1029 : _9123;
    assign _9126 = _1047 ? _1055 : _9124;
    assign _900 = _9126;
    always @(posedge _1038) begin
        if (_1036)
            _9123 <= _1055;
        else
            _9123 <= _900;
    end
    assign _9128 = _1062 == _4519;
    assign _9129 = _1059 & _9128;
    assign _9133 = _9129 ? _1029 : _9132;
    assign _9135 = _1047 ? _1055 : _9133;
    assign _901 = _9135;
    always @(posedge _1038) begin
        if (_1036)
            _9132 <= _1055;
        else
            _9132 <= _901;
    end
    assign _9137 = _1062 == _4528;
    assign _9138 = _1059 & _9137;
    assign _9142 = _9138 ? _1029 : _9141;
    assign _9144 = _1047 ? _1055 : _9142;
    assign _902 = _9144;
    always @(posedge _1038) begin
        if (_1036)
            _9141 <= _1055;
        else
            _9141 <= _902;
    end
    assign _9146 = _1062 == _4537;
    assign _9147 = _1059 & _9146;
    assign _9151 = _9147 ? _1029 : _9150;
    assign _9153 = _1047 ? _1055 : _9151;
    assign _903 = _9153;
    always @(posedge _1038) begin
        if (_1036)
            _9150 <= _1055;
        else
            _9150 <= _903;
    end
    assign _9155 = _1062 == _4546;
    assign _9156 = _1059 & _9155;
    assign _9160 = _9156 ? _1029 : _9159;
    assign _9162 = _1047 ? _1055 : _9160;
    assign _904 = _9162;
    always @(posedge _1038) begin
        if (_1036)
            _9159 <= _1055;
        else
            _9159 <= _904;
    end
    assign _9164 = _1062 == _4555;
    assign _9165 = _1059 & _9164;
    assign _9169 = _9165 ? _1029 : _9168;
    assign _9171 = _1047 ? _1055 : _9169;
    assign _905 = _9171;
    always @(posedge _1038) begin
        if (_1036)
            _9168 <= _1055;
        else
            _9168 <= _905;
    end
    assign _9173 = _1062 == _4564;
    assign _9174 = _1059 & _9173;
    assign _9178 = _9174 ? _1029 : _9177;
    assign _9180 = _1047 ? _1055 : _9178;
    assign _906 = _9180;
    always @(posedge _1038) begin
        if (_1036)
            _9177 <= _1055;
        else
            _9177 <= _906;
    end
    assign _9182 = _1062 == _4573;
    assign _9183 = _1059 & _9182;
    assign _9187 = _9183 ? _1029 : _9186;
    assign _9189 = _1047 ? _1055 : _9187;
    assign _907 = _9189;
    always @(posedge _1038) begin
        if (_1036)
            _9186 <= _1055;
        else
            _9186 <= _907;
    end
    assign _9191 = _1062 == _4582;
    assign _9192 = _1059 & _9191;
    assign _9196 = _9192 ? _1029 : _9195;
    assign _9198 = _1047 ? _1055 : _9196;
    assign _908 = _9198;
    always @(posedge _1038) begin
        if (_1036)
            _9195 <= _1055;
        else
            _9195 <= _908;
    end
    assign _9200 = _1062 == _4591;
    assign _9201 = _1059 & _9200;
    assign _9205 = _9201 ? _1029 : _9204;
    assign _9207 = _1047 ? _1055 : _9205;
    assign _909 = _9207;
    always @(posedge _1038) begin
        if (_1036)
            _9204 <= _1055;
        else
            _9204 <= _909;
    end
    assign _9209 = _1062 == _4600;
    assign _9210 = _1059 & _9209;
    assign _9214 = _9210 ? _1029 : _9213;
    assign _9216 = _1047 ? _1055 : _9214;
    assign _910 = _9216;
    always @(posedge _1038) begin
        if (_1036)
            _9213 <= _1055;
        else
            _9213 <= _910;
    end
    assign _9218 = _1062 == _4609;
    assign _9219 = _1059 & _9218;
    assign _9223 = _9219 ? _1029 : _9222;
    assign _9225 = _1047 ? _1055 : _9223;
    assign _911 = _9225;
    always @(posedge _1038) begin
        if (_1036)
            _9222 <= _1055;
        else
            _9222 <= _911;
    end
    assign _9227 = _1062 == _4618;
    assign _9228 = _1059 & _9227;
    assign _9232 = _9228 ? _1029 : _9231;
    assign _9234 = _1047 ? _1055 : _9232;
    assign _912 = _9234;
    always @(posedge _1038) begin
        if (_1036)
            _9231 <= _1055;
        else
            _9231 <= _912;
    end
    assign _9236 = _1062 == _4627;
    assign _9237 = _1059 & _9236;
    assign _9241 = _9237 ? _1029 : _9240;
    assign _9243 = _1047 ? _1055 : _9241;
    assign _913 = _9243;
    always @(posedge _1038) begin
        if (_1036)
            _9240 <= _1055;
        else
            _9240 <= _913;
    end
    assign _9245 = _1062 == _4636;
    assign _9246 = _1059 & _9245;
    assign _9250 = _9246 ? _1029 : _9249;
    assign _9252 = _1047 ? _1055 : _9250;
    assign _914 = _9252;
    always @(posedge _1038) begin
        if (_1036)
            _9249 <= _1055;
        else
            _9249 <= _914;
    end
    assign _9254 = _1062 == _4645;
    assign _9255 = _1059 & _9254;
    assign _9259 = _9255 ? _1029 : _9258;
    assign _9261 = _1047 ? _1055 : _9259;
    assign _915 = _9261;
    always @(posedge _1038) begin
        if (_1036)
            _9258 <= _1055;
        else
            _9258 <= _915;
    end
    assign _9263 = _1062 == _4654;
    assign _9264 = _1059 & _9263;
    assign _9268 = _9264 ? _1029 : _9267;
    assign _9270 = _1047 ? _1055 : _9268;
    assign _916 = _9270;
    always @(posedge _1038) begin
        if (_1036)
            _9267 <= _1055;
        else
            _9267 <= _916;
    end
    assign _9272 = _1062 == _4663;
    assign _9273 = _1059 & _9272;
    assign _9277 = _9273 ? _1029 : _9276;
    assign _9279 = _1047 ? _1055 : _9277;
    assign _917 = _9279;
    always @(posedge _1038) begin
        if (_1036)
            _9276 <= _1055;
        else
            _9276 <= _917;
    end
    assign _9281 = _1062 == _4672;
    assign _9282 = _1059 & _9281;
    assign _9286 = _9282 ? _1029 : _9285;
    assign _9288 = _1047 ? _1055 : _9286;
    assign _918 = _9288;
    always @(posedge _1038) begin
        if (_1036)
            _9285 <= _1055;
        else
            _9285 <= _918;
    end
    assign _9290 = _1062 == _4681;
    assign _9291 = _1059 & _9290;
    assign _9295 = _9291 ? _1029 : _9294;
    assign _9297 = _1047 ? _1055 : _9295;
    assign _919 = _9297;
    always @(posedge _1038) begin
        if (_1036)
            _9294 <= _1055;
        else
            _9294 <= _919;
    end
    assign _9299 = _1062 == _4690;
    assign _9300 = _1059 & _9299;
    assign _9304 = _9300 ? _1029 : _9303;
    assign _9306 = _1047 ? _1055 : _9304;
    assign _920 = _9306;
    always @(posedge _1038) begin
        if (_1036)
            _9303 <= _1055;
        else
            _9303 <= _920;
    end
    assign _9308 = _1062 == _4699;
    assign _9309 = _1059 & _9308;
    assign _9313 = _9309 ? _1029 : _9312;
    assign _9315 = _1047 ? _1055 : _9313;
    assign _921 = _9315;
    always @(posedge _1038) begin
        if (_1036)
            _9312 <= _1055;
        else
            _9312 <= _921;
    end
    assign _9317 = _1062 == _4708;
    assign _9318 = _1059 & _9317;
    assign _9322 = _9318 ? _1029 : _9321;
    assign _9324 = _1047 ? _1055 : _9322;
    assign _922 = _9324;
    always @(posedge _1038) begin
        if (_1036)
            _9321 <= _1055;
        else
            _9321 <= _922;
    end
    assign _9326 = _1062 == _4717;
    assign _9327 = _1059 & _9326;
    assign _9331 = _9327 ? _1029 : _9330;
    assign _9333 = _1047 ? _1055 : _9331;
    assign _923 = _9333;
    always @(posedge _1038) begin
        if (_1036)
            _9330 <= _1055;
        else
            _9330 <= _923;
    end
    assign _9335 = _1062 == _4726;
    assign _9336 = _1059 & _9335;
    assign _9340 = _9336 ? _1029 : _9339;
    assign _9342 = _1047 ? _1055 : _9340;
    assign _924 = _9342;
    always @(posedge _1038) begin
        if (_1036)
            _9339 <= _1055;
        else
            _9339 <= _924;
    end
    assign _9344 = _1062 == _4735;
    assign _9345 = _1059 & _9344;
    assign _9349 = _9345 ? _1029 : _9348;
    assign _9351 = _1047 ? _1055 : _9349;
    assign _925 = _9351;
    always @(posedge _1038) begin
        if (_1036)
            _9348 <= _1055;
        else
            _9348 <= _925;
    end
    assign _9353 = _1062 == _4744;
    assign _9354 = _1059 & _9353;
    assign _9358 = _9354 ? _1029 : _9357;
    assign _9360 = _1047 ? _1055 : _9358;
    assign _926 = _9360;
    always @(posedge _1038) begin
        if (_1036)
            _9357 <= _1055;
        else
            _9357 <= _926;
    end
    assign _9362 = _1062 == _4753;
    assign _9363 = _1059 & _9362;
    assign _9367 = _9363 ? _1029 : _9366;
    assign _9369 = _1047 ? _1055 : _9367;
    assign _927 = _9369;
    always @(posedge _1038) begin
        if (_1036)
            _9366 <= _1055;
        else
            _9366 <= _927;
    end
    assign _9371 = _1062 == _4762;
    assign _9372 = _1059 & _9371;
    assign _9376 = _9372 ? _1029 : _9375;
    assign _9378 = _1047 ? _1055 : _9376;
    assign _928 = _9378;
    always @(posedge _1038) begin
        if (_1036)
            _9375 <= _1055;
        else
            _9375 <= _928;
    end
    assign _9380 = _1062 == _4771;
    assign _9381 = _1059 & _9380;
    assign _9385 = _9381 ? _1029 : _9384;
    assign _9387 = _1047 ? _1055 : _9385;
    assign _929 = _9387;
    always @(posedge _1038) begin
        if (_1036)
            _9384 <= _1055;
        else
            _9384 <= _929;
    end
    assign _9389 = _1062 == _4780;
    assign _9390 = _1059 & _9389;
    assign _9394 = _9390 ? _1029 : _9393;
    assign _9396 = _1047 ? _1055 : _9394;
    assign _930 = _9396;
    always @(posedge _1038) begin
        if (_1036)
            _9393 <= _1055;
        else
            _9393 <= _930;
    end
    assign _9398 = _1062 == _4789;
    assign _9399 = _1059 & _9398;
    assign _9403 = _9399 ? _1029 : _9402;
    assign _9405 = _1047 ? _1055 : _9403;
    assign _931 = _9405;
    always @(posedge _1038) begin
        if (_1036)
            _9402 <= _1055;
        else
            _9402 <= _931;
    end
    assign _9407 = _1062 == _4798;
    assign _9408 = _1059 & _9407;
    assign _9412 = _9408 ? _1029 : _9411;
    assign _9414 = _1047 ? _1055 : _9412;
    assign _932 = _9414;
    always @(posedge _1038) begin
        if (_1036)
            _9411 <= _1055;
        else
            _9411 <= _932;
    end
    assign _9416 = _1062 == _4807;
    assign _9417 = _1059 & _9416;
    assign _9421 = _9417 ? _1029 : _9420;
    assign _9423 = _1047 ? _1055 : _9421;
    assign _933 = _9423;
    always @(posedge _1038) begin
        if (_1036)
            _9420 <= _1055;
        else
            _9420 <= _933;
    end
    assign _9425 = _1062 == _4816;
    assign _9426 = _1059 & _9425;
    assign _9430 = _9426 ? _1029 : _9429;
    assign _9432 = _1047 ? _1055 : _9430;
    assign _934 = _9432;
    always @(posedge _1038) begin
        if (_1036)
            _9429 <= _1055;
        else
            _9429 <= _934;
    end
    assign _9434 = _1062 == _4825;
    assign _9435 = _1059 & _9434;
    assign _9439 = _9435 ? _1029 : _9438;
    assign _9441 = _1047 ? _1055 : _9439;
    assign _935 = _9441;
    always @(posedge _1038) begin
        if (_1036)
            _9438 <= _1055;
        else
            _9438 <= _935;
    end
    assign _9443 = _1062 == _4834;
    assign _9444 = _1059 & _9443;
    assign _9448 = _9444 ? _1029 : _9447;
    assign _9450 = _1047 ? _1055 : _9448;
    assign _936 = _9450;
    always @(posedge _1038) begin
        if (_1036)
            _9447 <= _1055;
        else
            _9447 <= _936;
    end
    assign _9452 = _1062 == _4843;
    assign _9453 = _1059 & _9452;
    assign _9457 = _9453 ? _1029 : _9456;
    assign _9459 = _1047 ? _1055 : _9457;
    assign _937 = _9459;
    always @(posedge _1038) begin
        if (_1036)
            _9456 <= _1055;
        else
            _9456 <= _937;
    end
    assign _9461 = _1062 == _4852;
    assign _9462 = _1059 & _9461;
    assign _9466 = _9462 ? _1029 : _9465;
    assign _9468 = _1047 ? _1055 : _9466;
    assign _938 = _9468;
    always @(posedge _1038) begin
        if (_1036)
            _9465 <= _1055;
        else
            _9465 <= _938;
    end
    assign _9470 = _1062 == _4861;
    assign _9471 = _1059 & _9470;
    assign _9475 = _9471 ? _1029 : _9474;
    assign _9477 = _1047 ? _1055 : _9475;
    assign _939 = _9477;
    always @(posedge _1038) begin
        if (_1036)
            _9474 <= _1055;
        else
            _9474 <= _939;
    end
    assign _9479 = _1062 == _4870;
    assign _9480 = _1059 & _9479;
    assign _9484 = _9480 ? _1029 : _9483;
    assign _9486 = _1047 ? _1055 : _9484;
    assign _940 = _9486;
    always @(posedge _1038) begin
        if (_1036)
            _9483 <= _1055;
        else
            _9483 <= _940;
    end
    assign _9488 = _1062 == _4879;
    assign _9489 = _1059 & _9488;
    assign _9493 = _9489 ? _1029 : _9492;
    assign _9495 = _1047 ? _1055 : _9493;
    assign _941 = _9495;
    always @(posedge _1038) begin
        if (_1036)
            _9492 <= _1055;
        else
            _9492 <= _941;
    end
    assign _9497 = _1062 == _4888;
    assign _9498 = _1059 & _9497;
    assign _9502 = _9498 ? _1029 : _9501;
    assign _9504 = _1047 ? _1055 : _9502;
    assign _942 = _9504;
    always @(posedge _1038) begin
        if (_1036)
            _9501 <= _1055;
        else
            _9501 <= _942;
    end
    assign _9506 = _1062 == _4897;
    assign _9507 = _1059 & _9506;
    assign _9511 = _9507 ? _1029 : _9510;
    assign _9513 = _1047 ? _1055 : _9511;
    assign _943 = _9513;
    always @(posedge _1038) begin
        if (_1036)
            _9510 <= _1055;
        else
            _9510 <= _943;
    end
    assign _9515 = _1062 == _4906;
    assign _9516 = _1059 & _9515;
    assign _9520 = _9516 ? _1029 : _9519;
    assign _9522 = _1047 ? _1055 : _9520;
    assign _944 = _9522;
    always @(posedge _1038) begin
        if (_1036)
            _9519 <= _1055;
        else
            _9519 <= _944;
    end
    assign _9524 = _1062 == _4915;
    assign _9525 = _1059 & _9524;
    assign _9529 = _9525 ? _1029 : _9528;
    assign _9531 = _1047 ? _1055 : _9529;
    assign _945 = _9531;
    always @(posedge _1038) begin
        if (_1036)
            _9528 <= _1055;
        else
            _9528 <= _945;
    end
    assign _9533 = _1062 == _4924;
    assign _9534 = _1059 & _9533;
    assign _9538 = _9534 ? _1029 : _9537;
    assign _9540 = _1047 ? _1055 : _9538;
    assign _946 = _9540;
    always @(posedge _1038) begin
        if (_1036)
            _9537 <= _1055;
        else
            _9537 <= _946;
    end
    assign _9542 = _1062 == _4933;
    assign _9543 = _1059 & _9542;
    assign _9547 = _9543 ? _1029 : _9546;
    assign _9549 = _1047 ? _1055 : _9547;
    assign _947 = _9549;
    always @(posedge _1038) begin
        if (_1036)
            _9546 <= _1055;
        else
            _9546 <= _947;
    end
    assign _9551 = _1062 == _4942;
    assign _9552 = _1059 & _9551;
    assign _9556 = _9552 ? _1029 : _9555;
    assign _9558 = _1047 ? _1055 : _9556;
    assign _948 = _9558;
    always @(posedge _1038) begin
        if (_1036)
            _9555 <= _1055;
        else
            _9555 <= _948;
    end
    assign _9560 = _1062 == _4951;
    assign _9561 = _1059 & _9560;
    assign _9565 = _9561 ? _1029 : _9564;
    assign _9567 = _1047 ? _1055 : _9565;
    assign _949 = _9567;
    always @(posedge _1038) begin
        if (_1036)
            _9564 <= _1055;
        else
            _9564 <= _949;
    end
    assign _9569 = _1062 == _4960;
    assign _9570 = _1059 & _9569;
    assign _9574 = _9570 ? _1029 : _9573;
    assign _9576 = _1047 ? _1055 : _9574;
    assign _950 = _9576;
    always @(posedge _1038) begin
        if (_1036)
            _9573 <= _1055;
        else
            _9573 <= _950;
    end
    assign _9578 = _1062 == _4969;
    assign _9579 = _1059 & _9578;
    assign _9583 = _9579 ? _1029 : _9582;
    assign _9585 = _1047 ? _1055 : _9583;
    assign _951 = _9585;
    always @(posedge _1038) begin
        if (_1036)
            _9582 <= _1055;
        else
            _9582 <= _951;
    end
    assign _9587 = _1062 == _4978;
    assign _9588 = _1059 & _9587;
    assign _9592 = _9588 ? _1029 : _9591;
    assign _9594 = _1047 ? _1055 : _9592;
    assign _952 = _9594;
    always @(posedge _1038) begin
        if (_1036)
            _9591 <= _1055;
        else
            _9591 <= _952;
    end
    assign _9596 = _1062 == _4987;
    assign _9597 = _1059 & _9596;
    assign _9601 = _9597 ? _1029 : _9600;
    assign _9603 = _1047 ? _1055 : _9601;
    assign _953 = _9603;
    always @(posedge _1038) begin
        if (_1036)
            _9600 <= _1055;
        else
            _9600 <= _953;
    end
    assign _9605 = _1062 == _4996;
    assign _9606 = _1059 & _9605;
    assign _9610 = _9606 ? _1029 : _9609;
    assign _9612 = _1047 ? _1055 : _9610;
    assign _954 = _9612;
    always @(posedge _1038) begin
        if (_1036)
            _9609 <= _1055;
        else
            _9609 <= _954;
    end
    assign _9614 = _1062 == _5005;
    assign _9615 = _1059 & _9614;
    assign _9619 = _9615 ? _1029 : _9618;
    assign _9621 = _1047 ? _1055 : _9619;
    assign _955 = _9621;
    always @(posedge _1038) begin
        if (_1036)
            _9618 <= _1055;
        else
            _9618 <= _955;
    end
    assign _9623 = _1062 == _5014;
    assign _9624 = _1059 & _9623;
    assign _9628 = _9624 ? _1029 : _9627;
    assign _9630 = _1047 ? _1055 : _9628;
    assign _956 = _9630;
    always @(posedge _1038) begin
        if (_1036)
            _9627 <= _1055;
        else
            _9627 <= _956;
    end
    assign _9632 = _1062 == _5023;
    assign _9633 = _1059 & _9632;
    assign _9637 = _9633 ? _1029 : _9636;
    assign _9639 = _1047 ? _1055 : _9637;
    assign _957 = _9639;
    always @(posedge _1038) begin
        if (_1036)
            _9636 <= _1055;
        else
            _9636 <= _957;
    end
    assign _9641 = _1062 == _5032;
    assign _9642 = _1059 & _9641;
    assign _9646 = _9642 ? _1029 : _9645;
    assign _9648 = _1047 ? _1055 : _9646;
    assign _958 = _9648;
    always @(posedge _1038) begin
        if (_1036)
            _9645 <= _1055;
        else
            _9645 <= _958;
    end
    assign _9650 = _1062 == _5041;
    assign _9651 = _1059 & _9650;
    assign _9655 = _9651 ? _1029 : _9654;
    assign _9657 = _1047 ? _1055 : _9655;
    assign _959 = _9657;
    always @(posedge _1038) begin
        if (_1036)
            _9654 <= _1055;
        else
            _9654 <= _959;
    end
    assign _9659 = _1062 == _5050;
    assign _9660 = _1059 & _9659;
    assign _9664 = _9660 ? _1029 : _9663;
    assign _9666 = _1047 ? _1055 : _9664;
    assign _960 = _9666;
    always @(posedge _1038) begin
        if (_1036)
            _9663 <= _1055;
        else
            _9663 <= _960;
    end
    assign _9668 = _1062 == _5059;
    assign _9669 = _1059 & _9668;
    assign _9673 = _9669 ? _1029 : _9672;
    assign _9675 = _1047 ? _1055 : _9673;
    assign _961 = _9675;
    always @(posedge _1038) begin
        if (_1036)
            _9672 <= _1055;
        else
            _9672 <= _961;
    end
    assign _9677 = _1062 == _5068;
    assign _9678 = _1059 & _9677;
    assign _9682 = _9678 ? _1029 : _9681;
    assign _9684 = _1047 ? _1055 : _9682;
    assign _962 = _9684;
    always @(posedge _1038) begin
        if (_1036)
            _9681 <= _1055;
        else
            _9681 <= _962;
    end
    assign _9686 = _1062 == _5077;
    assign _9687 = _1059 & _9686;
    assign _9691 = _9687 ? _1029 : _9690;
    assign _9693 = _1047 ? _1055 : _9691;
    assign _963 = _9693;
    always @(posedge _1038) begin
        if (_1036)
            _9690 <= _1055;
        else
            _9690 <= _963;
    end
    assign _9695 = _1062 == _5086;
    assign _9696 = _1059 & _9695;
    assign _9700 = _9696 ? _1029 : _9699;
    assign _9702 = _1047 ? _1055 : _9700;
    assign _964 = _9702;
    always @(posedge _1038) begin
        if (_1036)
            _9699 <= _1055;
        else
            _9699 <= _964;
    end
    assign _9704 = _1062 == _5095;
    assign _9705 = _1059 & _9704;
    assign _9709 = _9705 ? _1029 : _9708;
    assign _9711 = _1047 ? _1055 : _9709;
    assign _965 = _9711;
    always @(posedge _1038) begin
        if (_1036)
            _9708 <= _1055;
        else
            _9708 <= _965;
    end
    assign _9713 = _1062 == _5104;
    assign _9714 = _1059 & _9713;
    assign _9718 = _9714 ? _1029 : _9717;
    assign _9720 = _1047 ? _1055 : _9718;
    assign _966 = _9720;
    always @(posedge _1038) begin
        if (_1036)
            _9717 <= _1055;
        else
            _9717 <= _966;
    end
    assign _9722 = _1062 == _5113;
    assign _9723 = _1059 & _9722;
    assign _9727 = _9723 ? _1029 : _9726;
    assign _9729 = _1047 ? _1055 : _9727;
    assign _967 = _9729;
    always @(posedge _1038) begin
        if (_1036)
            _9726 <= _1055;
        else
            _9726 <= _967;
    end
    assign _9731 = _1062 == _5122;
    assign _9732 = _1059 & _9731;
    assign _9736 = _9732 ? _1029 : _9735;
    assign _9738 = _1047 ? _1055 : _9736;
    assign _968 = _9738;
    always @(posedge _1038) begin
        if (_1036)
            _9735 <= _1055;
        else
            _9735 <= _968;
    end
    assign _9740 = _1062 == _5131;
    assign _9741 = _1059 & _9740;
    assign _9745 = _9741 ? _1029 : _9744;
    assign _9747 = _1047 ? _1055 : _9745;
    assign _969 = _9747;
    always @(posedge _1038) begin
        if (_1036)
            _9744 <= _1055;
        else
            _9744 <= _969;
    end
    assign _9749 = _1062 == _5140;
    assign _9750 = _1059 & _9749;
    assign _9754 = _9750 ? _1029 : _9753;
    assign _9756 = _1047 ? _1055 : _9754;
    assign _970 = _9756;
    always @(posedge _1038) begin
        if (_1036)
            _9753 <= _1055;
        else
            _9753 <= _970;
    end
    assign _9758 = _1062 == _5149;
    assign _9759 = _1059 & _9758;
    assign _9763 = _9759 ? _1029 : _9762;
    assign _9765 = _1047 ? _1055 : _9763;
    assign _971 = _9765;
    always @(posedge _1038) begin
        if (_1036)
            _9762 <= _1055;
        else
            _9762 <= _971;
    end
    assign _9767 = _1062 == _5158;
    assign _9768 = _1059 & _9767;
    assign _9772 = _9768 ? _1029 : _9771;
    assign _9774 = _1047 ? _1055 : _9772;
    assign _972 = _9774;
    always @(posedge _1038) begin
        if (_1036)
            _9771 <= _1055;
        else
            _9771 <= _972;
    end
    assign _9776 = _1062 == _5167;
    assign _9777 = _1059 & _9776;
    assign _9781 = _9777 ? _1029 : _9780;
    assign _9783 = _1047 ? _1055 : _9781;
    assign _973 = _9783;
    always @(posedge _1038) begin
        if (_1036)
            _9780 <= _1055;
        else
            _9780 <= _973;
    end
    assign _9785 = _1062 == _5176;
    assign _9786 = _1059 & _9785;
    assign _9790 = _9786 ? _1029 : _9789;
    assign _9792 = _1047 ? _1055 : _9790;
    assign _974 = _9792;
    always @(posedge _1038) begin
        if (_1036)
            _9789 <= _1055;
        else
            _9789 <= _974;
    end
    assign _9794 = _1062 == _5185;
    assign _9795 = _1059 & _9794;
    assign _9799 = _9795 ? _1029 : _9798;
    assign _9801 = _1047 ? _1055 : _9799;
    assign _975 = _9801;
    always @(posedge _1038) begin
        if (_1036)
            _9798 <= _1055;
        else
            _9798 <= _975;
    end
    assign _9803 = _1062 == _5194;
    assign _9804 = _1059 & _9803;
    assign _9808 = _9804 ? _1029 : _9807;
    assign _9810 = _1047 ? _1055 : _9808;
    assign _976 = _9810;
    always @(posedge _1038) begin
        if (_1036)
            _9807 <= _1055;
        else
            _9807 <= _976;
    end
    assign _9812 = _1062 == _5203;
    assign _9813 = _1059 & _9812;
    assign _9817 = _9813 ? _1029 : _9816;
    assign _9819 = _1047 ? _1055 : _9817;
    assign _977 = _9819;
    always @(posedge _1038) begin
        if (_1036)
            _9816 <= _1055;
        else
            _9816 <= _977;
    end
    assign _9821 = _1062 == _5212;
    assign _9822 = _1059 & _9821;
    assign _9826 = _9822 ? _1029 : _9825;
    assign _9828 = _1047 ? _1055 : _9826;
    assign _978 = _9828;
    always @(posedge _1038) begin
        if (_1036)
            _9825 <= _1055;
        else
            _9825 <= _978;
    end
    assign _9830 = _1062 == _5221;
    assign _9831 = _1059 & _9830;
    assign _9835 = _9831 ? _1029 : _9834;
    assign _9837 = _1047 ? _1055 : _9835;
    assign _979 = _9837;
    always @(posedge _1038) begin
        if (_1036)
            _9834 <= _1055;
        else
            _9834 <= _979;
    end
    assign _9839 = _1062 == _5230;
    assign _9840 = _1059 & _9839;
    assign _9844 = _9840 ? _1029 : _9843;
    assign _9846 = _1047 ? _1055 : _9844;
    assign _980 = _9846;
    always @(posedge _1038) begin
        if (_1036)
            _9843 <= _1055;
        else
            _9843 <= _980;
    end
    assign _9848 = _1062 == _5239;
    assign _9849 = _1059 & _9848;
    assign _9853 = _9849 ? _1029 : _9852;
    assign _9855 = _1047 ? _1055 : _9853;
    assign _981 = _9855;
    always @(posedge _1038) begin
        if (_1036)
            _9852 <= _1055;
        else
            _9852 <= _981;
    end
    assign _9857 = _1062 == _5248;
    assign _9858 = _1059 & _9857;
    assign _9862 = _9858 ? _1029 : _9861;
    assign _9864 = _1047 ? _1055 : _9862;
    assign _982 = _9864;
    always @(posedge _1038) begin
        if (_1036)
            _9861 <= _1055;
        else
            _9861 <= _982;
    end
    assign _9866 = _1062 == _5257;
    assign _9867 = _1059 & _9866;
    assign _9871 = _9867 ? _1029 : _9870;
    assign _9873 = _1047 ? _1055 : _9871;
    assign _983 = _9873;
    always @(posedge _1038) begin
        if (_1036)
            _9870 <= _1055;
        else
            _9870 <= _983;
    end
    assign _9875 = _1062 == _5266;
    assign _9876 = _1059 & _9875;
    assign _9880 = _9876 ? _1029 : _9879;
    assign _9882 = _1047 ? _1055 : _9880;
    assign _984 = _9882;
    always @(posedge _1038) begin
        if (_1036)
            _9879 <= _1055;
        else
            _9879 <= _984;
    end
    assign _9884 = _1062 == _5275;
    assign _9885 = _1059 & _9884;
    assign _9889 = _9885 ? _1029 : _9888;
    assign _9891 = _1047 ? _1055 : _9889;
    assign _985 = _9891;
    always @(posedge _1038) begin
        if (_1036)
            _9888 <= _1055;
        else
            _9888 <= _985;
    end
    assign _9893 = _1062 == _5284;
    assign _9894 = _1059 & _9893;
    assign _9898 = _9894 ? _1029 : _9897;
    assign _9900 = _1047 ? _1055 : _9898;
    assign _986 = _9900;
    always @(posedge _1038) begin
        if (_1036)
            _9897 <= _1055;
        else
            _9897 <= _986;
    end
    assign _9902 = _1062 == _5293;
    assign _9903 = _1059 & _9902;
    assign _9907 = _9903 ? _1029 : _9906;
    assign _9909 = _1047 ? _1055 : _9907;
    assign _987 = _9909;
    always @(posedge _1038) begin
        if (_1036)
            _9906 <= _1055;
        else
            _9906 <= _987;
    end
    assign _9911 = _1062 == _5302;
    assign _9912 = _1059 & _9911;
    assign _9916 = _9912 ? _1029 : _9915;
    assign _9918 = _1047 ? _1055 : _9916;
    assign _988 = _9918;
    always @(posedge _1038) begin
        if (_1036)
            _9915 <= _1055;
        else
            _9915 <= _988;
    end
    assign _9920 = _1062 == _5311;
    assign _9921 = _1059 & _9920;
    assign _9925 = _9921 ? _1029 : _9924;
    assign _9927 = _1047 ? _1055 : _9925;
    assign _989 = _9927;
    always @(posedge _1038) begin
        if (_1036)
            _9924 <= _1055;
        else
            _9924 <= _989;
    end
    assign _9929 = _1062 == _5320;
    assign _9930 = _1059 & _9929;
    assign _9934 = _9930 ? _1029 : _9933;
    assign _9936 = _1047 ? _1055 : _9934;
    assign _990 = _9936;
    always @(posedge _1038) begin
        if (_1036)
            _9933 <= _1055;
        else
            _9933 <= _990;
    end
    assign _9938 = _1062 == _5329;
    assign _9939 = _1059 & _9938;
    assign _9943 = _9939 ? _1029 : _9942;
    assign _9945 = _1047 ? _1055 : _9943;
    assign _991 = _9945;
    always @(posedge _1038) begin
        if (_1036)
            _9942 <= _1055;
        else
            _9942 <= _991;
    end
    assign _9947 = _1062 == _5338;
    assign _9948 = _1059 & _9947;
    assign _9952 = _9948 ? _1029 : _9951;
    assign _9954 = _1047 ? _1055 : _9952;
    assign _992 = _9954;
    always @(posedge _1038) begin
        if (_1036)
            _9951 <= _1055;
        else
            _9951 <= _992;
    end
    assign _9956 = _1062 == _5347;
    assign _9957 = _1059 & _9956;
    assign _9961 = _9957 ? _1029 : _9960;
    assign _9963 = _1047 ? _1055 : _9961;
    assign _993 = _9963;
    always @(posedge _1038) begin
        if (_1036)
            _9960 <= _1055;
        else
            _9960 <= _993;
    end
    assign _9965 = _1062 == _5356;
    assign _9966 = _1059 & _9965;
    assign _9970 = _9966 ? _1029 : _9969;
    assign _9972 = _1047 ? _1055 : _9970;
    assign _994 = _9972;
    always @(posedge _1038) begin
        if (_1036)
            _9969 <= _1055;
        else
            _9969 <= _994;
    end
    assign _9974 = _1062 == _5365;
    assign _9975 = _1059 & _9974;
    assign _9979 = _9975 ? _1029 : _9978;
    assign _9981 = _1047 ? _1055 : _9979;
    assign _995 = _9981;
    always @(posedge _1038) begin
        if (_1036)
            _9978 <= _1055;
        else
            _9978 <= _995;
    end
    assign _9983 = _1062 == _5374;
    assign _9984 = _1059 & _9983;
    assign _9988 = _9984 ? _1029 : _9987;
    assign _9990 = _1047 ? _1055 : _9988;
    assign _996 = _9990;
    always @(posedge _1038) begin
        if (_1036)
            _9987 <= _1055;
        else
            _9987 <= _996;
    end
    assign _9992 = _1062 == _5383;
    assign _9993 = _1059 & _9992;
    assign _9997 = _9993 ? _1029 : _9996;
    assign _9999 = _1047 ? _1055 : _9997;
    assign _997 = _9999;
    always @(posedge _1038) begin
        if (_1036)
            _9996 <= _1055;
        else
            _9996 <= _997;
    end
    assign _10001 = _1062 == _5392;
    assign _10002 = _1059 & _10001;
    assign _10006 = _10002 ? _1029 : _10005;
    assign _10008 = _1047 ? _1055 : _10006;
    assign _998 = _10008;
    always @(posedge _1038) begin
        if (_1036)
            _10005 <= _1055;
        else
            _10005 <= _998;
    end
    assign _10010 = _1062 == _5401;
    assign _10011 = _1059 & _10010;
    assign _10015 = _10011 ? _1029 : _10014;
    assign _10017 = _1047 ? _1055 : _10015;
    assign _999 = _10017;
    always @(posedge _1038) begin
        if (_1036)
            _10014 <= _1055;
        else
            _10014 <= _999;
    end
    assign _10019 = _1062 == _5410;
    assign _10020 = _1059 & _10019;
    assign _10024 = _10020 ? _1029 : _10023;
    assign _10026 = _1047 ? _1055 : _10024;
    assign _1000 = _10026;
    always @(posedge _1038) begin
        if (_1036)
            _10023 <= _1055;
        else
            _10023 <= _1000;
    end
    assign _10028 = _1062 == _5419;
    assign _10029 = _1059 & _10028;
    assign _10033 = _10029 ? _1029 : _10032;
    assign _10035 = _1047 ? _1055 : _10033;
    assign _1001 = _10035;
    always @(posedge _1038) begin
        if (_1036)
            _10032 <= _1055;
        else
            _10032 <= _1001;
    end
    assign _10037 = _1062 == _5428;
    assign _10038 = _1059 & _10037;
    assign _10042 = _10038 ? _1029 : _10041;
    assign _10044 = _1047 ? _1055 : _10042;
    assign _1002 = _10044;
    always @(posedge _1038) begin
        if (_1036)
            _10041 <= _1055;
        else
            _10041 <= _1002;
    end
    assign _10046 = _1062 == _5437;
    assign _10047 = _1059 & _10046;
    assign _10051 = _10047 ? _1029 : _10050;
    assign _10053 = _1047 ? _1055 : _10051;
    assign _1003 = _10053;
    always @(posedge _1038) begin
        if (_1036)
            _10050 <= _1055;
        else
            _10050 <= _1003;
    end
    assign _10055 = _1062 == _5446;
    assign _10056 = _1059 & _10055;
    assign _10060 = _10056 ? _1029 : _10059;
    assign _10062 = _1047 ? _1055 : _10060;
    assign _1004 = _10062;
    always @(posedge _1038) begin
        if (_1036)
            _10059 <= _1055;
        else
            _10059 <= _1004;
    end
    assign _10064 = _1062 == _5455;
    assign _10065 = _1059 & _10064;
    assign _10069 = _10065 ? _1029 : _10068;
    assign _10071 = _1047 ? _1055 : _10069;
    assign _1005 = _10071;
    always @(posedge _1038) begin
        if (_1036)
            _10068 <= _1055;
        else
            _10068 <= _1005;
    end
    assign _10073 = _1062 == _5464;
    assign _10074 = _1059 & _10073;
    assign _10078 = _10074 ? _1029 : _10077;
    assign _10080 = _1047 ? _1055 : _10078;
    assign _1006 = _10080;
    always @(posedge _1038) begin
        if (_1036)
            _10077 <= _1055;
        else
            _10077 <= _1006;
    end
    assign _10082 = _1062 == _5473;
    assign _10083 = _1059 & _10082;
    assign _10087 = _10083 ? _1029 : _10086;
    assign _10089 = _1047 ? _1055 : _10087;
    assign _1007 = _10089;
    always @(posedge _1038) begin
        if (_1036)
            _10086 <= _1055;
        else
            _10086 <= _1007;
    end
    assign _10091 = _1062 == _5482;
    assign _10092 = _1059 & _10091;
    assign _10096 = _10092 ? _1029 : _10095;
    assign _10098 = _1047 ? _1055 : _10096;
    assign _1008 = _10098;
    always @(posedge _1038) begin
        if (_1036)
            _10095 <= _1055;
        else
            _10095 <= _1008;
    end
    assign _10100 = _1062 == _5491;
    assign _10101 = _1059 & _10100;
    assign _10105 = _10101 ? _1029 : _10104;
    assign _10107 = _1047 ? _1055 : _10105;
    assign _1009 = _10107;
    always @(posedge _1038) begin
        if (_1036)
            _10104 <= _1055;
        else
            _10104 <= _1009;
    end
    assign _10109 = _1062 == _5500;
    assign _10110 = _1059 & _10109;
    assign _10114 = _10110 ? _1029 : _10113;
    assign _10116 = _1047 ? _1055 : _10114;
    assign _1010 = _10116;
    always @(posedge _1038) begin
        if (_1036)
            _10113 <= _1055;
        else
            _10113 <= _1010;
    end
    assign _10118 = _1062 == _5509;
    assign _10119 = _1059 & _10118;
    assign _10123 = _10119 ? _1029 : _10122;
    assign _10125 = _1047 ? _1055 : _10123;
    assign _1011 = _10125;
    always @(posedge _1038) begin
        if (_1036)
            _10122 <= _1055;
        else
            _10122 <= _1011;
    end
    assign _10127 = _1062 == _5518;
    assign _10128 = _1059 & _10127;
    assign _10132 = _10128 ? _1029 : _10131;
    assign _10134 = _1047 ? _1055 : _10132;
    assign _1012 = _10134;
    always @(posedge _1038) begin
        if (_1036)
            _10131 <= _1055;
        else
            _10131 <= _1012;
    end
    assign _10136 = _1062 == _5527;
    assign _10137 = _1059 & _10136;
    assign _10141 = _10137 ? _1029 : _10140;
    assign _10143 = _1047 ? _1055 : _10141;
    assign _1013 = _10143;
    always @(posedge _1038) begin
        if (_1036)
            _10140 <= _1055;
        else
            _10140 <= _1013;
    end
    assign _10145 = _1062 == _5536;
    assign _10146 = _1059 & _10145;
    assign _10150 = _10146 ? _1029 : _10149;
    assign _10152 = _1047 ? _1055 : _10150;
    assign _1014 = _10152;
    always @(posedge _1038) begin
        if (_1036)
            _10149 <= _1055;
        else
            _10149 <= _1014;
    end
    assign _10154 = _1062 == _5545;
    assign _10155 = _1059 & _10154;
    assign _10159 = _10155 ? _1029 : _10158;
    assign _10161 = _1047 ? _1055 : _10159;
    assign _1015 = _10161;
    always @(posedge _1038) begin
        if (_1036)
            _10158 <= _1055;
        else
            _10158 <= _1015;
    end
    assign _10163 = _1062 == _5554;
    assign _10164 = _1059 & _10163;
    assign _10168 = _10164 ? _1029 : _10167;
    assign _10170 = _1047 ? _1055 : _10168;
    assign _1016 = _10170;
    always @(posedge _1038) begin
        if (_1036)
            _10167 <= _1055;
        else
            _10167 <= _1016;
    end
    assign _10172 = _1062 == _5563;
    assign _10173 = _1059 & _10172;
    assign _10177 = _10173 ? _1029 : _10176;
    assign _10179 = _1047 ? _1055 : _10177;
    assign _1017 = _10179;
    always @(posedge _1038) begin
        if (_1036)
            _10176 <= _1055;
        else
            _10176 <= _1017;
    end
    assign _10181 = _1062 == _5572;
    assign _10182 = _1059 & _10181;
    assign _10186 = _10182 ? _1029 : _10185;
    assign _10188 = _1047 ? _1055 : _10186;
    assign _1018 = _10188;
    always @(posedge _1038) begin
        if (_1036)
            _10185 <= _1055;
        else
            _10185 <= _1018;
    end
    assign _10190 = _1062 == _5581;
    assign _10191 = _1059 & _10190;
    assign _10195 = _10191 ? _1029 : _10194;
    assign _10197 = _1047 ? _1055 : _10195;
    assign _1019 = _10197;
    always @(posedge _1038) begin
        if (_1036)
            _10194 <= _1055;
        else
            _10194 <= _1019;
    end
    assign _10199 = _1062 == _5590;
    assign _10200 = _1059 & _10199;
    assign _10204 = _10200 ? _1029 : _10203;
    assign _10206 = _1047 ? _1055 : _10204;
    assign _1020 = _10206;
    always @(posedge _1038) begin
        if (_1036)
            _10203 <= _1055;
        else
            _10203 <= _1020;
    end
    assign _10208 = _1062 == _5599;
    assign _10209 = _1059 & _10208;
    assign _10213 = _10209 ? _1029 : _10212;
    assign _10215 = _1047 ? _1055 : _10213;
    assign _1021 = _10215;
    always @(posedge _1038) begin
        if (_1036)
            _10212 <= _1055;
        else
            _10212 <= _1021;
    end
    assign _10217 = _1062 == _5608;
    assign _10218 = _1059 & _10217;
    assign _10222 = _10218 ? _1029 : _10221;
    assign _10224 = _1047 ? _1055 : _10222;
    assign _1022 = _10224;
    always @(posedge _1038) begin
        if (_1036)
            _10221 <= _1055;
        else
            _10221 <= _1022;
    end
    assign _10226 = _1062 == _5617;
    assign _10227 = _1059 & _10226;
    assign _10231 = _10227 ? _1029 : _10230;
    assign _10233 = _1047 ? _1055 : _10231;
    assign _1023 = _10233;
    always @(posedge _1038) begin
        if (_1036)
            _10230 <= _1055;
        else
            _10230 <= _1023;
    end
    assign _10235 = _1062 == _5626;
    assign _10236 = _1059 & _10235;
    assign _10240 = _10236 ? _1029 : _10239;
    assign _10242 = _1047 ? _1055 : _10240;
    assign _1024 = _10242;
    always @(posedge _1038) begin
        if (_1036)
            _10239 <= _1055;
        else
            _10239 <= _1024;
    end
    assign _10244 = _1062 == _5635;
    assign _10245 = _1059 & _10244;
    assign _10249 = _10245 ? _1029 : _10248;
    assign _10251 = _1047 ? _1055 : _10249;
    assign _1025 = _10251;
    always @(posedge _1038) begin
        if (_1036)
            _10248 <= _1055;
        else
            _10248 <= _1025;
    end
    assign _10253 = _1062 == _5644;
    assign _10254 = _1059 & _10253;
    assign _10258 = _10254 ? _1029 : _10257;
    assign _10260 = _1047 ? _1055 : _10258;
    assign _1026 = _10260;
    always @(posedge _1038) begin
        if (_1036)
            _10257 <= _1055;
        else
            _10257 <= _1026;
    end
    assign _10262 = _1062 == _5653;
    assign _10263 = _1059 & _10262;
    assign _10267 = _10263 ? _1029 : _10266;
    assign _10269 = _1047 ? _1055 : _10267;
    assign _1027 = _10269;
    always @(posedge _1038) begin
        if (_1036)
            _10266 <= _1055;
        else
            _10266 <= _1027;
    end
    assign _1029 = x;
    assign _10271 = _1062 == _5662;
    assign _10272 = _1059 & _10271;
    assign _10276 = _10272 ? _1029 : _10275;
    assign _10278 = _1047 ? _1055 : _10276;
    assign _1030 = _10278;
    always @(posedge _1038) begin
        if (_1036)
            _10275 <= _1055;
        else
            _10275 <= _1030;
    end
    always @* begin
        case (_10283)
        0:
            _10295 <= _10275;
        1:
            _10295 <= _10266;
        2:
            _10295 <= _10257;
        3:
            _10295 <= _10248;
        4:
            _10295 <= _10239;
        5:
            _10295 <= _10230;
        6:
            _10295 <= _10221;
        7:
            _10295 <= _10212;
        8:
            _10295 <= _10203;
        9:
            _10295 <= _10194;
        10:
            _10295 <= _10185;
        11:
            _10295 <= _10176;
        12:
            _10295 <= _10167;
        13:
            _10295 <= _10158;
        14:
            _10295 <= _10149;
        15:
            _10295 <= _10140;
        16:
            _10295 <= _10131;
        17:
            _10295 <= _10122;
        18:
            _10295 <= _10113;
        19:
            _10295 <= _10104;
        20:
            _10295 <= _10095;
        21:
            _10295 <= _10086;
        22:
            _10295 <= _10077;
        23:
            _10295 <= _10068;
        24:
            _10295 <= _10059;
        25:
            _10295 <= _10050;
        26:
            _10295 <= _10041;
        27:
            _10295 <= _10032;
        28:
            _10295 <= _10023;
        29:
            _10295 <= _10014;
        30:
            _10295 <= _10005;
        31:
            _10295 <= _9996;
        32:
            _10295 <= _9987;
        33:
            _10295 <= _9978;
        34:
            _10295 <= _9969;
        35:
            _10295 <= _9960;
        36:
            _10295 <= _9951;
        37:
            _10295 <= _9942;
        38:
            _10295 <= _9933;
        39:
            _10295 <= _9924;
        40:
            _10295 <= _9915;
        41:
            _10295 <= _9906;
        42:
            _10295 <= _9897;
        43:
            _10295 <= _9888;
        44:
            _10295 <= _9879;
        45:
            _10295 <= _9870;
        46:
            _10295 <= _9861;
        47:
            _10295 <= _9852;
        48:
            _10295 <= _9843;
        49:
            _10295 <= _9834;
        50:
            _10295 <= _9825;
        51:
            _10295 <= _9816;
        52:
            _10295 <= _9807;
        53:
            _10295 <= _9798;
        54:
            _10295 <= _9789;
        55:
            _10295 <= _9780;
        56:
            _10295 <= _9771;
        57:
            _10295 <= _9762;
        58:
            _10295 <= _9753;
        59:
            _10295 <= _9744;
        60:
            _10295 <= _9735;
        61:
            _10295 <= _9726;
        62:
            _10295 <= _9717;
        63:
            _10295 <= _9708;
        64:
            _10295 <= _9699;
        65:
            _10295 <= _9690;
        66:
            _10295 <= _9681;
        67:
            _10295 <= _9672;
        68:
            _10295 <= _9663;
        69:
            _10295 <= _9654;
        70:
            _10295 <= _9645;
        71:
            _10295 <= _9636;
        72:
            _10295 <= _9627;
        73:
            _10295 <= _9618;
        74:
            _10295 <= _9609;
        75:
            _10295 <= _9600;
        76:
            _10295 <= _9591;
        77:
            _10295 <= _9582;
        78:
            _10295 <= _9573;
        79:
            _10295 <= _9564;
        80:
            _10295 <= _9555;
        81:
            _10295 <= _9546;
        82:
            _10295 <= _9537;
        83:
            _10295 <= _9528;
        84:
            _10295 <= _9519;
        85:
            _10295 <= _9510;
        86:
            _10295 <= _9501;
        87:
            _10295 <= _9492;
        88:
            _10295 <= _9483;
        89:
            _10295 <= _9474;
        90:
            _10295 <= _9465;
        91:
            _10295 <= _9456;
        92:
            _10295 <= _9447;
        93:
            _10295 <= _9438;
        94:
            _10295 <= _9429;
        95:
            _10295 <= _9420;
        96:
            _10295 <= _9411;
        97:
            _10295 <= _9402;
        98:
            _10295 <= _9393;
        99:
            _10295 <= _9384;
        100:
            _10295 <= _9375;
        101:
            _10295 <= _9366;
        102:
            _10295 <= _9357;
        103:
            _10295 <= _9348;
        104:
            _10295 <= _9339;
        105:
            _10295 <= _9330;
        106:
            _10295 <= _9321;
        107:
            _10295 <= _9312;
        108:
            _10295 <= _9303;
        109:
            _10295 <= _9294;
        110:
            _10295 <= _9285;
        111:
            _10295 <= _9276;
        112:
            _10295 <= _9267;
        113:
            _10295 <= _9258;
        114:
            _10295 <= _9249;
        115:
            _10295 <= _9240;
        116:
            _10295 <= _9231;
        117:
            _10295 <= _9222;
        118:
            _10295 <= _9213;
        119:
            _10295 <= _9204;
        120:
            _10295 <= _9195;
        121:
            _10295 <= _9186;
        122:
            _10295 <= _9177;
        123:
            _10295 <= _9168;
        124:
            _10295 <= _9159;
        125:
            _10295 <= _9150;
        126:
            _10295 <= _9141;
        127:
            _10295 <= _9132;
        128:
            _10295 <= _9123;
        129:
            _10295 <= _9114;
        130:
            _10295 <= _9105;
        131:
            _10295 <= _9096;
        132:
            _10295 <= _9087;
        133:
            _10295 <= _9078;
        134:
            _10295 <= _9069;
        135:
            _10295 <= _9060;
        136:
            _10295 <= _9051;
        137:
            _10295 <= _9042;
        138:
            _10295 <= _9033;
        139:
            _10295 <= _9024;
        140:
            _10295 <= _9015;
        141:
            _10295 <= _9006;
        142:
            _10295 <= _8997;
        143:
            _10295 <= _8988;
        144:
            _10295 <= _8979;
        145:
            _10295 <= _8970;
        146:
            _10295 <= _8961;
        147:
            _10295 <= _8952;
        148:
            _10295 <= _8943;
        149:
            _10295 <= _8934;
        150:
            _10295 <= _8925;
        151:
            _10295 <= _8916;
        152:
            _10295 <= _8907;
        153:
            _10295 <= _8898;
        154:
            _10295 <= _8889;
        155:
            _10295 <= _8880;
        156:
            _10295 <= _8871;
        157:
            _10295 <= _8862;
        158:
            _10295 <= _8853;
        159:
            _10295 <= _8844;
        160:
            _10295 <= _8835;
        161:
            _10295 <= _8826;
        162:
            _10295 <= _8817;
        163:
            _10295 <= _8808;
        164:
            _10295 <= _8799;
        165:
            _10295 <= _8790;
        166:
            _10295 <= _8781;
        167:
            _10295 <= _8772;
        168:
            _10295 <= _8763;
        169:
            _10295 <= _8754;
        170:
            _10295 <= _8745;
        171:
            _10295 <= _8736;
        172:
            _10295 <= _8727;
        173:
            _10295 <= _8718;
        174:
            _10295 <= _8709;
        175:
            _10295 <= _8700;
        176:
            _10295 <= _8691;
        177:
            _10295 <= _8682;
        178:
            _10295 <= _8673;
        179:
            _10295 <= _8664;
        180:
            _10295 <= _8655;
        181:
            _10295 <= _8646;
        182:
            _10295 <= _8637;
        183:
            _10295 <= _8628;
        184:
            _10295 <= _8619;
        185:
            _10295 <= _8610;
        186:
            _10295 <= _8601;
        187:
            _10295 <= _8592;
        188:
            _10295 <= _8583;
        189:
            _10295 <= _8574;
        190:
            _10295 <= _8565;
        191:
            _10295 <= _8556;
        192:
            _10295 <= _8547;
        193:
            _10295 <= _8538;
        194:
            _10295 <= _8529;
        195:
            _10295 <= _8520;
        196:
            _10295 <= _8511;
        197:
            _10295 <= _8502;
        198:
            _10295 <= _8493;
        199:
            _10295 <= _8484;
        200:
            _10295 <= _8475;
        201:
            _10295 <= _8466;
        202:
            _10295 <= _8457;
        203:
            _10295 <= _8448;
        204:
            _10295 <= _8439;
        205:
            _10295 <= _8430;
        206:
            _10295 <= _8421;
        207:
            _10295 <= _8412;
        208:
            _10295 <= _8403;
        209:
            _10295 <= _8394;
        210:
            _10295 <= _8385;
        211:
            _10295 <= _8376;
        212:
            _10295 <= _8367;
        213:
            _10295 <= _8358;
        214:
            _10295 <= _8349;
        215:
            _10295 <= _8340;
        216:
            _10295 <= _8331;
        217:
            _10295 <= _8322;
        218:
            _10295 <= _8313;
        219:
            _10295 <= _8304;
        220:
            _10295 <= _8295;
        221:
            _10295 <= _8286;
        222:
            _10295 <= _8277;
        223:
            _10295 <= _8268;
        224:
            _10295 <= _8259;
        225:
            _10295 <= _8250;
        226:
            _10295 <= _8241;
        227:
            _10295 <= _8232;
        228:
            _10295 <= _8223;
        229:
            _10295 <= _8214;
        230:
            _10295 <= _8205;
        231:
            _10295 <= _8196;
        232:
            _10295 <= _8187;
        233:
            _10295 <= _8178;
        234:
            _10295 <= _8169;
        235:
            _10295 <= _8160;
        236:
            _10295 <= _8151;
        237:
            _10295 <= _8142;
        238:
            _10295 <= _8133;
        239:
            _10295 <= _8124;
        240:
            _10295 <= _8115;
        241:
            _10295 <= _8106;
        242:
            _10295 <= _8097;
        243:
            _10295 <= _8088;
        244:
            _10295 <= _8079;
        245:
            _10295 <= _8070;
        246:
            _10295 <= _8061;
        247:
            _10295 <= _8052;
        248:
            _10295 <= _8043;
        249:
            _10295 <= _8034;
        250:
            _10295 <= _8025;
        251:
            _10295 <= _8016;
        252:
            _10295 <= _8007;
        253:
            _10295 <= _7998;
        254:
            _10295 <= _7989;
        255:
            _10295 <= _7980;
        256:
            _10295 <= _7971;
        257:
            _10295 <= _7962;
        258:
            _10295 <= _7953;
        259:
            _10295 <= _7944;
        260:
            _10295 <= _7935;
        261:
            _10295 <= _7926;
        262:
            _10295 <= _7917;
        263:
            _10295 <= _7908;
        264:
            _10295 <= _7899;
        265:
            _10295 <= _7890;
        266:
            _10295 <= _7881;
        267:
            _10295 <= _7872;
        268:
            _10295 <= _7863;
        269:
            _10295 <= _7854;
        270:
            _10295 <= _7845;
        271:
            _10295 <= _7836;
        272:
            _10295 <= _7827;
        273:
            _10295 <= _7818;
        274:
            _10295 <= _7809;
        275:
            _10295 <= _7800;
        276:
            _10295 <= _7791;
        277:
            _10295 <= _7782;
        278:
            _10295 <= _7773;
        279:
            _10295 <= _7764;
        280:
            _10295 <= _7755;
        281:
            _10295 <= _7746;
        282:
            _10295 <= _7737;
        283:
            _10295 <= _7728;
        284:
            _10295 <= _7719;
        285:
            _10295 <= _7710;
        286:
            _10295 <= _7701;
        287:
            _10295 <= _7692;
        288:
            _10295 <= _7683;
        289:
            _10295 <= _7674;
        290:
            _10295 <= _7665;
        291:
            _10295 <= _7656;
        292:
            _10295 <= _7647;
        293:
            _10295 <= _7638;
        294:
            _10295 <= _7629;
        295:
            _10295 <= _7620;
        296:
            _10295 <= _7611;
        297:
            _10295 <= _7602;
        298:
            _10295 <= _7593;
        299:
            _10295 <= _7584;
        300:
            _10295 <= _7575;
        301:
            _10295 <= _7566;
        302:
            _10295 <= _7557;
        303:
            _10295 <= _7548;
        304:
            _10295 <= _7539;
        305:
            _10295 <= _7530;
        306:
            _10295 <= _7521;
        307:
            _10295 <= _7512;
        308:
            _10295 <= _7503;
        309:
            _10295 <= _7494;
        310:
            _10295 <= _7485;
        311:
            _10295 <= _7476;
        312:
            _10295 <= _7467;
        313:
            _10295 <= _7458;
        314:
            _10295 <= _7449;
        315:
            _10295 <= _7440;
        316:
            _10295 <= _7431;
        317:
            _10295 <= _7422;
        318:
            _10295 <= _7413;
        319:
            _10295 <= _7404;
        320:
            _10295 <= _7395;
        321:
            _10295 <= _7386;
        322:
            _10295 <= _7377;
        323:
            _10295 <= _7368;
        324:
            _10295 <= _7359;
        325:
            _10295 <= _7350;
        326:
            _10295 <= _7341;
        327:
            _10295 <= _7332;
        328:
            _10295 <= _7323;
        329:
            _10295 <= _7314;
        330:
            _10295 <= _7305;
        331:
            _10295 <= _7296;
        332:
            _10295 <= _7287;
        333:
            _10295 <= _7278;
        334:
            _10295 <= _7269;
        335:
            _10295 <= _7260;
        336:
            _10295 <= _7251;
        337:
            _10295 <= _7242;
        338:
            _10295 <= _7233;
        339:
            _10295 <= _7224;
        340:
            _10295 <= _7215;
        341:
            _10295 <= _7206;
        342:
            _10295 <= _7197;
        343:
            _10295 <= _7188;
        344:
            _10295 <= _7179;
        345:
            _10295 <= _7170;
        346:
            _10295 <= _7161;
        347:
            _10295 <= _7152;
        348:
            _10295 <= _7143;
        349:
            _10295 <= _7134;
        350:
            _10295 <= _7125;
        351:
            _10295 <= _7116;
        352:
            _10295 <= _7107;
        353:
            _10295 <= _7098;
        354:
            _10295 <= _7089;
        355:
            _10295 <= _7080;
        356:
            _10295 <= _7071;
        357:
            _10295 <= _7062;
        358:
            _10295 <= _7053;
        359:
            _10295 <= _7044;
        360:
            _10295 <= _7035;
        361:
            _10295 <= _7026;
        362:
            _10295 <= _7017;
        363:
            _10295 <= _7008;
        364:
            _10295 <= _6999;
        365:
            _10295 <= _6990;
        366:
            _10295 <= _6981;
        367:
            _10295 <= _6972;
        368:
            _10295 <= _6963;
        369:
            _10295 <= _6954;
        370:
            _10295 <= _6945;
        371:
            _10295 <= _6936;
        372:
            _10295 <= _6927;
        373:
            _10295 <= _6918;
        374:
            _10295 <= _6909;
        375:
            _10295 <= _6900;
        376:
            _10295 <= _6891;
        377:
            _10295 <= _6882;
        378:
            _10295 <= _6873;
        379:
            _10295 <= _6864;
        380:
            _10295 <= _6855;
        381:
            _10295 <= _6846;
        382:
            _10295 <= _6837;
        383:
            _10295 <= _6828;
        384:
            _10295 <= _6819;
        385:
            _10295 <= _6810;
        386:
            _10295 <= _6801;
        387:
            _10295 <= _6792;
        388:
            _10295 <= _6783;
        389:
            _10295 <= _6774;
        390:
            _10295 <= _6765;
        391:
            _10295 <= _6756;
        392:
            _10295 <= _6747;
        393:
            _10295 <= _6738;
        394:
            _10295 <= _6729;
        395:
            _10295 <= _6720;
        396:
            _10295 <= _6711;
        397:
            _10295 <= _6702;
        398:
            _10295 <= _6693;
        399:
            _10295 <= _6684;
        400:
            _10295 <= _6675;
        401:
            _10295 <= _6666;
        402:
            _10295 <= _6657;
        403:
            _10295 <= _6648;
        404:
            _10295 <= _6639;
        405:
            _10295 <= _6630;
        406:
            _10295 <= _6621;
        407:
            _10295 <= _6612;
        408:
            _10295 <= _6603;
        409:
            _10295 <= _6594;
        410:
            _10295 <= _6585;
        411:
            _10295 <= _6576;
        412:
            _10295 <= _6567;
        413:
            _10295 <= _6558;
        414:
            _10295 <= _6549;
        415:
            _10295 <= _6540;
        416:
            _10295 <= _6531;
        417:
            _10295 <= _6522;
        418:
            _10295 <= _6513;
        419:
            _10295 <= _6504;
        420:
            _10295 <= _6495;
        421:
            _10295 <= _6486;
        422:
            _10295 <= _6477;
        423:
            _10295 <= _6468;
        424:
            _10295 <= _6459;
        425:
            _10295 <= _6450;
        426:
            _10295 <= _6441;
        427:
            _10295 <= _6432;
        428:
            _10295 <= _6423;
        429:
            _10295 <= _6414;
        430:
            _10295 <= _6405;
        431:
            _10295 <= _6396;
        432:
            _10295 <= _6387;
        433:
            _10295 <= _6378;
        434:
            _10295 <= _6369;
        435:
            _10295 <= _6360;
        436:
            _10295 <= _6351;
        437:
            _10295 <= _6342;
        438:
            _10295 <= _6333;
        439:
            _10295 <= _6324;
        440:
            _10295 <= _6315;
        441:
            _10295 <= _6306;
        442:
            _10295 <= _6297;
        443:
            _10295 <= _6288;
        444:
            _10295 <= _6279;
        445:
            _10295 <= _6270;
        446:
            _10295 <= _6261;
        447:
            _10295 <= _6252;
        448:
            _10295 <= _6243;
        449:
            _10295 <= _6234;
        450:
            _10295 <= _6225;
        451:
            _10295 <= _6216;
        452:
            _10295 <= _6207;
        453:
            _10295 <= _6198;
        454:
            _10295 <= _6189;
        455:
            _10295 <= _6180;
        456:
            _10295 <= _6171;
        457:
            _10295 <= _6162;
        458:
            _10295 <= _6153;
        459:
            _10295 <= _6144;
        460:
            _10295 <= _6135;
        461:
            _10295 <= _6126;
        462:
            _10295 <= _6117;
        463:
            _10295 <= _6108;
        464:
            _10295 <= _6099;
        465:
            _10295 <= _6090;
        466:
            _10295 <= _6081;
        467:
            _10295 <= _6072;
        468:
            _10295 <= _6063;
        469:
            _10295 <= _6054;
        470:
            _10295 <= _6045;
        471:
            _10295 <= _6036;
        472:
            _10295 <= _6027;
        473:
            _10295 <= _6018;
        474:
            _10295 <= _6009;
        475:
            _10295 <= _6000;
        476:
            _10295 <= _5991;
        477:
            _10295 <= _5982;
        478:
            _10295 <= _5973;
        479:
            _10295 <= _5964;
        480:
            _10295 <= _5955;
        481:
            _10295 <= _5946;
        482:
            _10295 <= _5937;
        483:
            _10295 <= _5928;
        484:
            _10295 <= _5919;
        485:
            _10295 <= _5910;
        486:
            _10295 <= _5901;
        487:
            _10295 <= _5892;
        488:
            _10295 <= _5883;
        489:
            _10295 <= _5874;
        490:
            _10295 <= _5865;
        491:
            _10295 <= _5856;
        492:
            _10295 <= _5847;
        493:
            _10295 <= _5838;
        494:
            _10295 <= _5829;
        495:
            _10295 <= _5820;
        496:
            _10295 <= _5811;
        497:
            _10295 <= _5802;
        498:
            _10295 <= _5793;
        499:
            _10295 <= _5784;
        500:
            _10295 <= _5775;
        501:
            _10295 <= _5766;
        502:
            _10295 <= _5757;
        503:
            _10295 <= _5748;
        504:
            _10295 <= _5739;
        505:
            _10295 <= _5730;
        506:
            _10295 <= _5721;
        507:
            _10295 <= _5712;
        508:
            _10295 <= _5703;
        509:
            _10295 <= _5694;
        510:
            _10295 <= _5685;
        default:
            _10295 <= _5676;
        endcase
    end
    assign _10297 = _10295 < _10296;
    assign _10298 = ~ _10297;
    assign _10301 = _10298 ? _10300 : _10299;
    assign _10303 = _10301 + _10311;
    assign _10313 = _10303 * _10312;
    assign _10314 = _10313[63:0];
    assign _10315 = _1056 < _10314;
    assign _10294 = _10280 & _10293;
    assign _10316 = _10294 & _10315;
    assign _10322 = _10316 ? _10314 : _10321;
    assign _1031 = _10322;
    always @(posedge _1038) begin
        if (_1036)
            _1056 <= _1055;
        else
            _1056 <= _1031;
    end
    assign _10324 = _1053 == _10323;
    assign _1051 = 2'b00;
    assign _10323 = 2'b10;
    assign _10363 = _10286 - _5644;
    assign _10359 = _10283 + _5653;
    assign _10355 = _1047 ? _5662 : _10283;
    assign _10353 = _1059 & _1043;
    assign _10357 = _10353 ? _5662 : _10355;
    assign _10337 = _10283 + _5644;
    assign _10335 = _10291 + _5653;
    assign _10332 = _10286 - _5653;
    assign _10333 = _10291 == _10332;
    assign _10338 = _10333 ? _10337 : _10335;
    assign _10328 = _1047 ? _5662 : _10291;
    assign _10326 = _1059 & _1043;
    assign _10330 = _10326 ? _5653 : _10328;
    assign _10325 = _10280 & _10293;
    assign _10339 = _10325 ? _10338 : _10330;
    assign _1034 = _10339;
    always @(posedge _1038) begin
        if (_1036)
            _10291 <= _5662;
        else
            _10291 <= _1034;
    end
    assign _10292 = _10291 < _10286;
    assign vdd = 1'b1;
    assign _1036 = clear;
    assign _1038 = clock;
    assign _10343 = _1062 + _5653;
    assign _10341 = _1047 ? _5662 : _1062;
    assign _10344 = _1059 ? _10343 : _10341;
    assign _1039 = _10344;
    always @(posedge _1038) begin
        if (_1036)
            _1062 <= _5662;
        else
            _1062 <= _1039;
    end
    assign _10349 = _1062 + _5653;
    assign _10347 = _1047 ? _5662 : _10286;
    assign _10345 = _1059 & _1043;
    assign _10350 = _10345 ? _10349 : _10347;
    assign _1040 = _10350;
    always @(posedge _1038) begin
        if (_1036)
            _10286 <= _5662;
        else
            _10286 <= _1040;
    end
    assign _10287 = _10283 < _10286;
    assign _10288 = _10280 & _10287;
    assign _10293 = _10288 & _10292;
    assign _10351 = _10280 & _10293;
    assign _10352 = _10351 & _10333;
    assign _10360 = _10352 ? _10359 : _10357;
    assign _1041 = _10360;
    always @(posedge _1038) begin
        if (_1036)
            _10283 <= _5662;
        else
            _10283 <= _1041;
    end
    assign _10364 = _10283 == _10363;
    assign _10279 = 2'b01;
    assign _10280 = _1053 == _10279;
    assign _10365 = _10280 & _10364;
    assign _10366 = _10365 & _10333;
    assign _10367 = _10366 ? _10323 : _1053;
    assign _1043 = tile_last;
    assign _1045 = tile_valid;
    assign _1059 = _1058 & _1045;
    assign _10361 = _1059 & _1043;
    assign _10368 = _10361 ? _10279 : _10367;
    assign _1047 = load;
    assign _10369 = _1047 ? _1051 : _10368;
    assign _1048 = _10369;
    always @(posedge _1038) begin
        if (_1036)
            _1053 <= _1051;
        else
            _1053 <= _1048;
    end
    assign _1058 = _1053 == _1051;
    assign ready = _1058;
    assign done_ = _10324;
    assign part1_result = _1056;
    assign part2_result = _1056;
    assign state = _1053;

endmodule
