module day5_opt_a (
    id,
    range_to,
    range_from,
    id_last,
    id_valid,
    clear,
    clock,
    range_last,
    range_valid,
    load,
    part1_result,
    part2_result,
    range_ready,
    id_ready,
    done_,
    phase
);

    input [63:0] id;
    input [63:0] range_to;
    input [63:0] range_from;
    input id_last;
    input id_valid;
    input clear;
    input clock;
    input range_last;
    input range_valid;
    input load;
    output [63:0] part1_result;
    output [63:0] part2_result;
    output range_ready;
    output id_ready;
    output done_;
    output [1:0] phase;

    wire _556;
    wire [63:0] _567;
    wire [63:0] _600;
    wire [63:0] _601;
    wire [63:0] _584;
    wire [63:0] _585;
    wire [63:0] _586;
    wire [63:0] _602;
    wire [63:0] _603;
    wire [63:0] _605;
    wire [63:0] _5;
    reg [63:0] _568;
    wire [63:0] _7353;
    wire [63:0] _7354;
    wire _7347;
    wire [7:0] _617;
    wire _618;
    wire _613;
    wire _619;
    wire [63:0] _623;
    wire _611;
    wire _606;
    wire _612;
    wire [63:0] _624;
    wire [63:0] _7;
    reg [63:0] _622;
    wire [7:0] _630;
    wire _631;
    wire _629;
    wire _632;
    wire [63:0] _636;
    wire _627;
    wire _625;
    wire _628;
    wire [63:0] _637;
    wire [63:0] _8;
    reg [63:0] _635;
    wire [7:0] _643;
    wire _644;
    wire _642;
    wire _645;
    wire [63:0] _649;
    wire _640;
    wire _638;
    wire _641;
    wire [63:0] _650;
    wire [63:0] _9;
    reg [63:0] _648;
    wire [7:0] _656;
    wire _657;
    wire _655;
    wire _658;
    wire [63:0] _662;
    wire _653;
    wire _651;
    wire _654;
    wire [63:0] _663;
    wire [63:0] _10;
    reg [63:0] _661;
    wire [7:0] _669;
    wire _670;
    wire _668;
    wire _671;
    wire [63:0] _675;
    wire _666;
    wire _664;
    wire _667;
    wire [63:0] _676;
    wire [63:0] _11;
    reg [63:0] _674;
    wire [7:0] _682;
    wire _683;
    wire _681;
    wire _684;
    wire [63:0] _688;
    wire _679;
    wire _677;
    wire _680;
    wire [63:0] _689;
    wire [63:0] _12;
    reg [63:0] _687;
    wire [7:0] _695;
    wire _696;
    wire _694;
    wire _697;
    wire [63:0] _701;
    wire _692;
    wire _690;
    wire _693;
    wire [63:0] _702;
    wire [63:0] _13;
    reg [63:0] _700;
    wire [7:0] _708;
    wire _709;
    wire _707;
    wire _710;
    wire [63:0] _714;
    wire _705;
    wire _703;
    wire _706;
    wire [63:0] _715;
    wire [63:0] _14;
    reg [63:0] _713;
    wire [7:0] _721;
    wire _722;
    wire _720;
    wire _723;
    wire [63:0] _727;
    wire _718;
    wire _716;
    wire _719;
    wire [63:0] _728;
    wire [63:0] _15;
    reg [63:0] _726;
    wire [7:0] _734;
    wire _735;
    wire _733;
    wire _736;
    wire [63:0] _740;
    wire _731;
    wire _729;
    wire _732;
    wire [63:0] _741;
    wire [63:0] _16;
    reg [63:0] _739;
    wire [7:0] _747;
    wire _748;
    wire _746;
    wire _749;
    wire [63:0] _753;
    wire _744;
    wire _742;
    wire _745;
    wire [63:0] _754;
    wire [63:0] _17;
    reg [63:0] _752;
    wire [7:0] _760;
    wire _761;
    wire _759;
    wire _762;
    wire [63:0] _766;
    wire _757;
    wire _755;
    wire _758;
    wire [63:0] _767;
    wire [63:0] _18;
    reg [63:0] _765;
    wire [7:0] _773;
    wire _774;
    wire _772;
    wire _775;
    wire [63:0] _779;
    wire _770;
    wire _768;
    wire _771;
    wire [63:0] _780;
    wire [63:0] _19;
    reg [63:0] _778;
    wire [7:0] _786;
    wire _787;
    wire _785;
    wire _788;
    wire [63:0] _792;
    wire _783;
    wire _781;
    wire _784;
    wire [63:0] _793;
    wire [63:0] _20;
    reg [63:0] _791;
    wire [7:0] _799;
    wire _800;
    wire _798;
    wire _801;
    wire [63:0] _805;
    wire _796;
    wire _794;
    wire _797;
    wire [63:0] _806;
    wire [63:0] _21;
    reg [63:0] _804;
    wire [7:0] _812;
    wire _813;
    wire _811;
    wire _814;
    wire [63:0] _818;
    wire _809;
    wire _807;
    wire _810;
    wire [63:0] _819;
    wire [63:0] _22;
    reg [63:0] _817;
    wire [7:0] _825;
    wire _826;
    wire _824;
    wire _827;
    wire [63:0] _831;
    wire _822;
    wire _820;
    wire _823;
    wire [63:0] _832;
    wire [63:0] _23;
    reg [63:0] _830;
    wire [7:0] _838;
    wire _839;
    wire _837;
    wire _840;
    wire [63:0] _844;
    wire _835;
    wire _833;
    wire _836;
    wire [63:0] _845;
    wire [63:0] _24;
    reg [63:0] _843;
    wire [7:0] _851;
    wire _852;
    wire _850;
    wire _853;
    wire [63:0] _857;
    wire _848;
    wire _846;
    wire _849;
    wire [63:0] _858;
    wire [63:0] _25;
    reg [63:0] _856;
    wire [7:0] _864;
    wire _865;
    wire _863;
    wire _866;
    wire [63:0] _870;
    wire _861;
    wire _859;
    wire _862;
    wire [63:0] _871;
    wire [63:0] _26;
    reg [63:0] _869;
    wire [7:0] _877;
    wire _878;
    wire _876;
    wire _879;
    wire [63:0] _883;
    wire _874;
    wire _872;
    wire _875;
    wire [63:0] _884;
    wire [63:0] _27;
    reg [63:0] _882;
    wire [7:0] _890;
    wire _891;
    wire _889;
    wire _892;
    wire [63:0] _896;
    wire _887;
    wire _885;
    wire _888;
    wire [63:0] _897;
    wire [63:0] _28;
    reg [63:0] _895;
    wire [7:0] _903;
    wire _904;
    wire _902;
    wire _905;
    wire [63:0] _909;
    wire _900;
    wire _898;
    wire _901;
    wire [63:0] _910;
    wire [63:0] _29;
    reg [63:0] _908;
    wire [7:0] _916;
    wire _917;
    wire _915;
    wire _918;
    wire [63:0] _922;
    wire _913;
    wire _911;
    wire _914;
    wire [63:0] _923;
    wire [63:0] _30;
    reg [63:0] _921;
    wire [7:0] _929;
    wire _930;
    wire _928;
    wire _931;
    wire [63:0] _935;
    wire _926;
    wire _924;
    wire _927;
    wire [63:0] _936;
    wire [63:0] _31;
    reg [63:0] _934;
    wire [7:0] _942;
    wire _943;
    wire _941;
    wire _944;
    wire [63:0] _948;
    wire _939;
    wire _937;
    wire _940;
    wire [63:0] _949;
    wire [63:0] _32;
    reg [63:0] _947;
    wire [7:0] _955;
    wire _956;
    wire _954;
    wire _957;
    wire [63:0] _961;
    wire _952;
    wire _950;
    wire _953;
    wire [63:0] _962;
    wire [63:0] _33;
    reg [63:0] _960;
    wire [7:0] _968;
    wire _969;
    wire _967;
    wire _970;
    wire [63:0] _974;
    wire _965;
    wire _963;
    wire _966;
    wire [63:0] _975;
    wire [63:0] _34;
    reg [63:0] _973;
    wire [7:0] _981;
    wire _982;
    wire _980;
    wire _983;
    wire [63:0] _987;
    wire _978;
    wire _976;
    wire _979;
    wire [63:0] _988;
    wire [63:0] _35;
    reg [63:0] _986;
    wire [7:0] _994;
    wire _995;
    wire _993;
    wire _996;
    wire [63:0] _1000;
    wire _991;
    wire _989;
    wire _992;
    wire [63:0] _1001;
    wire [63:0] _36;
    reg [63:0] _999;
    wire [7:0] _1007;
    wire _1008;
    wire _1006;
    wire _1009;
    wire [63:0] _1013;
    wire _1004;
    wire _1002;
    wire _1005;
    wire [63:0] _1014;
    wire [63:0] _37;
    reg [63:0] _1012;
    wire [7:0] _1020;
    wire _1021;
    wire _1019;
    wire _1022;
    wire [63:0] _1026;
    wire _1017;
    wire _1015;
    wire _1018;
    wire [63:0] _1027;
    wire [63:0] _38;
    reg [63:0] _1025;
    wire [7:0] _1033;
    wire _1034;
    wire _1032;
    wire _1035;
    wire [63:0] _1039;
    wire _1030;
    wire _1028;
    wire _1031;
    wire [63:0] _1040;
    wire [63:0] _39;
    reg [63:0] _1038;
    wire [7:0] _1046;
    wire _1047;
    wire _1045;
    wire _1048;
    wire [63:0] _1052;
    wire _1043;
    wire _1041;
    wire _1044;
    wire [63:0] _1053;
    wire [63:0] _40;
    reg [63:0] _1051;
    wire [7:0] _1059;
    wire _1060;
    wire _1058;
    wire _1061;
    wire [63:0] _1065;
    wire _1056;
    wire _1054;
    wire _1057;
    wire [63:0] _1066;
    wire [63:0] _41;
    reg [63:0] _1064;
    wire [7:0] _1072;
    wire _1073;
    wire _1071;
    wire _1074;
    wire [63:0] _1078;
    wire _1069;
    wire _1067;
    wire _1070;
    wire [63:0] _1079;
    wire [63:0] _42;
    reg [63:0] _1077;
    wire [7:0] _1085;
    wire _1086;
    wire _1084;
    wire _1087;
    wire [63:0] _1091;
    wire _1082;
    wire _1080;
    wire _1083;
    wire [63:0] _1092;
    wire [63:0] _43;
    reg [63:0] _1090;
    wire [7:0] _1098;
    wire _1099;
    wire _1097;
    wire _1100;
    wire [63:0] _1104;
    wire _1095;
    wire _1093;
    wire _1096;
    wire [63:0] _1105;
    wire [63:0] _44;
    reg [63:0] _1103;
    wire [7:0] _1111;
    wire _1112;
    wire _1110;
    wire _1113;
    wire [63:0] _1117;
    wire _1108;
    wire _1106;
    wire _1109;
    wire [63:0] _1118;
    wire [63:0] _45;
    reg [63:0] _1116;
    wire [7:0] _1124;
    wire _1125;
    wire _1123;
    wire _1126;
    wire [63:0] _1130;
    wire _1121;
    wire _1119;
    wire _1122;
    wire [63:0] _1131;
    wire [63:0] _46;
    reg [63:0] _1129;
    wire [7:0] _1137;
    wire _1138;
    wire _1136;
    wire _1139;
    wire [63:0] _1143;
    wire _1134;
    wire _1132;
    wire _1135;
    wire [63:0] _1144;
    wire [63:0] _47;
    reg [63:0] _1142;
    wire [7:0] _1150;
    wire _1151;
    wire _1149;
    wire _1152;
    wire [63:0] _1156;
    wire _1147;
    wire _1145;
    wire _1148;
    wire [63:0] _1157;
    wire [63:0] _48;
    reg [63:0] _1155;
    wire [7:0] _1163;
    wire _1164;
    wire _1162;
    wire _1165;
    wire [63:0] _1169;
    wire _1160;
    wire _1158;
    wire _1161;
    wire [63:0] _1170;
    wire [63:0] _49;
    reg [63:0] _1168;
    wire [7:0] _1176;
    wire _1177;
    wire _1175;
    wire _1178;
    wire [63:0] _1182;
    wire _1173;
    wire _1171;
    wire _1174;
    wire [63:0] _1183;
    wire [63:0] _50;
    reg [63:0] _1181;
    wire [7:0] _1189;
    wire _1190;
    wire _1188;
    wire _1191;
    wire [63:0] _1195;
    wire _1186;
    wire _1184;
    wire _1187;
    wire [63:0] _1196;
    wire [63:0] _51;
    reg [63:0] _1194;
    wire [7:0] _1202;
    wire _1203;
    wire _1201;
    wire _1204;
    wire [63:0] _1208;
    wire _1199;
    wire _1197;
    wire _1200;
    wire [63:0] _1209;
    wire [63:0] _52;
    reg [63:0] _1207;
    wire [7:0] _1215;
    wire _1216;
    wire _1214;
    wire _1217;
    wire [63:0] _1221;
    wire _1212;
    wire _1210;
    wire _1213;
    wire [63:0] _1222;
    wire [63:0] _53;
    reg [63:0] _1220;
    wire [7:0] _1228;
    wire _1229;
    wire _1227;
    wire _1230;
    wire [63:0] _1234;
    wire _1225;
    wire _1223;
    wire _1226;
    wire [63:0] _1235;
    wire [63:0] _54;
    reg [63:0] _1233;
    wire [7:0] _1241;
    wire _1242;
    wire _1240;
    wire _1243;
    wire [63:0] _1247;
    wire _1238;
    wire _1236;
    wire _1239;
    wire [63:0] _1248;
    wire [63:0] _55;
    reg [63:0] _1246;
    wire [7:0] _1254;
    wire _1255;
    wire _1253;
    wire _1256;
    wire [63:0] _1260;
    wire _1251;
    wire _1249;
    wire _1252;
    wire [63:0] _1261;
    wire [63:0] _56;
    reg [63:0] _1259;
    wire [7:0] _1267;
    wire _1268;
    wire _1266;
    wire _1269;
    wire [63:0] _1273;
    wire _1264;
    wire _1262;
    wire _1265;
    wire [63:0] _1274;
    wire [63:0] _57;
    reg [63:0] _1272;
    wire [7:0] _1280;
    wire _1281;
    wire _1279;
    wire _1282;
    wire [63:0] _1286;
    wire _1277;
    wire _1275;
    wire _1278;
    wire [63:0] _1287;
    wire [63:0] _58;
    reg [63:0] _1285;
    wire [7:0] _1293;
    wire _1294;
    wire _1292;
    wire _1295;
    wire [63:0] _1299;
    wire _1290;
    wire _1288;
    wire _1291;
    wire [63:0] _1300;
    wire [63:0] _59;
    reg [63:0] _1298;
    wire [7:0] _1306;
    wire _1307;
    wire _1305;
    wire _1308;
    wire [63:0] _1312;
    wire _1303;
    wire _1301;
    wire _1304;
    wire [63:0] _1313;
    wire [63:0] _60;
    reg [63:0] _1311;
    wire [7:0] _1319;
    wire _1320;
    wire _1318;
    wire _1321;
    wire [63:0] _1325;
    wire _1316;
    wire _1314;
    wire _1317;
    wire [63:0] _1326;
    wire [63:0] _61;
    reg [63:0] _1324;
    wire [7:0] _1332;
    wire _1333;
    wire _1331;
    wire _1334;
    wire [63:0] _1338;
    wire _1329;
    wire _1327;
    wire _1330;
    wire [63:0] _1339;
    wire [63:0] _62;
    reg [63:0] _1337;
    wire [7:0] _1345;
    wire _1346;
    wire _1344;
    wire _1347;
    wire [63:0] _1351;
    wire _1342;
    wire _1340;
    wire _1343;
    wire [63:0] _1352;
    wire [63:0] _63;
    reg [63:0] _1350;
    wire [7:0] _1358;
    wire _1359;
    wire _1357;
    wire _1360;
    wire [63:0] _1364;
    wire _1355;
    wire _1353;
    wire _1356;
    wire [63:0] _1365;
    wire [63:0] _64;
    reg [63:0] _1363;
    wire [7:0] _1371;
    wire _1372;
    wire _1370;
    wire _1373;
    wire [63:0] _1377;
    wire _1368;
    wire _1366;
    wire _1369;
    wire [63:0] _1378;
    wire [63:0] _65;
    reg [63:0] _1376;
    wire [7:0] _1384;
    wire _1385;
    wire _1383;
    wire _1386;
    wire [63:0] _1390;
    wire _1381;
    wire _1379;
    wire _1382;
    wire [63:0] _1391;
    wire [63:0] _66;
    reg [63:0] _1389;
    wire [7:0] _1397;
    wire _1398;
    wire _1396;
    wire _1399;
    wire [63:0] _1403;
    wire _1394;
    wire _1392;
    wire _1395;
    wire [63:0] _1404;
    wire [63:0] _67;
    reg [63:0] _1402;
    wire [7:0] _1410;
    wire _1411;
    wire _1409;
    wire _1412;
    wire [63:0] _1416;
    wire _1407;
    wire _1405;
    wire _1408;
    wire [63:0] _1417;
    wire [63:0] _68;
    reg [63:0] _1415;
    wire [7:0] _1423;
    wire _1424;
    wire _1422;
    wire _1425;
    wire [63:0] _1429;
    wire _1420;
    wire _1418;
    wire _1421;
    wire [63:0] _1430;
    wire [63:0] _69;
    reg [63:0] _1428;
    wire [7:0] _1436;
    wire _1437;
    wire _1435;
    wire _1438;
    wire [63:0] _1442;
    wire _1433;
    wire _1431;
    wire _1434;
    wire [63:0] _1443;
    wire [63:0] _70;
    reg [63:0] _1441;
    wire [7:0] _1449;
    wire _1450;
    wire _1448;
    wire _1451;
    wire [63:0] _1455;
    wire _1446;
    wire _1444;
    wire _1447;
    wire [63:0] _1456;
    wire [63:0] _71;
    reg [63:0] _1454;
    wire [7:0] _1462;
    wire _1463;
    wire _1461;
    wire _1464;
    wire [63:0] _1468;
    wire _1459;
    wire _1457;
    wire _1460;
    wire [63:0] _1469;
    wire [63:0] _72;
    reg [63:0] _1467;
    wire [7:0] _1475;
    wire _1476;
    wire _1474;
    wire _1477;
    wire [63:0] _1481;
    wire _1472;
    wire _1470;
    wire _1473;
    wire [63:0] _1482;
    wire [63:0] _73;
    reg [63:0] _1480;
    wire [7:0] _1488;
    wire _1489;
    wire _1487;
    wire _1490;
    wire [63:0] _1494;
    wire _1485;
    wire _1483;
    wire _1486;
    wire [63:0] _1495;
    wire [63:0] _74;
    reg [63:0] _1493;
    wire [7:0] _1501;
    wire _1502;
    wire _1500;
    wire _1503;
    wire [63:0] _1507;
    wire _1498;
    wire _1496;
    wire _1499;
    wire [63:0] _1508;
    wire [63:0] _75;
    reg [63:0] _1506;
    wire [7:0] _1514;
    wire _1515;
    wire _1513;
    wire _1516;
    wire [63:0] _1520;
    wire _1511;
    wire _1509;
    wire _1512;
    wire [63:0] _1521;
    wire [63:0] _76;
    reg [63:0] _1519;
    wire [7:0] _1527;
    wire _1528;
    wire _1526;
    wire _1529;
    wire [63:0] _1533;
    wire _1524;
    wire _1522;
    wire _1525;
    wire [63:0] _1534;
    wire [63:0] _77;
    reg [63:0] _1532;
    wire [7:0] _1540;
    wire _1541;
    wire _1539;
    wire _1542;
    wire [63:0] _1546;
    wire _1537;
    wire _1535;
    wire _1538;
    wire [63:0] _1547;
    wire [63:0] _78;
    reg [63:0] _1545;
    wire [7:0] _1553;
    wire _1554;
    wire _1552;
    wire _1555;
    wire [63:0] _1559;
    wire _1550;
    wire _1548;
    wire _1551;
    wire [63:0] _1560;
    wire [63:0] _79;
    reg [63:0] _1558;
    wire [7:0] _1566;
    wire _1567;
    wire _1565;
    wire _1568;
    wire [63:0] _1572;
    wire _1563;
    wire _1561;
    wire _1564;
    wire [63:0] _1573;
    wire [63:0] _80;
    reg [63:0] _1571;
    wire [7:0] _1579;
    wire _1580;
    wire _1578;
    wire _1581;
    wire [63:0] _1585;
    wire _1576;
    wire _1574;
    wire _1577;
    wire [63:0] _1586;
    wire [63:0] _81;
    reg [63:0] _1584;
    wire [7:0] _1592;
    wire _1593;
    wire _1591;
    wire _1594;
    wire [63:0] _1598;
    wire _1589;
    wire _1587;
    wire _1590;
    wire [63:0] _1599;
    wire [63:0] _82;
    reg [63:0] _1597;
    wire [7:0] _1605;
    wire _1606;
    wire _1604;
    wire _1607;
    wire [63:0] _1611;
    wire _1602;
    wire _1600;
    wire _1603;
    wire [63:0] _1612;
    wire [63:0] _83;
    reg [63:0] _1610;
    wire [7:0] _1618;
    wire _1619;
    wire _1617;
    wire _1620;
    wire [63:0] _1624;
    wire _1615;
    wire _1613;
    wire _1616;
    wire [63:0] _1625;
    wire [63:0] _84;
    reg [63:0] _1623;
    wire [7:0] _1631;
    wire _1632;
    wire _1630;
    wire _1633;
    wire [63:0] _1637;
    wire _1628;
    wire _1626;
    wire _1629;
    wire [63:0] _1638;
    wire [63:0] _85;
    reg [63:0] _1636;
    wire [7:0] _1644;
    wire _1645;
    wire _1643;
    wire _1646;
    wire [63:0] _1650;
    wire _1641;
    wire _1639;
    wire _1642;
    wire [63:0] _1651;
    wire [63:0] _86;
    reg [63:0] _1649;
    wire [7:0] _1657;
    wire _1658;
    wire _1656;
    wire _1659;
    wire [63:0] _1663;
    wire _1654;
    wire _1652;
    wire _1655;
    wire [63:0] _1664;
    wire [63:0] _87;
    reg [63:0] _1662;
    wire [7:0] _1670;
    wire _1671;
    wire _1669;
    wire _1672;
    wire [63:0] _1676;
    wire _1667;
    wire _1665;
    wire _1668;
    wire [63:0] _1677;
    wire [63:0] _88;
    reg [63:0] _1675;
    wire [7:0] _1683;
    wire _1684;
    wire _1682;
    wire _1685;
    wire [63:0] _1689;
    wire _1680;
    wire _1678;
    wire _1681;
    wire [63:0] _1690;
    wire [63:0] _89;
    reg [63:0] _1688;
    wire [7:0] _1696;
    wire _1697;
    wire _1695;
    wire _1698;
    wire [63:0] _1702;
    wire _1693;
    wire _1691;
    wire _1694;
    wire [63:0] _1703;
    wire [63:0] _90;
    reg [63:0] _1701;
    wire [7:0] _1709;
    wire _1710;
    wire _1708;
    wire _1711;
    wire [63:0] _1715;
    wire _1706;
    wire _1704;
    wire _1707;
    wire [63:0] _1716;
    wire [63:0] _91;
    reg [63:0] _1714;
    wire [7:0] _1722;
    wire _1723;
    wire _1721;
    wire _1724;
    wire [63:0] _1728;
    wire _1719;
    wire _1717;
    wire _1720;
    wire [63:0] _1729;
    wire [63:0] _92;
    reg [63:0] _1727;
    wire [7:0] _1735;
    wire _1736;
    wire _1734;
    wire _1737;
    wire [63:0] _1741;
    wire _1732;
    wire _1730;
    wire _1733;
    wire [63:0] _1742;
    wire [63:0] _93;
    reg [63:0] _1740;
    wire [7:0] _1748;
    wire _1749;
    wire _1747;
    wire _1750;
    wire [63:0] _1754;
    wire _1745;
    wire _1743;
    wire _1746;
    wire [63:0] _1755;
    wire [63:0] _94;
    reg [63:0] _1753;
    wire [7:0] _1761;
    wire _1762;
    wire _1760;
    wire _1763;
    wire [63:0] _1767;
    wire _1758;
    wire _1756;
    wire _1759;
    wire [63:0] _1768;
    wire [63:0] _95;
    reg [63:0] _1766;
    wire [7:0] _1774;
    wire _1775;
    wire _1773;
    wire _1776;
    wire [63:0] _1780;
    wire _1771;
    wire _1769;
    wire _1772;
    wire [63:0] _1781;
    wire [63:0] _96;
    reg [63:0] _1779;
    wire [7:0] _1787;
    wire _1788;
    wire _1786;
    wire _1789;
    wire [63:0] _1793;
    wire _1784;
    wire _1782;
    wire _1785;
    wire [63:0] _1794;
    wire [63:0] _97;
    reg [63:0] _1792;
    wire [7:0] _1800;
    wire _1801;
    wire _1799;
    wire _1802;
    wire [63:0] _1806;
    wire _1797;
    wire _1795;
    wire _1798;
    wire [63:0] _1807;
    wire [63:0] _98;
    reg [63:0] _1805;
    wire [7:0] _1813;
    wire _1814;
    wire _1812;
    wire _1815;
    wire [63:0] _1819;
    wire _1810;
    wire _1808;
    wire _1811;
    wire [63:0] _1820;
    wire [63:0] _99;
    reg [63:0] _1818;
    wire [7:0] _1826;
    wire _1827;
    wire _1825;
    wire _1828;
    wire [63:0] _1832;
    wire _1823;
    wire _1821;
    wire _1824;
    wire [63:0] _1833;
    wire [63:0] _100;
    reg [63:0] _1831;
    wire [7:0] _1839;
    wire _1840;
    wire _1838;
    wire _1841;
    wire [63:0] _1845;
    wire _1836;
    wire _1834;
    wire _1837;
    wire [63:0] _1846;
    wire [63:0] _101;
    reg [63:0] _1844;
    wire [7:0] _1852;
    wire _1853;
    wire _1851;
    wire _1854;
    wire [63:0] _1858;
    wire _1849;
    wire _1847;
    wire _1850;
    wire [63:0] _1859;
    wire [63:0] _102;
    reg [63:0] _1857;
    wire [7:0] _1865;
    wire _1866;
    wire _1864;
    wire _1867;
    wire [63:0] _1871;
    wire _1862;
    wire _1860;
    wire _1863;
    wire [63:0] _1872;
    wire [63:0] _103;
    reg [63:0] _1870;
    wire [7:0] _1878;
    wire _1879;
    wire _1877;
    wire _1880;
    wire [63:0] _1884;
    wire _1875;
    wire _1873;
    wire _1876;
    wire [63:0] _1885;
    wire [63:0] _104;
    reg [63:0] _1883;
    wire [7:0] _1891;
    wire _1892;
    wire _1890;
    wire _1893;
    wire [63:0] _1897;
    wire _1888;
    wire _1886;
    wire _1889;
    wire [63:0] _1898;
    wire [63:0] _105;
    reg [63:0] _1896;
    wire [7:0] _1904;
    wire _1905;
    wire _1903;
    wire _1906;
    wire [63:0] _1910;
    wire _1901;
    wire _1899;
    wire _1902;
    wire [63:0] _1911;
    wire [63:0] _106;
    reg [63:0] _1909;
    wire [7:0] _1917;
    wire _1918;
    wire _1916;
    wire _1919;
    wire [63:0] _1923;
    wire _1914;
    wire _1912;
    wire _1915;
    wire [63:0] _1924;
    wire [63:0] _107;
    reg [63:0] _1922;
    wire [7:0] _1930;
    wire _1931;
    wire _1929;
    wire _1932;
    wire [63:0] _1936;
    wire _1927;
    wire _1925;
    wire _1928;
    wire [63:0] _1937;
    wire [63:0] _108;
    reg [63:0] _1935;
    wire [7:0] _1943;
    wire _1944;
    wire _1942;
    wire _1945;
    wire [63:0] _1949;
    wire _1940;
    wire _1938;
    wire _1941;
    wire [63:0] _1950;
    wire [63:0] _109;
    reg [63:0] _1948;
    wire [7:0] _1956;
    wire _1957;
    wire _1955;
    wire _1958;
    wire [63:0] _1962;
    wire _1953;
    wire _1951;
    wire _1954;
    wire [63:0] _1963;
    wire [63:0] _110;
    reg [63:0] _1961;
    wire [7:0] _1969;
    wire _1970;
    wire _1968;
    wire _1971;
    wire [63:0] _1975;
    wire _1966;
    wire _1964;
    wire _1967;
    wire [63:0] _1976;
    wire [63:0] _111;
    reg [63:0] _1974;
    wire [7:0] _1982;
    wire _1983;
    wire _1981;
    wire _1984;
    wire [63:0] _1988;
    wire _1979;
    wire _1977;
    wire _1980;
    wire [63:0] _1989;
    wire [63:0] _112;
    reg [63:0] _1987;
    wire [7:0] _1995;
    wire _1996;
    wire _1994;
    wire _1997;
    wire [63:0] _2001;
    wire _1992;
    wire _1990;
    wire _1993;
    wire [63:0] _2002;
    wire [63:0] _113;
    reg [63:0] _2000;
    wire [7:0] _2008;
    wire _2009;
    wire _2007;
    wire _2010;
    wire [63:0] _2014;
    wire _2005;
    wire _2003;
    wire _2006;
    wire [63:0] _2015;
    wire [63:0] _114;
    reg [63:0] _2013;
    wire [7:0] _2021;
    wire _2022;
    wire _2020;
    wire _2023;
    wire [63:0] _2027;
    wire _2018;
    wire _2016;
    wire _2019;
    wire [63:0] _2028;
    wire [63:0] _115;
    reg [63:0] _2026;
    wire [7:0] _2034;
    wire _2035;
    wire _2033;
    wire _2036;
    wire [63:0] _2040;
    wire _2031;
    wire _2029;
    wire _2032;
    wire [63:0] _2041;
    wire [63:0] _116;
    reg [63:0] _2039;
    wire [7:0] _2047;
    wire _2048;
    wire _2046;
    wire _2049;
    wire [63:0] _2053;
    wire _2044;
    wire _2042;
    wire _2045;
    wire [63:0] _2054;
    wire [63:0] _117;
    reg [63:0] _2052;
    wire [7:0] _2060;
    wire _2061;
    wire _2059;
    wire _2062;
    wire [63:0] _2066;
    wire _2057;
    wire _2055;
    wire _2058;
    wire [63:0] _2067;
    wire [63:0] _118;
    reg [63:0] _2065;
    wire [7:0] _2073;
    wire _2074;
    wire _2072;
    wire _2075;
    wire [63:0] _2079;
    wire _2070;
    wire _2068;
    wire _2071;
    wire [63:0] _2080;
    wire [63:0] _119;
    reg [63:0] _2078;
    wire [7:0] _2086;
    wire _2087;
    wire _2085;
    wire _2088;
    wire [63:0] _2092;
    wire _2083;
    wire _2081;
    wire _2084;
    wire [63:0] _2093;
    wire [63:0] _120;
    reg [63:0] _2091;
    wire [7:0] _2099;
    wire _2100;
    wire _2098;
    wire _2101;
    wire [63:0] _2105;
    wire _2096;
    wire _2094;
    wire _2097;
    wire [63:0] _2106;
    wire [63:0] _121;
    reg [63:0] _2104;
    wire [7:0] _2112;
    wire _2113;
    wire _2111;
    wire _2114;
    wire [63:0] _2118;
    wire _2109;
    wire _2107;
    wire _2110;
    wire [63:0] _2119;
    wire [63:0] _122;
    reg [63:0] _2117;
    wire [7:0] _2125;
    wire _2126;
    wire _2124;
    wire _2127;
    wire [63:0] _2131;
    wire _2122;
    wire _2120;
    wire _2123;
    wire [63:0] _2132;
    wire [63:0] _123;
    reg [63:0] _2130;
    wire [7:0] _2138;
    wire _2139;
    wire _2137;
    wire _2140;
    wire [63:0] _2144;
    wire _2135;
    wire _2133;
    wire _2136;
    wire [63:0] _2145;
    wire [63:0] _124;
    reg [63:0] _2143;
    wire [7:0] _2151;
    wire _2152;
    wire _2150;
    wire _2153;
    wire [63:0] _2157;
    wire _2148;
    wire _2146;
    wire _2149;
    wire [63:0] _2158;
    wire [63:0] _125;
    reg [63:0] _2156;
    wire [7:0] _2164;
    wire _2165;
    wire _2163;
    wire _2166;
    wire [63:0] _2170;
    wire _2161;
    wire _2159;
    wire _2162;
    wire [63:0] _2171;
    wire [63:0] _126;
    reg [63:0] _2169;
    wire [7:0] _2177;
    wire _2178;
    wire _2176;
    wire _2179;
    wire [63:0] _2183;
    wire _2174;
    wire _2172;
    wire _2175;
    wire [63:0] _2184;
    wire [63:0] _127;
    reg [63:0] _2182;
    wire [7:0] _2190;
    wire _2191;
    wire _2189;
    wire _2192;
    wire [63:0] _2196;
    wire _2187;
    wire _2185;
    wire _2188;
    wire [63:0] _2197;
    wire [63:0] _128;
    reg [63:0] _2195;
    wire [7:0] _2203;
    wire _2204;
    wire _2202;
    wire _2205;
    wire [63:0] _2209;
    wire _2200;
    wire _2198;
    wire _2201;
    wire [63:0] _2210;
    wire [63:0] _129;
    reg [63:0] _2208;
    wire [7:0] _2216;
    wire _2217;
    wire _2215;
    wire _2218;
    wire [63:0] _2222;
    wire _2213;
    wire _2211;
    wire _2214;
    wire [63:0] _2223;
    wire [63:0] _130;
    reg [63:0] _2221;
    wire [7:0] _2229;
    wire _2230;
    wire _2228;
    wire _2231;
    wire [63:0] _2235;
    wire _2226;
    wire _2224;
    wire _2227;
    wire [63:0] _2236;
    wire [63:0] _131;
    reg [63:0] _2234;
    wire [7:0] _2242;
    wire _2243;
    wire _2241;
    wire _2244;
    wire [63:0] _2248;
    wire _2239;
    wire _2237;
    wire _2240;
    wire [63:0] _2249;
    wire [63:0] _132;
    reg [63:0] _2247;
    wire [7:0] _2255;
    wire _2256;
    wire _2254;
    wire _2257;
    wire [63:0] _2261;
    wire _2252;
    wire _2250;
    wire _2253;
    wire [63:0] _2262;
    wire [63:0] _133;
    reg [63:0] _2260;
    wire [7:0] _2268;
    wire _2269;
    wire _2267;
    wire _2270;
    wire [63:0] _2274;
    wire _2265;
    wire _2263;
    wire _2266;
    wire [63:0] _2275;
    wire [63:0] _134;
    reg [63:0] _2273;
    wire [7:0] _2281;
    wire _2282;
    wire _2280;
    wire _2283;
    wire [63:0] _2287;
    wire _2278;
    wire _2276;
    wire _2279;
    wire [63:0] _2288;
    wire [63:0] _135;
    reg [63:0] _2286;
    wire [7:0] _2294;
    wire _2295;
    wire _2293;
    wire _2296;
    wire [63:0] _2300;
    wire _2291;
    wire _2289;
    wire _2292;
    wire [63:0] _2301;
    wire [63:0] _136;
    reg [63:0] _2299;
    wire [7:0] _2307;
    wire _2308;
    wire _2306;
    wire _2309;
    wire [63:0] _2313;
    wire _2304;
    wire _2302;
    wire _2305;
    wire [63:0] _2314;
    wire [63:0] _137;
    reg [63:0] _2312;
    wire [7:0] _2320;
    wire _2321;
    wire _2319;
    wire _2322;
    wire [63:0] _2326;
    wire _2317;
    wire _2315;
    wire _2318;
    wire [63:0] _2327;
    wire [63:0] _138;
    reg [63:0] _2325;
    wire [7:0] _2333;
    wire _2334;
    wire _2332;
    wire _2335;
    wire [63:0] _2339;
    wire _2330;
    wire _2328;
    wire _2331;
    wire [63:0] _2340;
    wire [63:0] _139;
    reg [63:0] _2338;
    wire [7:0] _2346;
    wire _2347;
    wire _2345;
    wire _2348;
    wire [63:0] _2352;
    wire _2343;
    wire _2341;
    wire _2344;
    wire [63:0] _2353;
    wire [63:0] _140;
    reg [63:0] _2351;
    wire [7:0] _2359;
    wire _2360;
    wire _2358;
    wire _2361;
    wire [63:0] _2365;
    wire _2356;
    wire _2354;
    wire _2357;
    wire [63:0] _2366;
    wire [63:0] _141;
    reg [63:0] _2364;
    wire [7:0] _2372;
    wire _2373;
    wire _2371;
    wire _2374;
    wire [63:0] _2378;
    wire _2369;
    wire _2367;
    wire _2370;
    wire [63:0] _2379;
    wire [63:0] _142;
    reg [63:0] _2377;
    wire [7:0] _2385;
    wire _2386;
    wire _2384;
    wire _2387;
    wire [63:0] _2391;
    wire _2382;
    wire _2380;
    wire _2383;
    wire [63:0] _2392;
    wire [63:0] _143;
    reg [63:0] _2390;
    wire [7:0] _2398;
    wire _2399;
    wire _2397;
    wire _2400;
    wire [63:0] _2404;
    wire _2395;
    wire _2393;
    wire _2396;
    wire [63:0] _2405;
    wire [63:0] _144;
    reg [63:0] _2403;
    wire [7:0] _2411;
    wire _2412;
    wire _2410;
    wire _2413;
    wire [63:0] _2417;
    wire _2408;
    wire _2406;
    wire _2409;
    wire [63:0] _2418;
    wire [63:0] _145;
    reg [63:0] _2416;
    wire [7:0] _2424;
    wire _2425;
    wire _2423;
    wire _2426;
    wire [63:0] _2430;
    wire _2421;
    wire _2419;
    wire _2422;
    wire [63:0] _2431;
    wire [63:0] _146;
    reg [63:0] _2429;
    wire [7:0] _2437;
    wire _2438;
    wire _2436;
    wire _2439;
    wire [63:0] _2443;
    wire _2434;
    wire _2432;
    wire _2435;
    wire [63:0] _2444;
    wire [63:0] _147;
    reg [63:0] _2442;
    wire [7:0] _2450;
    wire _2451;
    wire _2449;
    wire _2452;
    wire [63:0] _2456;
    wire _2447;
    wire _2445;
    wire _2448;
    wire [63:0] _2457;
    wire [63:0] _148;
    reg [63:0] _2455;
    wire [7:0] _2463;
    wire _2464;
    wire _2462;
    wire _2465;
    wire [63:0] _2469;
    wire _2460;
    wire _2458;
    wire _2461;
    wire [63:0] _2470;
    wire [63:0] _149;
    reg [63:0] _2468;
    wire [7:0] _2476;
    wire _2477;
    wire _2475;
    wire _2478;
    wire [63:0] _2482;
    wire _2473;
    wire _2471;
    wire _2474;
    wire [63:0] _2483;
    wire [63:0] _150;
    reg [63:0] _2481;
    wire [7:0] _2489;
    wire _2490;
    wire _2488;
    wire _2491;
    wire [63:0] _2495;
    wire _2486;
    wire _2484;
    wire _2487;
    wire [63:0] _2496;
    wire [63:0] _151;
    reg [63:0] _2494;
    wire [7:0] _2502;
    wire _2503;
    wire _2501;
    wire _2504;
    wire [63:0] _2508;
    wire _2499;
    wire _2497;
    wire _2500;
    wire [63:0] _2509;
    wire [63:0] _152;
    reg [63:0] _2507;
    wire [7:0] _2515;
    wire _2516;
    wire _2514;
    wire _2517;
    wire [63:0] _2521;
    wire _2512;
    wire _2510;
    wire _2513;
    wire [63:0] _2522;
    wire [63:0] _153;
    reg [63:0] _2520;
    wire [7:0] _2528;
    wire _2529;
    wire _2527;
    wire _2530;
    wire [63:0] _2534;
    wire _2525;
    wire _2523;
    wire _2526;
    wire [63:0] _2535;
    wire [63:0] _154;
    reg [63:0] _2533;
    wire [7:0] _2541;
    wire _2542;
    wire _2540;
    wire _2543;
    wire [63:0] _2547;
    wire _2538;
    wire _2536;
    wire _2539;
    wire [63:0] _2548;
    wire [63:0] _155;
    reg [63:0] _2546;
    wire [7:0] _2554;
    wire _2555;
    wire _2553;
    wire _2556;
    wire [63:0] _2560;
    wire _2551;
    wire _2549;
    wire _2552;
    wire [63:0] _2561;
    wire [63:0] _156;
    reg [63:0] _2559;
    wire [7:0] _2567;
    wire _2568;
    wire _2566;
    wire _2569;
    wire [63:0] _2573;
    wire _2564;
    wire _2562;
    wire _2565;
    wire [63:0] _2574;
    wire [63:0] _157;
    reg [63:0] _2572;
    wire [7:0] _2580;
    wire _2581;
    wire _2579;
    wire _2582;
    wire [63:0] _2586;
    wire _2577;
    wire _2575;
    wire _2578;
    wire [63:0] _2587;
    wire [63:0] _158;
    reg [63:0] _2585;
    wire [7:0] _2593;
    wire _2594;
    wire _2592;
    wire _2595;
    wire [63:0] _2599;
    wire _2590;
    wire _2588;
    wire _2591;
    wire [63:0] _2600;
    wire [63:0] _159;
    reg [63:0] _2598;
    wire [7:0] _2606;
    wire _2607;
    wire _2605;
    wire _2608;
    wire [63:0] _2612;
    wire _2603;
    wire _2601;
    wire _2604;
    wire [63:0] _2613;
    wire [63:0] _160;
    reg [63:0] _2611;
    wire [7:0] _2619;
    wire _2620;
    wire _2618;
    wire _2621;
    wire [63:0] _2625;
    wire _2616;
    wire _2614;
    wire _2617;
    wire [63:0] _2626;
    wire [63:0] _161;
    reg [63:0] _2624;
    wire [7:0] _2632;
    wire _2633;
    wire _2631;
    wire _2634;
    wire [63:0] _2638;
    wire _2629;
    wire _2627;
    wire _2630;
    wire [63:0] _2639;
    wire [63:0] _162;
    reg [63:0] _2637;
    wire [7:0] _2645;
    wire _2646;
    wire _2644;
    wire _2647;
    wire [63:0] _2651;
    wire _2642;
    wire _2640;
    wire _2643;
    wire [63:0] _2652;
    wire [63:0] _163;
    reg [63:0] _2650;
    wire [7:0] _2658;
    wire _2659;
    wire _2657;
    wire _2660;
    wire [63:0] _2664;
    wire _2655;
    wire _2653;
    wire _2656;
    wire [63:0] _2665;
    wire [63:0] _164;
    reg [63:0] _2663;
    wire [7:0] _2671;
    wire _2672;
    wire _2670;
    wire _2673;
    wire [63:0] _2677;
    wire _2668;
    wire _2666;
    wire _2669;
    wire [63:0] _2678;
    wire [63:0] _165;
    reg [63:0] _2676;
    wire [7:0] _2684;
    wire _2685;
    wire _2683;
    wire _2686;
    wire [63:0] _2690;
    wire _2681;
    wire _2679;
    wire _2682;
    wire [63:0] _2691;
    wire [63:0] _166;
    reg [63:0] _2689;
    wire [7:0] _2697;
    wire _2698;
    wire _2696;
    wire _2699;
    wire [63:0] _2703;
    wire _2694;
    wire _2692;
    wire _2695;
    wire [63:0] _2704;
    wire [63:0] _167;
    reg [63:0] _2702;
    wire [7:0] _2710;
    wire _2711;
    wire _2709;
    wire _2712;
    wire [63:0] _2716;
    wire _2707;
    wire _2705;
    wire _2708;
    wire [63:0] _2717;
    wire [63:0] _168;
    reg [63:0] _2715;
    wire [7:0] _2723;
    wire _2724;
    wire _2722;
    wire _2725;
    wire [63:0] _2729;
    wire _2720;
    wire _2718;
    wire _2721;
    wire [63:0] _2730;
    wire [63:0] _169;
    reg [63:0] _2728;
    wire [7:0] _2736;
    wire _2737;
    wire _2735;
    wire _2738;
    wire [63:0] _2742;
    wire _2733;
    wire _2731;
    wire _2734;
    wire [63:0] _2743;
    wire [63:0] _170;
    reg [63:0] _2741;
    wire [7:0] _2749;
    wire _2750;
    wire _2748;
    wire _2751;
    wire [63:0] _2755;
    wire _2746;
    wire _2744;
    wire _2747;
    wire [63:0] _2756;
    wire [63:0] _171;
    reg [63:0] _2754;
    wire [7:0] _2762;
    wire _2763;
    wire _2761;
    wire _2764;
    wire [63:0] _2768;
    wire _2759;
    wire _2757;
    wire _2760;
    wire [63:0] _2769;
    wire [63:0] _172;
    reg [63:0] _2767;
    wire [7:0] _2775;
    wire _2776;
    wire _2774;
    wire _2777;
    wire [63:0] _2781;
    wire _2772;
    wire _2770;
    wire _2773;
    wire [63:0] _2782;
    wire [63:0] _173;
    reg [63:0] _2780;
    wire [7:0] _2788;
    wire _2789;
    wire _2787;
    wire _2790;
    wire [63:0] _2794;
    wire _2785;
    wire _2783;
    wire _2786;
    wire [63:0] _2795;
    wire [63:0] _174;
    reg [63:0] _2793;
    wire [7:0] _2801;
    wire _2802;
    wire _2800;
    wire _2803;
    wire [63:0] _2807;
    wire _2798;
    wire _2796;
    wire _2799;
    wire [63:0] _2808;
    wire [63:0] _175;
    reg [63:0] _2806;
    wire [7:0] _2814;
    wire _2815;
    wire _2813;
    wire _2816;
    wire [63:0] _2820;
    wire _2811;
    wire _2809;
    wire _2812;
    wire [63:0] _2821;
    wire [63:0] _176;
    reg [63:0] _2819;
    wire [7:0] _2827;
    wire _2828;
    wire _2826;
    wire _2829;
    wire [63:0] _2833;
    wire _2824;
    wire _2822;
    wire _2825;
    wire [63:0] _2834;
    wire [63:0] _177;
    reg [63:0] _2832;
    wire [7:0] _2840;
    wire _2841;
    wire _2839;
    wire _2842;
    wire [63:0] _2846;
    wire _2837;
    wire _2835;
    wire _2838;
    wire [63:0] _2847;
    wire [63:0] _178;
    reg [63:0] _2845;
    wire [7:0] _2853;
    wire _2854;
    wire _2852;
    wire _2855;
    wire [63:0] _2859;
    wire _2850;
    wire _2848;
    wire _2851;
    wire [63:0] _2860;
    wire [63:0] _179;
    reg [63:0] _2858;
    wire [7:0] _2866;
    wire _2867;
    wire _2865;
    wire _2868;
    wire [63:0] _2872;
    wire _2863;
    wire _2861;
    wire _2864;
    wire [63:0] _2873;
    wire [63:0] _180;
    reg [63:0] _2871;
    wire [7:0] _2879;
    wire _2880;
    wire _2878;
    wire _2881;
    wire [63:0] _2885;
    wire _2876;
    wire _2874;
    wire _2877;
    wire [63:0] _2886;
    wire [63:0] _181;
    reg [63:0] _2884;
    wire [7:0] _2892;
    wire _2893;
    wire _2891;
    wire _2894;
    wire [63:0] _2898;
    wire _2889;
    wire _2887;
    wire _2890;
    wire [63:0] _2899;
    wire [63:0] _182;
    reg [63:0] _2897;
    wire [7:0] _2905;
    wire _2906;
    wire _2904;
    wire _2907;
    wire [63:0] _2911;
    wire _2902;
    wire _2900;
    wire _2903;
    wire [63:0] _2912;
    wire [63:0] _183;
    reg [63:0] _2910;
    wire [7:0] _2918;
    wire _2919;
    wire _2917;
    wire _2920;
    wire [63:0] _2924;
    wire _2915;
    wire _2913;
    wire _2916;
    wire [63:0] _2925;
    wire [63:0] _184;
    reg [63:0] _2923;
    wire [7:0] _2931;
    wire _2932;
    wire _2930;
    wire _2933;
    wire [63:0] _2937;
    wire _2928;
    wire _2926;
    wire _2929;
    wire [63:0] _2938;
    wire [63:0] _185;
    reg [63:0] _2936;
    wire [7:0] _2944;
    wire _2945;
    wire _2943;
    wire _2946;
    wire [63:0] _2950;
    wire _2941;
    wire _2939;
    wire _2942;
    wire [63:0] _2951;
    wire [63:0] _186;
    reg [63:0] _2949;
    wire [7:0] _2957;
    wire _2958;
    wire _2956;
    wire _2959;
    wire [63:0] _2963;
    wire _2954;
    wire _2952;
    wire _2955;
    wire [63:0] _2964;
    wire [63:0] _187;
    reg [63:0] _2962;
    wire [7:0] _2970;
    wire _2971;
    wire _2969;
    wire _2972;
    wire [63:0] _2976;
    wire _2967;
    wire _2965;
    wire _2968;
    wire [63:0] _2977;
    wire [63:0] _188;
    reg [63:0] _2975;
    wire [7:0] _2983;
    wire _2984;
    wire _2982;
    wire _2985;
    wire [63:0] _2989;
    wire _2980;
    wire _2978;
    wire _2981;
    wire [63:0] _2990;
    wire [63:0] _189;
    reg [63:0] _2988;
    wire [7:0] _2996;
    wire _2997;
    wire _2995;
    wire _2998;
    wire [63:0] _3002;
    wire _2993;
    wire _2991;
    wire _2994;
    wire [63:0] _3003;
    wire [63:0] _190;
    reg [63:0] _3001;
    wire [7:0] _3009;
    wire _3010;
    wire _3008;
    wire _3011;
    wire [63:0] _3015;
    wire _3006;
    wire _3004;
    wire _3007;
    wire [63:0] _3016;
    wire [63:0] _191;
    reg [63:0] _3014;
    wire [7:0] _3022;
    wire _3023;
    wire _3021;
    wire _3024;
    wire [63:0] _3028;
    wire _3019;
    wire _3017;
    wire _3020;
    wire [63:0] _3029;
    wire [63:0] _192;
    reg [63:0] _3027;
    wire [7:0] _3035;
    wire _3036;
    wire _3034;
    wire _3037;
    wire [63:0] _3041;
    wire _3032;
    wire _3030;
    wire _3033;
    wire [63:0] _3042;
    wire [63:0] _193;
    reg [63:0] _3040;
    wire [7:0] _3048;
    wire _3049;
    wire _3047;
    wire _3050;
    wire [63:0] _3054;
    wire _3045;
    wire _3043;
    wire _3046;
    wire [63:0] _3055;
    wire [63:0] _194;
    reg [63:0] _3053;
    wire [7:0] _3061;
    wire _3062;
    wire _3060;
    wire _3063;
    wire [63:0] _3067;
    wire _3058;
    wire _3056;
    wire _3059;
    wire [63:0] _3068;
    wire [63:0] _195;
    reg [63:0] _3066;
    wire [7:0] _3074;
    wire _3075;
    wire _3073;
    wire _3076;
    wire [63:0] _3080;
    wire _3071;
    wire _3069;
    wire _3072;
    wire [63:0] _3081;
    wire [63:0] _196;
    reg [63:0] _3079;
    wire [7:0] _3087;
    wire _3088;
    wire _3086;
    wire _3089;
    wire [63:0] _3093;
    wire _3084;
    wire _3082;
    wire _3085;
    wire [63:0] _3094;
    wire [63:0] _197;
    reg [63:0] _3092;
    wire [7:0] _3100;
    wire _3101;
    wire _3099;
    wire _3102;
    wire [63:0] _3106;
    wire _3097;
    wire _3095;
    wire _3098;
    wire [63:0] _3107;
    wire [63:0] _198;
    reg [63:0] _3105;
    wire [7:0] _3113;
    wire _3114;
    wire _3112;
    wire _3115;
    wire [63:0] _3119;
    wire _3110;
    wire _3108;
    wire _3111;
    wire [63:0] _3120;
    wire [63:0] _199;
    reg [63:0] _3118;
    wire [7:0] _3126;
    wire _3127;
    wire _3125;
    wire _3128;
    wire [63:0] _3132;
    wire _3123;
    wire _3121;
    wire _3124;
    wire [63:0] _3133;
    wire [63:0] _200;
    reg [63:0] _3131;
    wire [7:0] _3139;
    wire _3140;
    wire _3138;
    wire _3141;
    wire [63:0] _3145;
    wire _3136;
    wire _3134;
    wire _3137;
    wire [63:0] _3146;
    wire [63:0] _201;
    reg [63:0] _3144;
    wire [7:0] _3152;
    wire _3153;
    wire _3151;
    wire _3154;
    wire [63:0] _3158;
    wire _3149;
    wire _3147;
    wire _3150;
    wire [63:0] _3159;
    wire [63:0] _202;
    reg [63:0] _3157;
    wire [7:0] _3165;
    wire _3166;
    wire _3164;
    wire _3167;
    wire [63:0] _3171;
    wire _3162;
    wire _3160;
    wire _3163;
    wire [63:0] _3172;
    wire [63:0] _203;
    reg [63:0] _3170;
    wire [7:0] _3178;
    wire _3179;
    wire _3177;
    wire _3180;
    wire [63:0] _3184;
    wire _3175;
    wire _3173;
    wire _3176;
    wire [63:0] _3185;
    wire [63:0] _204;
    reg [63:0] _3183;
    wire [7:0] _3191;
    wire _3192;
    wire _3190;
    wire _3193;
    wire [63:0] _3197;
    wire _3188;
    wire _3186;
    wire _3189;
    wire [63:0] _3198;
    wire [63:0] _205;
    reg [63:0] _3196;
    wire [7:0] _3204;
    wire _3205;
    wire _3203;
    wire _3206;
    wire [63:0] _3210;
    wire _3201;
    wire _3199;
    wire _3202;
    wire [63:0] _3211;
    wire [63:0] _206;
    reg [63:0] _3209;
    wire [7:0] _3217;
    wire _3218;
    wire _3216;
    wire _3219;
    wire [63:0] _3223;
    wire _3214;
    wire _3212;
    wire _3215;
    wire [63:0] _3224;
    wire [63:0] _207;
    reg [63:0] _3222;
    wire [7:0] _3230;
    wire _3231;
    wire _3229;
    wire _3232;
    wire [63:0] _3236;
    wire _3227;
    wire _3225;
    wire _3228;
    wire [63:0] _3237;
    wire [63:0] _208;
    reg [63:0] _3235;
    wire [7:0] _3243;
    wire _3244;
    wire _3242;
    wire _3245;
    wire [63:0] _3249;
    wire _3240;
    wire _3238;
    wire _3241;
    wire [63:0] _3250;
    wire [63:0] _209;
    reg [63:0] _3248;
    wire [7:0] _3256;
    wire _3257;
    wire _3255;
    wire _3258;
    wire [63:0] _3262;
    wire _3253;
    wire _3251;
    wire _3254;
    wire [63:0] _3263;
    wire [63:0] _210;
    reg [63:0] _3261;
    wire [7:0] _3269;
    wire _3270;
    wire _3268;
    wire _3271;
    wire [63:0] _3275;
    wire _3266;
    wire _3264;
    wire _3267;
    wire [63:0] _3276;
    wire [63:0] _211;
    reg [63:0] _3274;
    wire [7:0] _3282;
    wire _3283;
    wire _3281;
    wire _3284;
    wire [63:0] _3288;
    wire _3279;
    wire _3277;
    wire _3280;
    wire [63:0] _3289;
    wire [63:0] _212;
    reg [63:0] _3287;
    wire [7:0] _3295;
    wire _3296;
    wire _3294;
    wire _3297;
    wire [63:0] _3301;
    wire _3292;
    wire _3290;
    wire _3293;
    wire [63:0] _3302;
    wire [63:0] _213;
    reg [63:0] _3300;
    wire [7:0] _3308;
    wire _3309;
    wire _3307;
    wire _3310;
    wire [63:0] _3314;
    wire _3305;
    wire _3303;
    wire _3306;
    wire [63:0] _3315;
    wire [63:0] _214;
    reg [63:0] _3313;
    wire [7:0] _3321;
    wire _3322;
    wire _3320;
    wire _3323;
    wire [63:0] _3327;
    wire _3318;
    wire _3316;
    wire _3319;
    wire [63:0] _3328;
    wire [63:0] _215;
    reg [63:0] _3326;
    wire [7:0] _3334;
    wire _3335;
    wire _3333;
    wire _3336;
    wire [63:0] _3340;
    wire _3331;
    wire _3329;
    wire _3332;
    wire [63:0] _3341;
    wire [63:0] _216;
    reg [63:0] _3339;
    wire [7:0] _3347;
    wire _3348;
    wire _3346;
    wire _3349;
    wire [63:0] _3353;
    wire _3344;
    wire _3342;
    wire _3345;
    wire [63:0] _3354;
    wire [63:0] _217;
    reg [63:0] _3352;
    wire [7:0] _3360;
    wire _3361;
    wire _3359;
    wire _3362;
    wire [63:0] _3366;
    wire _3357;
    wire _3355;
    wire _3358;
    wire [63:0] _3367;
    wire [63:0] _218;
    reg [63:0] _3365;
    wire [7:0] _3373;
    wire _3374;
    wire _3372;
    wire _3375;
    wire [63:0] _3379;
    wire _3370;
    wire _3368;
    wire _3371;
    wire [63:0] _3380;
    wire [63:0] _219;
    reg [63:0] _3378;
    wire [7:0] _3386;
    wire _3387;
    wire _3385;
    wire _3388;
    wire [63:0] _3392;
    wire _3383;
    wire _3381;
    wire _3384;
    wire [63:0] _3393;
    wire [63:0] _220;
    reg [63:0] _3391;
    wire [7:0] _3399;
    wire _3400;
    wire _3398;
    wire _3401;
    wire [63:0] _3405;
    wire _3396;
    wire _3394;
    wire _3397;
    wire [63:0] _3406;
    wire [63:0] _221;
    reg [63:0] _3404;
    wire [7:0] _3412;
    wire _3413;
    wire _3411;
    wire _3414;
    wire [63:0] _3418;
    wire _3409;
    wire _3407;
    wire _3410;
    wire [63:0] _3419;
    wire [63:0] _222;
    reg [63:0] _3417;
    wire [7:0] _3425;
    wire _3426;
    wire _3424;
    wire _3427;
    wire [63:0] _3431;
    wire _3422;
    wire _3420;
    wire _3423;
    wire [63:0] _3432;
    wire [63:0] _223;
    reg [63:0] _3430;
    wire [7:0] _3438;
    wire _3439;
    wire _3437;
    wire _3440;
    wire [63:0] _3444;
    wire _3435;
    wire _3433;
    wire _3436;
    wire [63:0] _3445;
    wire [63:0] _224;
    reg [63:0] _3443;
    wire [7:0] _3451;
    wire _3452;
    wire _3450;
    wire _3453;
    wire [63:0] _3457;
    wire _3448;
    wire _3446;
    wire _3449;
    wire [63:0] _3458;
    wire [63:0] _225;
    reg [63:0] _3456;
    wire [7:0] _3464;
    wire _3465;
    wire _3463;
    wire _3466;
    wire [63:0] _3470;
    wire _3461;
    wire _3459;
    wire _3462;
    wire [63:0] _3471;
    wire [63:0] _226;
    reg [63:0] _3469;
    wire [7:0] _3477;
    wire _3478;
    wire _3476;
    wire _3479;
    wire [63:0] _3483;
    wire _3474;
    wire _3472;
    wire _3475;
    wire [63:0] _3484;
    wire [63:0] _227;
    reg [63:0] _3482;
    wire [7:0] _3490;
    wire _3491;
    wire _3489;
    wire _3492;
    wire [63:0] _3496;
    wire _3487;
    wire _3485;
    wire _3488;
    wire [63:0] _3497;
    wire [63:0] _228;
    reg [63:0] _3495;
    wire [7:0] _3503;
    wire _3504;
    wire _3502;
    wire _3505;
    wire [63:0] _3509;
    wire _3500;
    wire _3498;
    wire _3501;
    wire [63:0] _3510;
    wire [63:0] _229;
    reg [63:0] _3508;
    wire [7:0] _3516;
    wire _3517;
    wire _3515;
    wire _3518;
    wire [63:0] _3522;
    wire _3513;
    wire _3511;
    wire _3514;
    wire [63:0] _3523;
    wire [63:0] _230;
    reg [63:0] _3521;
    wire [7:0] _3529;
    wire _3530;
    wire _3528;
    wire _3531;
    wire [63:0] _3535;
    wire _3526;
    wire _3524;
    wire _3527;
    wire [63:0] _3536;
    wire [63:0] _231;
    reg [63:0] _3534;
    wire [7:0] _3542;
    wire _3543;
    wire _3541;
    wire _3544;
    wire [63:0] _3548;
    wire _3539;
    wire _3537;
    wire _3540;
    wire [63:0] _3549;
    wire [63:0] _232;
    reg [63:0] _3547;
    wire [7:0] _3555;
    wire _3556;
    wire _3554;
    wire _3557;
    wire [63:0] _3561;
    wire _3552;
    wire _3550;
    wire _3553;
    wire [63:0] _3562;
    wire [63:0] _233;
    reg [63:0] _3560;
    wire [7:0] _3568;
    wire _3569;
    wire _3567;
    wire _3570;
    wire [63:0] _3574;
    wire _3565;
    wire _3563;
    wire _3566;
    wire [63:0] _3575;
    wire [63:0] _234;
    reg [63:0] _3573;
    wire [7:0] _3581;
    wire _3582;
    wire _3580;
    wire _3583;
    wire [63:0] _3587;
    wire _3578;
    wire _3576;
    wire _3579;
    wire [63:0] _3588;
    wire [63:0] _235;
    reg [63:0] _3586;
    wire [7:0] _3594;
    wire _3595;
    wire _3593;
    wire _3596;
    wire [63:0] _3600;
    wire _3591;
    wire _3589;
    wire _3592;
    wire [63:0] _3601;
    wire [63:0] _236;
    reg [63:0] _3599;
    wire [7:0] _3607;
    wire _3608;
    wire _3606;
    wire _3609;
    wire [63:0] _3613;
    wire _3604;
    wire _3602;
    wire _3605;
    wire [63:0] _3614;
    wire [63:0] _237;
    reg [63:0] _3612;
    wire [7:0] _3620;
    wire _3621;
    wire _3619;
    wire _3622;
    wire [63:0] _3626;
    wire _3617;
    wire _3615;
    wire _3618;
    wire [63:0] _3627;
    wire [63:0] _238;
    reg [63:0] _3625;
    wire [7:0] _3633;
    wire _3634;
    wire _3632;
    wire _3635;
    wire [63:0] _3639;
    wire _3630;
    wire _3628;
    wire _3631;
    wire [63:0] _3640;
    wire [63:0] _239;
    reg [63:0] _3638;
    wire [7:0] _3646;
    wire _3647;
    wire _3645;
    wire _3648;
    wire [63:0] _3652;
    wire _3643;
    wire _3641;
    wire _3644;
    wire [63:0] _3653;
    wire [63:0] _240;
    reg [63:0] _3651;
    wire [7:0] _3659;
    wire _3660;
    wire _3658;
    wire _3661;
    wire [63:0] _3665;
    wire _3656;
    wire _3654;
    wire _3657;
    wire [63:0] _3666;
    wire [63:0] _241;
    reg [63:0] _3664;
    wire [7:0] _3672;
    wire _3673;
    wire _3671;
    wire _3674;
    wire [63:0] _3678;
    wire _3669;
    wire _3667;
    wire _3670;
    wire [63:0] _3679;
    wire [63:0] _242;
    reg [63:0] _3677;
    wire [7:0] _3685;
    wire _3686;
    wire _3684;
    wire _3687;
    wire [63:0] _3691;
    wire _3682;
    wire _3680;
    wire _3683;
    wire [63:0] _3692;
    wire [63:0] _243;
    reg [63:0] _3690;
    wire [7:0] _3698;
    wire _3699;
    wire _3697;
    wire _3700;
    wire [63:0] _3704;
    wire _3695;
    wire _3693;
    wire _3696;
    wire [63:0] _3705;
    wire [63:0] _244;
    reg [63:0] _3703;
    wire [7:0] _3711;
    wire _3712;
    wire _3710;
    wire _3713;
    wire [63:0] _3717;
    wire _3708;
    wire _3706;
    wire _3709;
    wire [63:0] _3718;
    wire [63:0] _245;
    reg [63:0] _3716;
    wire [7:0] _3724;
    wire _3725;
    wire _3723;
    wire _3726;
    wire [63:0] _3730;
    wire _3721;
    wire _3719;
    wire _3722;
    wire [63:0] _3731;
    wire [63:0] _246;
    reg [63:0] _3729;
    wire [7:0] _3737;
    wire _3738;
    wire _3736;
    wire _3739;
    wire [63:0] _3743;
    wire _3734;
    wire _3732;
    wire _3735;
    wire [63:0] _3744;
    wire [63:0] _247;
    reg [63:0] _3742;
    wire [7:0] _3750;
    wire _3751;
    wire _3749;
    wire _3752;
    wire [63:0] _3756;
    wire _3747;
    wire _3745;
    wire _3748;
    wire [63:0] _3757;
    wire [63:0] _248;
    reg [63:0] _3755;
    wire [7:0] _3763;
    wire _3764;
    wire _3762;
    wire _3765;
    wire [63:0] _3769;
    wire _3760;
    wire _3758;
    wire _3761;
    wire [63:0] _3770;
    wire [63:0] _249;
    reg [63:0] _3768;
    wire [7:0] _3776;
    wire _3777;
    wire _3775;
    wire _3778;
    wire [63:0] _3782;
    wire _3773;
    wire _3771;
    wire _3774;
    wire [63:0] _3783;
    wire [63:0] _250;
    reg [63:0] _3781;
    wire [7:0] _3789;
    wire _3790;
    wire _3788;
    wire _3791;
    wire [63:0] _3795;
    wire _3786;
    wire _3784;
    wire _3787;
    wire [63:0] _3796;
    wire [63:0] _251;
    reg [63:0] _3794;
    wire [7:0] _3802;
    wire _3803;
    wire _3801;
    wire _3804;
    wire [63:0] _3808;
    wire _3799;
    wire _3797;
    wire _3800;
    wire [63:0] _3809;
    wire [63:0] _252;
    reg [63:0] _3807;
    wire [7:0] _3815;
    wire _3816;
    wire _3814;
    wire _3817;
    wire [63:0] _3821;
    wire _3812;
    wire _3810;
    wire _3813;
    wire [63:0] _3822;
    wire [63:0] _253;
    reg [63:0] _3820;
    wire [7:0] _3828;
    wire _3829;
    wire _3827;
    wire _3830;
    wire [63:0] _3834;
    wire _3825;
    wire _3823;
    wire _3826;
    wire [63:0] _3835;
    wire [63:0] _254;
    reg [63:0] _3833;
    wire [7:0] _3841;
    wire _3842;
    wire _3840;
    wire _3843;
    wire [63:0] _3847;
    wire _3838;
    wire _3836;
    wire _3839;
    wire [63:0] _3848;
    wire [63:0] _255;
    reg [63:0] _3846;
    wire [7:0] _3854;
    wire _3855;
    wire _3853;
    wire _3856;
    wire [63:0] _3860;
    wire _3851;
    wire _3849;
    wire _3852;
    wire [63:0] _3861;
    wire [63:0] _256;
    reg [63:0] _3859;
    wire [7:0] _3867;
    wire _3868;
    wire _3866;
    wire _3869;
    wire [63:0] _3873;
    wire _3864;
    wire _3862;
    wire _3865;
    wire [63:0] _3874;
    wire [63:0] _257;
    reg [63:0] _3872;
    wire [7:0] _3880;
    wire _3881;
    wire _3879;
    wire _3882;
    wire [63:0] _3886;
    wire _3877;
    wire _3875;
    wire _3878;
    wire [63:0] _3887;
    wire [63:0] _258;
    reg [63:0] _3885;
    wire [7:0] _3893;
    wire _3894;
    wire _3892;
    wire _3895;
    wire [63:0] _3899;
    wire _3890;
    wire _3888;
    wire _3891;
    wire [63:0] _3900;
    wire [63:0] _259;
    reg [63:0] _3898;
    wire [7:0] _3906;
    wire _3907;
    wire _3905;
    wire _3908;
    wire [63:0] _3912;
    wire _3903;
    wire _3901;
    wire _3904;
    wire [63:0] _3913;
    wire [63:0] _260;
    reg [63:0] _3911;
    wire [7:0] _3919;
    wire _3920;
    wire _3918;
    wire _3921;
    wire [63:0] _3925;
    wire _3916;
    wire _3914;
    wire _3917;
    wire [63:0] _3926;
    wire [63:0] _261;
    reg [63:0] _3924;
    wire [63:0] _3927;
    wire [63:0] _3929;
    wire [63:0] _262;
    reg [63:0] _583;
    wire [63:0] _598;
    wire [63:0] _599;
    wire [7:0] _3935;
    wire _3936;
    wire _3934;
    wire _3937;
    wire [63:0] _3941;
    wire _3932;
    wire _3930;
    wire _3933;
    wire [63:0] _3942;
    wire [63:0] _263;
    reg [63:0] _3940;
    reg [63:0] _7343;
    wire _7344;
    wire _7345;
    wire _7346;
    wire _7348;
    wire [7:0] _7292;
    wire [7:0] _7293;
    wire _7294;
    wire _3949;
    wire _3947;
    wire _3950;
    wire [63:0] _3954;
    wire _3945;
    wire _3943;
    wire _3946;
    wire [63:0] _3955;
    wire [63:0] _264;
    reg [63:0] _3953;
    wire _3962;
    wire _3960;
    wire _3963;
    wire [63:0] _3967;
    wire _3958;
    wire _3956;
    wire _3959;
    wire [63:0] _3968;
    wire [63:0] _265;
    reg [63:0] _3966;
    wire _3975;
    wire _3973;
    wire _3976;
    wire [63:0] _3980;
    wire _3971;
    wire _3969;
    wire _3972;
    wire [63:0] _3981;
    wire [63:0] _266;
    reg [63:0] _3979;
    wire _3988;
    wire _3986;
    wire _3989;
    wire [63:0] _3993;
    wire _3984;
    wire _3982;
    wire _3985;
    wire [63:0] _3994;
    wire [63:0] _267;
    reg [63:0] _3992;
    wire _4001;
    wire _3999;
    wire _4002;
    wire [63:0] _4006;
    wire _3997;
    wire _3995;
    wire _3998;
    wire [63:0] _4007;
    wire [63:0] _268;
    reg [63:0] _4005;
    wire _4014;
    wire _4012;
    wire _4015;
    wire [63:0] _4019;
    wire _4010;
    wire _4008;
    wire _4011;
    wire [63:0] _4020;
    wire [63:0] _269;
    reg [63:0] _4018;
    wire _4027;
    wire _4025;
    wire _4028;
    wire [63:0] _4032;
    wire _4023;
    wire _4021;
    wire _4024;
    wire [63:0] _4033;
    wire [63:0] _270;
    reg [63:0] _4031;
    wire _4040;
    wire _4038;
    wire _4041;
    wire [63:0] _4045;
    wire _4036;
    wire _4034;
    wire _4037;
    wire [63:0] _4046;
    wire [63:0] _271;
    reg [63:0] _4044;
    wire _4053;
    wire _4051;
    wire _4054;
    wire [63:0] _4058;
    wire _4049;
    wire _4047;
    wire _4050;
    wire [63:0] _4059;
    wire [63:0] _272;
    reg [63:0] _4057;
    wire _4066;
    wire _4064;
    wire _4067;
    wire [63:0] _4071;
    wire _4062;
    wire _4060;
    wire _4063;
    wire [63:0] _4072;
    wire [63:0] _273;
    reg [63:0] _4070;
    wire _4079;
    wire _4077;
    wire _4080;
    wire [63:0] _4084;
    wire _4075;
    wire _4073;
    wire _4076;
    wire [63:0] _4085;
    wire [63:0] _274;
    reg [63:0] _4083;
    wire _4092;
    wire _4090;
    wire _4093;
    wire [63:0] _4097;
    wire _4088;
    wire _4086;
    wire _4089;
    wire [63:0] _4098;
    wire [63:0] _275;
    reg [63:0] _4096;
    wire _4105;
    wire _4103;
    wire _4106;
    wire [63:0] _4110;
    wire _4101;
    wire _4099;
    wire _4102;
    wire [63:0] _4111;
    wire [63:0] _276;
    reg [63:0] _4109;
    wire _4118;
    wire _4116;
    wire _4119;
    wire [63:0] _4123;
    wire _4114;
    wire _4112;
    wire _4115;
    wire [63:0] _4124;
    wire [63:0] _277;
    reg [63:0] _4122;
    wire _4131;
    wire _4129;
    wire _4132;
    wire [63:0] _4136;
    wire _4127;
    wire _4125;
    wire _4128;
    wire [63:0] _4137;
    wire [63:0] _278;
    reg [63:0] _4135;
    wire _4144;
    wire _4142;
    wire _4145;
    wire [63:0] _4149;
    wire _4140;
    wire _4138;
    wire _4141;
    wire [63:0] _4150;
    wire [63:0] _279;
    reg [63:0] _4148;
    wire _4157;
    wire _4155;
    wire _4158;
    wire [63:0] _4162;
    wire _4153;
    wire _4151;
    wire _4154;
    wire [63:0] _4163;
    wire [63:0] _280;
    reg [63:0] _4161;
    wire _4170;
    wire _4168;
    wire _4171;
    wire [63:0] _4175;
    wire _4166;
    wire _4164;
    wire _4167;
    wire [63:0] _4176;
    wire [63:0] _281;
    reg [63:0] _4174;
    wire _4183;
    wire _4181;
    wire _4184;
    wire [63:0] _4188;
    wire _4179;
    wire _4177;
    wire _4180;
    wire [63:0] _4189;
    wire [63:0] _282;
    reg [63:0] _4187;
    wire _4196;
    wire _4194;
    wire _4197;
    wire [63:0] _4201;
    wire _4192;
    wire _4190;
    wire _4193;
    wire [63:0] _4202;
    wire [63:0] _283;
    reg [63:0] _4200;
    wire _4209;
    wire _4207;
    wire _4210;
    wire [63:0] _4214;
    wire _4205;
    wire _4203;
    wire _4206;
    wire [63:0] _4215;
    wire [63:0] _284;
    reg [63:0] _4213;
    wire _4222;
    wire _4220;
    wire _4223;
    wire [63:0] _4227;
    wire _4218;
    wire _4216;
    wire _4219;
    wire [63:0] _4228;
    wire [63:0] _285;
    reg [63:0] _4226;
    wire _4235;
    wire _4233;
    wire _4236;
    wire [63:0] _4240;
    wire _4231;
    wire _4229;
    wire _4232;
    wire [63:0] _4241;
    wire [63:0] _286;
    reg [63:0] _4239;
    wire _4248;
    wire _4246;
    wire _4249;
    wire [63:0] _4253;
    wire _4244;
    wire _4242;
    wire _4245;
    wire [63:0] _4254;
    wire [63:0] _287;
    reg [63:0] _4252;
    wire _4261;
    wire _4259;
    wire _4262;
    wire [63:0] _4266;
    wire _4257;
    wire _4255;
    wire _4258;
    wire [63:0] _4267;
    wire [63:0] _288;
    reg [63:0] _4265;
    wire _4274;
    wire _4272;
    wire _4275;
    wire [63:0] _4279;
    wire _4270;
    wire _4268;
    wire _4271;
    wire [63:0] _4280;
    wire [63:0] _289;
    reg [63:0] _4278;
    wire _4287;
    wire _4285;
    wire _4288;
    wire [63:0] _4292;
    wire _4283;
    wire _4281;
    wire _4284;
    wire [63:0] _4293;
    wire [63:0] _290;
    reg [63:0] _4291;
    wire _4300;
    wire _4298;
    wire _4301;
    wire [63:0] _4305;
    wire _4296;
    wire _4294;
    wire _4297;
    wire [63:0] _4306;
    wire [63:0] _291;
    reg [63:0] _4304;
    wire _4313;
    wire _4311;
    wire _4314;
    wire [63:0] _4318;
    wire _4309;
    wire _4307;
    wire _4310;
    wire [63:0] _4319;
    wire [63:0] _292;
    reg [63:0] _4317;
    wire _4326;
    wire _4324;
    wire _4327;
    wire [63:0] _4331;
    wire _4322;
    wire _4320;
    wire _4323;
    wire [63:0] _4332;
    wire [63:0] _293;
    reg [63:0] _4330;
    wire _4339;
    wire _4337;
    wire _4340;
    wire [63:0] _4344;
    wire _4335;
    wire _4333;
    wire _4336;
    wire [63:0] _4345;
    wire [63:0] _294;
    reg [63:0] _4343;
    wire _4352;
    wire _4350;
    wire _4353;
    wire [63:0] _4357;
    wire _4348;
    wire _4346;
    wire _4349;
    wire [63:0] _4358;
    wire [63:0] _295;
    reg [63:0] _4356;
    wire _4365;
    wire _4363;
    wire _4366;
    wire [63:0] _4370;
    wire _4361;
    wire _4359;
    wire _4362;
    wire [63:0] _4371;
    wire [63:0] _296;
    reg [63:0] _4369;
    wire _4378;
    wire _4376;
    wire _4379;
    wire [63:0] _4383;
    wire _4374;
    wire _4372;
    wire _4375;
    wire [63:0] _4384;
    wire [63:0] _297;
    reg [63:0] _4382;
    wire _4391;
    wire _4389;
    wire _4392;
    wire [63:0] _4396;
    wire _4387;
    wire _4385;
    wire _4388;
    wire [63:0] _4397;
    wire [63:0] _298;
    reg [63:0] _4395;
    wire _4404;
    wire _4402;
    wire _4405;
    wire [63:0] _4409;
    wire _4400;
    wire _4398;
    wire _4401;
    wire [63:0] _4410;
    wire [63:0] _299;
    reg [63:0] _4408;
    wire _4417;
    wire _4415;
    wire _4418;
    wire [63:0] _4422;
    wire _4413;
    wire _4411;
    wire _4414;
    wire [63:0] _4423;
    wire [63:0] _300;
    reg [63:0] _4421;
    wire _4430;
    wire _4428;
    wire _4431;
    wire [63:0] _4435;
    wire _4426;
    wire _4424;
    wire _4427;
    wire [63:0] _4436;
    wire [63:0] _301;
    reg [63:0] _4434;
    wire _4443;
    wire _4441;
    wire _4444;
    wire [63:0] _4448;
    wire _4439;
    wire _4437;
    wire _4440;
    wire [63:0] _4449;
    wire [63:0] _302;
    reg [63:0] _4447;
    wire _4456;
    wire _4454;
    wire _4457;
    wire [63:0] _4461;
    wire _4452;
    wire _4450;
    wire _4453;
    wire [63:0] _4462;
    wire [63:0] _303;
    reg [63:0] _4460;
    wire _4469;
    wire _4467;
    wire _4470;
    wire [63:0] _4474;
    wire _4465;
    wire _4463;
    wire _4466;
    wire [63:0] _4475;
    wire [63:0] _304;
    reg [63:0] _4473;
    wire _4482;
    wire _4480;
    wire _4483;
    wire [63:0] _4487;
    wire _4478;
    wire _4476;
    wire _4479;
    wire [63:0] _4488;
    wire [63:0] _305;
    reg [63:0] _4486;
    wire _4495;
    wire _4493;
    wire _4496;
    wire [63:0] _4500;
    wire _4491;
    wire _4489;
    wire _4492;
    wire [63:0] _4501;
    wire [63:0] _306;
    reg [63:0] _4499;
    wire _4508;
    wire _4506;
    wire _4509;
    wire [63:0] _4513;
    wire _4504;
    wire _4502;
    wire _4505;
    wire [63:0] _4514;
    wire [63:0] _307;
    reg [63:0] _4512;
    wire _4521;
    wire _4519;
    wire _4522;
    wire [63:0] _4526;
    wire _4517;
    wire _4515;
    wire _4518;
    wire [63:0] _4527;
    wire [63:0] _308;
    reg [63:0] _4525;
    wire _4534;
    wire _4532;
    wire _4535;
    wire [63:0] _4539;
    wire _4530;
    wire _4528;
    wire _4531;
    wire [63:0] _4540;
    wire [63:0] _309;
    reg [63:0] _4538;
    wire _4547;
    wire _4545;
    wire _4548;
    wire [63:0] _4552;
    wire _4543;
    wire _4541;
    wire _4544;
    wire [63:0] _4553;
    wire [63:0] _310;
    reg [63:0] _4551;
    wire _4560;
    wire _4558;
    wire _4561;
    wire [63:0] _4565;
    wire _4556;
    wire _4554;
    wire _4557;
    wire [63:0] _4566;
    wire [63:0] _311;
    reg [63:0] _4564;
    wire _4573;
    wire _4571;
    wire _4574;
    wire [63:0] _4578;
    wire _4569;
    wire _4567;
    wire _4570;
    wire [63:0] _4579;
    wire [63:0] _312;
    reg [63:0] _4577;
    wire _4586;
    wire _4584;
    wire _4587;
    wire [63:0] _4591;
    wire _4582;
    wire _4580;
    wire _4583;
    wire [63:0] _4592;
    wire [63:0] _313;
    reg [63:0] _4590;
    wire _4599;
    wire _4597;
    wire _4600;
    wire [63:0] _4604;
    wire _4595;
    wire _4593;
    wire _4596;
    wire [63:0] _4605;
    wire [63:0] _314;
    reg [63:0] _4603;
    wire _4612;
    wire _4610;
    wire _4613;
    wire [63:0] _4617;
    wire _4608;
    wire _4606;
    wire _4609;
    wire [63:0] _4618;
    wire [63:0] _315;
    reg [63:0] _4616;
    wire _4625;
    wire _4623;
    wire _4626;
    wire [63:0] _4630;
    wire _4621;
    wire _4619;
    wire _4622;
    wire [63:0] _4631;
    wire [63:0] _316;
    reg [63:0] _4629;
    wire _4638;
    wire _4636;
    wire _4639;
    wire [63:0] _4643;
    wire _4634;
    wire _4632;
    wire _4635;
    wire [63:0] _4644;
    wire [63:0] _317;
    reg [63:0] _4642;
    wire _4651;
    wire _4649;
    wire _4652;
    wire [63:0] _4656;
    wire _4647;
    wire _4645;
    wire _4648;
    wire [63:0] _4657;
    wire [63:0] _318;
    reg [63:0] _4655;
    wire _4664;
    wire _4662;
    wire _4665;
    wire [63:0] _4669;
    wire _4660;
    wire _4658;
    wire _4661;
    wire [63:0] _4670;
    wire [63:0] _319;
    reg [63:0] _4668;
    wire _4677;
    wire _4675;
    wire _4678;
    wire [63:0] _4682;
    wire _4673;
    wire _4671;
    wire _4674;
    wire [63:0] _4683;
    wire [63:0] _320;
    reg [63:0] _4681;
    wire _4690;
    wire _4688;
    wire _4691;
    wire [63:0] _4695;
    wire _4686;
    wire _4684;
    wire _4687;
    wire [63:0] _4696;
    wire [63:0] _321;
    reg [63:0] _4694;
    wire _4703;
    wire _4701;
    wire _4704;
    wire [63:0] _4708;
    wire _4699;
    wire _4697;
    wire _4700;
    wire [63:0] _4709;
    wire [63:0] _322;
    reg [63:0] _4707;
    wire _4716;
    wire _4714;
    wire _4717;
    wire [63:0] _4721;
    wire _4712;
    wire _4710;
    wire _4713;
    wire [63:0] _4722;
    wire [63:0] _323;
    reg [63:0] _4720;
    wire _4729;
    wire _4727;
    wire _4730;
    wire [63:0] _4734;
    wire _4725;
    wire _4723;
    wire _4726;
    wire [63:0] _4735;
    wire [63:0] _324;
    reg [63:0] _4733;
    wire _4742;
    wire _4740;
    wire _4743;
    wire [63:0] _4747;
    wire _4738;
    wire _4736;
    wire _4739;
    wire [63:0] _4748;
    wire [63:0] _325;
    reg [63:0] _4746;
    wire _4755;
    wire _4753;
    wire _4756;
    wire [63:0] _4760;
    wire _4751;
    wire _4749;
    wire _4752;
    wire [63:0] _4761;
    wire [63:0] _326;
    reg [63:0] _4759;
    wire _4768;
    wire _4766;
    wire _4769;
    wire [63:0] _4773;
    wire _4764;
    wire _4762;
    wire _4765;
    wire [63:0] _4774;
    wire [63:0] _327;
    reg [63:0] _4772;
    wire _4781;
    wire _4779;
    wire _4782;
    wire [63:0] _4786;
    wire _4777;
    wire _4775;
    wire _4778;
    wire [63:0] _4787;
    wire [63:0] _328;
    reg [63:0] _4785;
    wire _4794;
    wire _4792;
    wire _4795;
    wire [63:0] _4799;
    wire _4790;
    wire _4788;
    wire _4791;
    wire [63:0] _4800;
    wire [63:0] _329;
    reg [63:0] _4798;
    wire _4807;
    wire _4805;
    wire _4808;
    wire [63:0] _4812;
    wire _4803;
    wire _4801;
    wire _4804;
    wire [63:0] _4813;
    wire [63:0] _330;
    reg [63:0] _4811;
    wire _4820;
    wire _4818;
    wire _4821;
    wire [63:0] _4825;
    wire _4816;
    wire _4814;
    wire _4817;
    wire [63:0] _4826;
    wire [63:0] _331;
    reg [63:0] _4824;
    wire _4833;
    wire _4831;
    wire _4834;
    wire [63:0] _4838;
    wire _4829;
    wire _4827;
    wire _4830;
    wire [63:0] _4839;
    wire [63:0] _332;
    reg [63:0] _4837;
    wire _4846;
    wire _4844;
    wire _4847;
    wire [63:0] _4851;
    wire _4842;
    wire _4840;
    wire _4843;
    wire [63:0] _4852;
    wire [63:0] _333;
    reg [63:0] _4850;
    wire _4859;
    wire _4857;
    wire _4860;
    wire [63:0] _4864;
    wire _4855;
    wire _4853;
    wire _4856;
    wire [63:0] _4865;
    wire [63:0] _334;
    reg [63:0] _4863;
    wire _4872;
    wire _4870;
    wire _4873;
    wire [63:0] _4877;
    wire _4868;
    wire _4866;
    wire _4869;
    wire [63:0] _4878;
    wire [63:0] _335;
    reg [63:0] _4876;
    wire _4885;
    wire _4883;
    wire _4886;
    wire [63:0] _4890;
    wire _4881;
    wire _4879;
    wire _4882;
    wire [63:0] _4891;
    wire [63:0] _336;
    reg [63:0] _4889;
    wire _4898;
    wire _4896;
    wire _4899;
    wire [63:0] _4903;
    wire _4894;
    wire _4892;
    wire _4895;
    wire [63:0] _4904;
    wire [63:0] _337;
    reg [63:0] _4902;
    wire _4911;
    wire _4909;
    wire _4912;
    wire [63:0] _4916;
    wire _4907;
    wire _4905;
    wire _4908;
    wire [63:0] _4917;
    wire [63:0] _338;
    reg [63:0] _4915;
    wire _4924;
    wire _4922;
    wire _4925;
    wire [63:0] _4929;
    wire _4920;
    wire _4918;
    wire _4921;
    wire [63:0] _4930;
    wire [63:0] _339;
    reg [63:0] _4928;
    wire _4937;
    wire _4935;
    wire _4938;
    wire [63:0] _4942;
    wire _4933;
    wire _4931;
    wire _4934;
    wire [63:0] _4943;
    wire [63:0] _340;
    reg [63:0] _4941;
    wire _4950;
    wire _4948;
    wire _4951;
    wire [63:0] _4955;
    wire _4946;
    wire _4944;
    wire _4947;
    wire [63:0] _4956;
    wire [63:0] _341;
    reg [63:0] _4954;
    wire _4963;
    wire _4961;
    wire _4964;
    wire [63:0] _4968;
    wire _4959;
    wire _4957;
    wire _4960;
    wire [63:0] _4969;
    wire [63:0] _342;
    reg [63:0] _4967;
    wire _4976;
    wire _4974;
    wire _4977;
    wire [63:0] _4981;
    wire _4972;
    wire _4970;
    wire _4973;
    wire [63:0] _4982;
    wire [63:0] _343;
    reg [63:0] _4980;
    wire _4989;
    wire _4987;
    wire _4990;
    wire [63:0] _4994;
    wire _4985;
    wire _4983;
    wire _4986;
    wire [63:0] _4995;
    wire [63:0] _344;
    reg [63:0] _4993;
    wire _5002;
    wire _5000;
    wire _5003;
    wire [63:0] _5007;
    wire _4998;
    wire _4996;
    wire _4999;
    wire [63:0] _5008;
    wire [63:0] _345;
    reg [63:0] _5006;
    wire _5015;
    wire _5013;
    wire _5016;
    wire [63:0] _5020;
    wire _5011;
    wire _5009;
    wire _5012;
    wire [63:0] _5021;
    wire [63:0] _346;
    reg [63:0] _5019;
    wire _5028;
    wire _5026;
    wire _5029;
    wire [63:0] _5033;
    wire _5024;
    wire _5022;
    wire _5025;
    wire [63:0] _5034;
    wire [63:0] _347;
    reg [63:0] _5032;
    wire _5041;
    wire _5039;
    wire _5042;
    wire [63:0] _5046;
    wire _5037;
    wire _5035;
    wire _5038;
    wire [63:0] _5047;
    wire [63:0] _348;
    reg [63:0] _5045;
    wire _5054;
    wire _5052;
    wire _5055;
    wire [63:0] _5059;
    wire _5050;
    wire _5048;
    wire _5051;
    wire [63:0] _5060;
    wire [63:0] _349;
    reg [63:0] _5058;
    wire _5067;
    wire _5065;
    wire _5068;
    wire [63:0] _5072;
    wire _5063;
    wire _5061;
    wire _5064;
    wire [63:0] _5073;
    wire [63:0] _350;
    reg [63:0] _5071;
    wire _5080;
    wire _5078;
    wire _5081;
    wire [63:0] _5085;
    wire _5076;
    wire _5074;
    wire _5077;
    wire [63:0] _5086;
    wire [63:0] _351;
    reg [63:0] _5084;
    wire _5093;
    wire _5091;
    wire _5094;
    wire [63:0] _5098;
    wire _5089;
    wire _5087;
    wire _5090;
    wire [63:0] _5099;
    wire [63:0] _352;
    reg [63:0] _5097;
    wire _5106;
    wire _5104;
    wire _5107;
    wire [63:0] _5111;
    wire _5102;
    wire _5100;
    wire _5103;
    wire [63:0] _5112;
    wire [63:0] _353;
    reg [63:0] _5110;
    wire _5119;
    wire _5117;
    wire _5120;
    wire [63:0] _5124;
    wire _5115;
    wire _5113;
    wire _5116;
    wire [63:0] _5125;
    wire [63:0] _354;
    reg [63:0] _5123;
    wire _5132;
    wire _5130;
    wire _5133;
    wire [63:0] _5137;
    wire _5128;
    wire _5126;
    wire _5129;
    wire [63:0] _5138;
    wire [63:0] _355;
    reg [63:0] _5136;
    wire _5145;
    wire _5143;
    wire _5146;
    wire [63:0] _5150;
    wire _5141;
    wire _5139;
    wire _5142;
    wire [63:0] _5151;
    wire [63:0] _356;
    reg [63:0] _5149;
    wire _5158;
    wire _5156;
    wire _5159;
    wire [63:0] _5163;
    wire _5154;
    wire _5152;
    wire _5155;
    wire [63:0] _5164;
    wire [63:0] _357;
    reg [63:0] _5162;
    wire _5171;
    wire _5169;
    wire _5172;
    wire [63:0] _5176;
    wire _5167;
    wire _5165;
    wire _5168;
    wire [63:0] _5177;
    wire [63:0] _358;
    reg [63:0] _5175;
    wire _5184;
    wire _5182;
    wire _5185;
    wire [63:0] _5189;
    wire _5180;
    wire _5178;
    wire _5181;
    wire [63:0] _5190;
    wire [63:0] _359;
    reg [63:0] _5188;
    wire _5197;
    wire _5195;
    wire _5198;
    wire [63:0] _5202;
    wire _5193;
    wire _5191;
    wire _5194;
    wire [63:0] _5203;
    wire [63:0] _360;
    reg [63:0] _5201;
    wire _5210;
    wire _5208;
    wire _5211;
    wire [63:0] _5215;
    wire _5206;
    wire _5204;
    wire _5207;
    wire [63:0] _5216;
    wire [63:0] _361;
    reg [63:0] _5214;
    wire _5223;
    wire _5221;
    wire _5224;
    wire [63:0] _5228;
    wire _5219;
    wire _5217;
    wire _5220;
    wire [63:0] _5229;
    wire [63:0] _362;
    reg [63:0] _5227;
    wire _5236;
    wire _5234;
    wire _5237;
    wire [63:0] _5241;
    wire _5232;
    wire _5230;
    wire _5233;
    wire [63:0] _5242;
    wire [63:0] _363;
    reg [63:0] _5240;
    wire _5249;
    wire _5247;
    wire _5250;
    wire [63:0] _5254;
    wire _5245;
    wire _5243;
    wire _5246;
    wire [63:0] _5255;
    wire [63:0] _364;
    reg [63:0] _5253;
    wire _5262;
    wire _5260;
    wire _5263;
    wire [63:0] _5267;
    wire _5258;
    wire _5256;
    wire _5259;
    wire [63:0] _5268;
    wire [63:0] _365;
    reg [63:0] _5266;
    wire _5275;
    wire _5273;
    wire _5276;
    wire [63:0] _5280;
    wire _5271;
    wire _5269;
    wire _5272;
    wire [63:0] _5281;
    wire [63:0] _366;
    reg [63:0] _5279;
    wire _5288;
    wire _5286;
    wire _5289;
    wire [63:0] _5293;
    wire _5284;
    wire _5282;
    wire _5285;
    wire [63:0] _5294;
    wire [63:0] _367;
    reg [63:0] _5292;
    wire _5301;
    wire _5299;
    wire _5302;
    wire [63:0] _5306;
    wire _5297;
    wire _5295;
    wire _5298;
    wire [63:0] _5307;
    wire [63:0] _368;
    reg [63:0] _5305;
    wire _5314;
    wire _5312;
    wire _5315;
    wire [63:0] _5319;
    wire _5310;
    wire _5308;
    wire _5311;
    wire [63:0] _5320;
    wire [63:0] _369;
    reg [63:0] _5318;
    wire _5327;
    wire _5325;
    wire _5328;
    wire [63:0] _5332;
    wire _5323;
    wire _5321;
    wire _5324;
    wire [63:0] _5333;
    wire [63:0] _370;
    reg [63:0] _5331;
    wire _5340;
    wire _5338;
    wire _5341;
    wire [63:0] _5345;
    wire _5336;
    wire _5334;
    wire _5337;
    wire [63:0] _5346;
    wire [63:0] _371;
    reg [63:0] _5344;
    wire _5353;
    wire _5351;
    wire _5354;
    wire [63:0] _5358;
    wire _5349;
    wire _5347;
    wire _5350;
    wire [63:0] _5359;
    wire [63:0] _372;
    reg [63:0] _5357;
    wire _5366;
    wire _5364;
    wire _5367;
    wire [63:0] _5371;
    wire _5362;
    wire _5360;
    wire _5363;
    wire [63:0] _5372;
    wire [63:0] _373;
    reg [63:0] _5370;
    wire _5379;
    wire _5377;
    wire _5380;
    wire [63:0] _5384;
    wire _5375;
    wire _5373;
    wire _5376;
    wire [63:0] _5385;
    wire [63:0] _374;
    reg [63:0] _5383;
    wire _5392;
    wire _5390;
    wire _5393;
    wire [63:0] _5397;
    wire _5388;
    wire _5386;
    wire _5389;
    wire [63:0] _5398;
    wire [63:0] _375;
    reg [63:0] _5396;
    wire _5405;
    wire _5403;
    wire _5406;
    wire [63:0] _5410;
    wire _5401;
    wire _5399;
    wire _5402;
    wire [63:0] _5411;
    wire [63:0] _376;
    reg [63:0] _5409;
    wire _5418;
    wire _5416;
    wire _5419;
    wire [63:0] _5423;
    wire _5414;
    wire _5412;
    wire _5415;
    wire [63:0] _5424;
    wire [63:0] _377;
    reg [63:0] _5422;
    wire _5431;
    wire _5429;
    wire _5432;
    wire [63:0] _5436;
    wire _5427;
    wire _5425;
    wire _5428;
    wire [63:0] _5437;
    wire [63:0] _378;
    reg [63:0] _5435;
    wire _5444;
    wire _5442;
    wire _5445;
    wire [63:0] _5449;
    wire _5440;
    wire _5438;
    wire _5441;
    wire [63:0] _5450;
    wire [63:0] _379;
    reg [63:0] _5448;
    wire _5457;
    wire _5455;
    wire _5458;
    wire [63:0] _5462;
    wire _5453;
    wire _5451;
    wire _5454;
    wire [63:0] _5463;
    wire [63:0] _380;
    reg [63:0] _5461;
    wire _5470;
    wire _5468;
    wire _5471;
    wire [63:0] _5475;
    wire _5466;
    wire _5464;
    wire _5467;
    wire [63:0] _5476;
    wire [63:0] _381;
    reg [63:0] _5474;
    wire _5483;
    wire _5481;
    wire _5484;
    wire [63:0] _5488;
    wire _5479;
    wire _5477;
    wire _5480;
    wire [63:0] _5489;
    wire [63:0] _382;
    reg [63:0] _5487;
    wire _5496;
    wire _5494;
    wire _5497;
    wire [63:0] _5501;
    wire _5492;
    wire _5490;
    wire _5493;
    wire [63:0] _5502;
    wire [63:0] _383;
    reg [63:0] _5500;
    wire _5509;
    wire _5507;
    wire _5510;
    wire [63:0] _5514;
    wire _5505;
    wire _5503;
    wire _5506;
    wire [63:0] _5515;
    wire [63:0] _384;
    reg [63:0] _5513;
    wire _5522;
    wire _5520;
    wire _5523;
    wire [63:0] _5527;
    wire _5518;
    wire _5516;
    wire _5519;
    wire [63:0] _5528;
    wire [63:0] _385;
    reg [63:0] _5526;
    wire _5535;
    wire _5533;
    wire _5536;
    wire [63:0] _5540;
    wire _5531;
    wire _5529;
    wire _5532;
    wire [63:0] _5541;
    wire [63:0] _386;
    reg [63:0] _5539;
    wire _5548;
    wire _5546;
    wire _5549;
    wire [63:0] _5553;
    wire _5544;
    wire _5542;
    wire _5545;
    wire [63:0] _5554;
    wire [63:0] _387;
    reg [63:0] _5552;
    wire _5561;
    wire _5559;
    wire _5562;
    wire [63:0] _5566;
    wire _5557;
    wire _5555;
    wire _5558;
    wire [63:0] _5567;
    wire [63:0] _388;
    reg [63:0] _5565;
    wire _5574;
    wire _5572;
    wire _5575;
    wire [63:0] _5579;
    wire _5570;
    wire _5568;
    wire _5571;
    wire [63:0] _5580;
    wire [63:0] _389;
    reg [63:0] _5578;
    wire _5587;
    wire _5585;
    wire _5588;
    wire [63:0] _5592;
    wire _5583;
    wire _5581;
    wire _5584;
    wire [63:0] _5593;
    wire [63:0] _390;
    reg [63:0] _5591;
    wire _5600;
    wire _5598;
    wire _5601;
    wire [63:0] _5605;
    wire _5596;
    wire _5594;
    wire _5597;
    wire [63:0] _5606;
    wire [63:0] _391;
    reg [63:0] _5604;
    wire _5613;
    wire _5611;
    wire _5614;
    wire [63:0] _5618;
    wire _5609;
    wire _5607;
    wire _5610;
    wire [63:0] _5619;
    wire [63:0] _392;
    reg [63:0] _5617;
    wire _5626;
    wire _5624;
    wire _5627;
    wire [63:0] _5631;
    wire _5622;
    wire _5620;
    wire _5623;
    wire [63:0] _5632;
    wire [63:0] _393;
    reg [63:0] _5630;
    wire _5639;
    wire _5637;
    wire _5640;
    wire [63:0] _5644;
    wire _5635;
    wire _5633;
    wire _5636;
    wire [63:0] _5645;
    wire [63:0] _394;
    reg [63:0] _5643;
    wire _5652;
    wire _5650;
    wire _5653;
    wire [63:0] _5657;
    wire _5648;
    wire _5646;
    wire _5649;
    wire [63:0] _5658;
    wire [63:0] _395;
    reg [63:0] _5656;
    wire _5665;
    wire _5663;
    wire _5666;
    wire [63:0] _5670;
    wire _5661;
    wire _5659;
    wire _5662;
    wire [63:0] _5671;
    wire [63:0] _396;
    reg [63:0] _5669;
    wire _5678;
    wire _5676;
    wire _5679;
    wire [63:0] _5683;
    wire _5674;
    wire _5672;
    wire _5675;
    wire [63:0] _5684;
    wire [63:0] _397;
    reg [63:0] _5682;
    wire _5691;
    wire _5689;
    wire _5692;
    wire [63:0] _5696;
    wire _5687;
    wire _5685;
    wire _5688;
    wire [63:0] _5697;
    wire [63:0] _398;
    reg [63:0] _5695;
    wire _5704;
    wire _5702;
    wire _5705;
    wire [63:0] _5709;
    wire _5700;
    wire _5698;
    wire _5701;
    wire [63:0] _5710;
    wire [63:0] _399;
    reg [63:0] _5708;
    wire _5717;
    wire _5715;
    wire _5718;
    wire [63:0] _5722;
    wire _5713;
    wire _5711;
    wire _5714;
    wire [63:0] _5723;
    wire [63:0] _400;
    reg [63:0] _5721;
    wire _5730;
    wire _5728;
    wire _5731;
    wire [63:0] _5735;
    wire _5726;
    wire _5724;
    wire _5727;
    wire [63:0] _5736;
    wire [63:0] _401;
    reg [63:0] _5734;
    wire _5743;
    wire _5741;
    wire _5744;
    wire [63:0] _5748;
    wire _5739;
    wire _5737;
    wire _5740;
    wire [63:0] _5749;
    wire [63:0] _402;
    reg [63:0] _5747;
    wire _5756;
    wire _5754;
    wire _5757;
    wire [63:0] _5761;
    wire _5752;
    wire _5750;
    wire _5753;
    wire [63:0] _5762;
    wire [63:0] _403;
    reg [63:0] _5760;
    wire _5769;
    wire _5767;
    wire _5770;
    wire [63:0] _5774;
    wire _5765;
    wire _5763;
    wire _5766;
    wire [63:0] _5775;
    wire [63:0] _404;
    reg [63:0] _5773;
    wire _5782;
    wire _5780;
    wire _5783;
    wire [63:0] _5787;
    wire _5778;
    wire _5776;
    wire _5779;
    wire [63:0] _5788;
    wire [63:0] _405;
    reg [63:0] _5786;
    wire _5795;
    wire _5793;
    wire _5796;
    wire [63:0] _5800;
    wire _5791;
    wire _5789;
    wire _5792;
    wire [63:0] _5801;
    wire [63:0] _406;
    reg [63:0] _5799;
    wire _5808;
    wire _5806;
    wire _5809;
    wire [63:0] _5813;
    wire _5804;
    wire _5802;
    wire _5805;
    wire [63:0] _5814;
    wire [63:0] _407;
    reg [63:0] _5812;
    wire _5821;
    wire _5819;
    wire _5822;
    wire [63:0] _5826;
    wire _5817;
    wire _5815;
    wire _5818;
    wire [63:0] _5827;
    wire [63:0] _408;
    reg [63:0] _5825;
    wire _5834;
    wire _5832;
    wire _5835;
    wire [63:0] _5839;
    wire _5830;
    wire _5828;
    wire _5831;
    wire [63:0] _5840;
    wire [63:0] _409;
    reg [63:0] _5838;
    wire _5847;
    wire _5845;
    wire _5848;
    wire [63:0] _5852;
    wire _5843;
    wire _5841;
    wire _5844;
    wire [63:0] _5853;
    wire [63:0] _410;
    reg [63:0] _5851;
    wire _5860;
    wire _5858;
    wire _5861;
    wire [63:0] _5865;
    wire _5856;
    wire _5854;
    wire _5857;
    wire [63:0] _5866;
    wire [63:0] _411;
    reg [63:0] _5864;
    wire _5873;
    wire _5871;
    wire _5874;
    wire [63:0] _5878;
    wire _5869;
    wire _5867;
    wire _5870;
    wire [63:0] _5879;
    wire [63:0] _412;
    reg [63:0] _5877;
    wire _5886;
    wire _5884;
    wire _5887;
    wire [63:0] _5891;
    wire _5882;
    wire _5880;
    wire _5883;
    wire [63:0] _5892;
    wire [63:0] _413;
    reg [63:0] _5890;
    wire _5899;
    wire _5897;
    wire _5900;
    wire [63:0] _5904;
    wire _5895;
    wire _5893;
    wire _5896;
    wire [63:0] _5905;
    wire [63:0] _414;
    reg [63:0] _5903;
    wire _5912;
    wire _5910;
    wire _5913;
    wire [63:0] _5917;
    wire _5908;
    wire _5906;
    wire _5909;
    wire [63:0] _5918;
    wire [63:0] _415;
    reg [63:0] _5916;
    wire _5925;
    wire _5923;
    wire _5926;
    wire [63:0] _5930;
    wire _5921;
    wire _5919;
    wire _5922;
    wire [63:0] _5931;
    wire [63:0] _416;
    reg [63:0] _5929;
    wire _5938;
    wire _5936;
    wire _5939;
    wire [63:0] _5943;
    wire _5934;
    wire _5932;
    wire _5935;
    wire [63:0] _5944;
    wire [63:0] _417;
    reg [63:0] _5942;
    wire _5951;
    wire _5949;
    wire _5952;
    wire [63:0] _5956;
    wire _5947;
    wire _5945;
    wire _5948;
    wire [63:0] _5957;
    wire [63:0] _418;
    reg [63:0] _5955;
    wire _5964;
    wire _5962;
    wire _5965;
    wire [63:0] _5969;
    wire _5960;
    wire _5958;
    wire _5961;
    wire [63:0] _5970;
    wire [63:0] _419;
    reg [63:0] _5968;
    wire _5977;
    wire _5975;
    wire _5978;
    wire [63:0] _5982;
    wire _5973;
    wire _5971;
    wire _5974;
    wire [63:0] _5983;
    wire [63:0] _420;
    reg [63:0] _5981;
    wire _5990;
    wire _5988;
    wire _5991;
    wire [63:0] _5995;
    wire _5986;
    wire _5984;
    wire _5987;
    wire [63:0] _5996;
    wire [63:0] _421;
    reg [63:0] _5994;
    wire _6003;
    wire _6001;
    wire _6004;
    wire [63:0] _6008;
    wire _5999;
    wire _5997;
    wire _6000;
    wire [63:0] _6009;
    wire [63:0] _422;
    reg [63:0] _6007;
    wire _6016;
    wire _6014;
    wire _6017;
    wire [63:0] _6021;
    wire _6012;
    wire _6010;
    wire _6013;
    wire [63:0] _6022;
    wire [63:0] _423;
    reg [63:0] _6020;
    wire _6029;
    wire _6027;
    wire _6030;
    wire [63:0] _6034;
    wire _6025;
    wire _6023;
    wire _6026;
    wire [63:0] _6035;
    wire [63:0] _424;
    reg [63:0] _6033;
    wire _6042;
    wire _6040;
    wire _6043;
    wire [63:0] _6047;
    wire _6038;
    wire _6036;
    wire _6039;
    wire [63:0] _6048;
    wire [63:0] _425;
    reg [63:0] _6046;
    wire _6055;
    wire _6053;
    wire _6056;
    wire [63:0] _6060;
    wire _6051;
    wire _6049;
    wire _6052;
    wire [63:0] _6061;
    wire [63:0] _426;
    reg [63:0] _6059;
    wire _6068;
    wire _6066;
    wire _6069;
    wire [63:0] _6073;
    wire _6064;
    wire _6062;
    wire _6065;
    wire [63:0] _6074;
    wire [63:0] _427;
    reg [63:0] _6072;
    wire _6081;
    wire _6079;
    wire _6082;
    wire [63:0] _6086;
    wire _6077;
    wire _6075;
    wire _6078;
    wire [63:0] _6087;
    wire [63:0] _428;
    reg [63:0] _6085;
    wire _6094;
    wire _6092;
    wire _6095;
    wire [63:0] _6099;
    wire _6090;
    wire _6088;
    wire _6091;
    wire [63:0] _6100;
    wire [63:0] _429;
    reg [63:0] _6098;
    wire _6107;
    wire _6105;
    wire _6108;
    wire [63:0] _6112;
    wire _6103;
    wire _6101;
    wire _6104;
    wire [63:0] _6113;
    wire [63:0] _430;
    reg [63:0] _6111;
    wire _6120;
    wire _6118;
    wire _6121;
    wire [63:0] _6125;
    wire _6116;
    wire _6114;
    wire _6117;
    wire [63:0] _6126;
    wire [63:0] _431;
    reg [63:0] _6124;
    wire _6133;
    wire _6131;
    wire _6134;
    wire [63:0] _6138;
    wire _6129;
    wire _6127;
    wire _6130;
    wire [63:0] _6139;
    wire [63:0] _432;
    reg [63:0] _6137;
    wire _6146;
    wire _6144;
    wire _6147;
    wire [63:0] _6151;
    wire _6142;
    wire _6140;
    wire _6143;
    wire [63:0] _6152;
    wire [63:0] _433;
    reg [63:0] _6150;
    wire _6159;
    wire _6157;
    wire _6160;
    wire [63:0] _6164;
    wire _6155;
    wire _6153;
    wire _6156;
    wire [63:0] _6165;
    wire [63:0] _434;
    reg [63:0] _6163;
    wire _6172;
    wire _6170;
    wire _6173;
    wire [63:0] _6177;
    wire _6168;
    wire _6166;
    wire _6169;
    wire [63:0] _6178;
    wire [63:0] _435;
    reg [63:0] _6176;
    wire _6185;
    wire _6183;
    wire _6186;
    wire [63:0] _6190;
    wire _6181;
    wire _6179;
    wire _6182;
    wire [63:0] _6191;
    wire [63:0] _436;
    reg [63:0] _6189;
    wire _6198;
    wire _6196;
    wire _6199;
    wire [63:0] _6203;
    wire _6194;
    wire _6192;
    wire _6195;
    wire [63:0] _6204;
    wire [63:0] _437;
    reg [63:0] _6202;
    wire _6211;
    wire _6209;
    wire _6212;
    wire [63:0] _6216;
    wire _6207;
    wire _6205;
    wire _6208;
    wire [63:0] _6217;
    wire [63:0] _438;
    reg [63:0] _6215;
    wire _6224;
    wire _6222;
    wire _6225;
    wire [63:0] _6229;
    wire _6220;
    wire _6218;
    wire _6221;
    wire [63:0] _6230;
    wire [63:0] _439;
    reg [63:0] _6228;
    wire _6237;
    wire _6235;
    wire _6238;
    wire [63:0] _6242;
    wire _6233;
    wire _6231;
    wire _6234;
    wire [63:0] _6243;
    wire [63:0] _440;
    reg [63:0] _6241;
    wire _6250;
    wire _6248;
    wire _6251;
    wire [63:0] _6255;
    wire _6246;
    wire _6244;
    wire _6247;
    wire [63:0] _6256;
    wire [63:0] _441;
    reg [63:0] _6254;
    wire _6263;
    wire _6261;
    wire _6264;
    wire [63:0] _6268;
    wire _6259;
    wire _6257;
    wire _6260;
    wire [63:0] _6269;
    wire [63:0] _442;
    reg [63:0] _6267;
    wire _6276;
    wire _6274;
    wire _6277;
    wire [63:0] _6281;
    wire _6272;
    wire _6270;
    wire _6273;
    wire [63:0] _6282;
    wire [63:0] _443;
    reg [63:0] _6280;
    wire _6289;
    wire _6287;
    wire _6290;
    wire [63:0] _6294;
    wire _6285;
    wire _6283;
    wire _6286;
    wire [63:0] _6295;
    wire [63:0] _444;
    reg [63:0] _6293;
    wire _6302;
    wire _6300;
    wire _6303;
    wire [63:0] _6307;
    wire _6298;
    wire _6296;
    wire _6299;
    wire [63:0] _6308;
    wire [63:0] _445;
    reg [63:0] _6306;
    wire _6315;
    wire _6313;
    wire _6316;
    wire [63:0] _6320;
    wire _6311;
    wire _6309;
    wire _6312;
    wire [63:0] _6321;
    wire [63:0] _446;
    reg [63:0] _6319;
    wire _6328;
    wire _6326;
    wire _6329;
    wire [63:0] _6333;
    wire _6324;
    wire _6322;
    wire _6325;
    wire [63:0] _6334;
    wire [63:0] _447;
    reg [63:0] _6332;
    wire _6341;
    wire _6339;
    wire _6342;
    wire [63:0] _6346;
    wire _6337;
    wire _6335;
    wire _6338;
    wire [63:0] _6347;
    wire [63:0] _448;
    reg [63:0] _6345;
    wire _6354;
    wire _6352;
    wire _6355;
    wire [63:0] _6359;
    wire _6350;
    wire _6348;
    wire _6351;
    wire [63:0] _6360;
    wire [63:0] _449;
    reg [63:0] _6358;
    wire _6367;
    wire _6365;
    wire _6368;
    wire [63:0] _6372;
    wire _6363;
    wire _6361;
    wire _6364;
    wire [63:0] _6373;
    wire [63:0] _450;
    reg [63:0] _6371;
    wire _6380;
    wire _6378;
    wire _6381;
    wire [63:0] _6385;
    wire _6376;
    wire _6374;
    wire _6377;
    wire [63:0] _6386;
    wire [63:0] _451;
    reg [63:0] _6384;
    wire _6393;
    wire _6391;
    wire _6394;
    wire [63:0] _6398;
    wire _6389;
    wire _6387;
    wire _6390;
    wire [63:0] _6399;
    wire [63:0] _452;
    reg [63:0] _6397;
    wire _6406;
    wire _6404;
    wire _6407;
    wire [63:0] _6411;
    wire _6402;
    wire _6400;
    wire _6403;
    wire [63:0] _6412;
    wire [63:0] _453;
    reg [63:0] _6410;
    wire _6419;
    wire _6417;
    wire _6420;
    wire [63:0] _6424;
    wire _6415;
    wire _6413;
    wire _6416;
    wire [63:0] _6425;
    wire [63:0] _454;
    reg [63:0] _6423;
    wire _6432;
    wire _6430;
    wire _6433;
    wire [63:0] _6437;
    wire _6428;
    wire _6426;
    wire _6429;
    wire [63:0] _6438;
    wire [63:0] _455;
    reg [63:0] _6436;
    wire _6445;
    wire _6443;
    wire _6446;
    wire [63:0] _6450;
    wire _6441;
    wire _6439;
    wire _6442;
    wire [63:0] _6451;
    wire [63:0] _456;
    reg [63:0] _6449;
    wire _6458;
    wire _6456;
    wire _6459;
    wire [63:0] _6463;
    wire _6454;
    wire _6452;
    wire _6455;
    wire [63:0] _6464;
    wire [63:0] _457;
    reg [63:0] _6462;
    wire _6471;
    wire _6469;
    wire _6472;
    wire [63:0] _6476;
    wire _6467;
    wire _6465;
    wire _6468;
    wire [63:0] _6477;
    wire [63:0] _458;
    reg [63:0] _6475;
    wire _6484;
    wire _6482;
    wire _6485;
    wire [63:0] _6489;
    wire _6480;
    wire _6478;
    wire _6481;
    wire [63:0] _6490;
    wire [63:0] _459;
    reg [63:0] _6488;
    wire _6497;
    wire _6495;
    wire _6498;
    wire [63:0] _6502;
    wire _6493;
    wire _6491;
    wire _6494;
    wire [63:0] _6503;
    wire [63:0] _460;
    reg [63:0] _6501;
    wire _6510;
    wire _6508;
    wire _6511;
    wire [63:0] _6515;
    wire _6506;
    wire _6504;
    wire _6507;
    wire [63:0] _6516;
    wire [63:0] _461;
    reg [63:0] _6514;
    wire _6523;
    wire _6521;
    wire _6524;
    wire [63:0] _6528;
    wire _6519;
    wire _6517;
    wire _6520;
    wire [63:0] _6529;
    wire [63:0] _462;
    reg [63:0] _6527;
    wire _6536;
    wire _6534;
    wire _6537;
    wire [63:0] _6541;
    wire _6532;
    wire _6530;
    wire _6533;
    wire [63:0] _6542;
    wire [63:0] _463;
    reg [63:0] _6540;
    wire _6549;
    wire _6547;
    wire _6550;
    wire [63:0] _6554;
    wire _6545;
    wire _6543;
    wire _6546;
    wire [63:0] _6555;
    wire [63:0] _464;
    reg [63:0] _6553;
    wire _6562;
    wire _6560;
    wire _6563;
    wire [63:0] _6567;
    wire _6558;
    wire _6556;
    wire _6559;
    wire [63:0] _6568;
    wire [63:0] _465;
    reg [63:0] _6566;
    wire _6575;
    wire _6573;
    wire _6576;
    wire [63:0] _6580;
    wire _6571;
    wire _6569;
    wire _6572;
    wire [63:0] _6581;
    wire [63:0] _466;
    reg [63:0] _6579;
    wire _6588;
    wire _6586;
    wire _6589;
    wire [63:0] _6593;
    wire _6584;
    wire _6582;
    wire _6585;
    wire [63:0] _6594;
    wire [63:0] _467;
    reg [63:0] _6592;
    wire _6601;
    wire _6599;
    wire _6602;
    wire [63:0] _6606;
    wire _6597;
    wire _6595;
    wire _6598;
    wire [63:0] _6607;
    wire [63:0] _468;
    reg [63:0] _6605;
    wire _6614;
    wire _6612;
    wire _6615;
    wire [63:0] _6619;
    wire _6610;
    wire _6608;
    wire _6611;
    wire [63:0] _6620;
    wire [63:0] _469;
    reg [63:0] _6618;
    wire _6627;
    wire _6625;
    wire _6628;
    wire [63:0] _6632;
    wire _6623;
    wire _6621;
    wire _6624;
    wire [63:0] _6633;
    wire [63:0] _470;
    reg [63:0] _6631;
    wire _6640;
    wire _6638;
    wire _6641;
    wire [63:0] _6645;
    wire _6636;
    wire _6634;
    wire _6637;
    wire [63:0] _6646;
    wire [63:0] _471;
    reg [63:0] _6644;
    wire _6653;
    wire _6651;
    wire _6654;
    wire [63:0] _6658;
    wire _6649;
    wire _6647;
    wire _6650;
    wire [63:0] _6659;
    wire [63:0] _472;
    reg [63:0] _6657;
    wire _6666;
    wire _6664;
    wire _6667;
    wire [63:0] _6671;
    wire _6662;
    wire _6660;
    wire _6663;
    wire [63:0] _6672;
    wire [63:0] _473;
    reg [63:0] _6670;
    wire _6679;
    wire _6677;
    wire _6680;
    wire [63:0] _6684;
    wire _6675;
    wire _6673;
    wire _6676;
    wire [63:0] _6685;
    wire [63:0] _474;
    reg [63:0] _6683;
    wire _6692;
    wire _6690;
    wire _6693;
    wire [63:0] _6697;
    wire _6688;
    wire _6686;
    wire _6689;
    wire [63:0] _6698;
    wire [63:0] _475;
    reg [63:0] _6696;
    wire _6705;
    wire _6703;
    wire _6706;
    wire [63:0] _6710;
    wire _6701;
    wire _6699;
    wire _6702;
    wire [63:0] _6711;
    wire [63:0] _476;
    reg [63:0] _6709;
    wire _6718;
    wire _6716;
    wire _6719;
    wire [63:0] _6723;
    wire _6714;
    wire _6712;
    wire _6715;
    wire [63:0] _6724;
    wire [63:0] _477;
    reg [63:0] _6722;
    wire _6731;
    wire _6729;
    wire _6732;
    wire [63:0] _6736;
    wire _6727;
    wire _6725;
    wire _6728;
    wire [63:0] _6737;
    wire [63:0] _478;
    reg [63:0] _6735;
    wire _6744;
    wire _6742;
    wire _6745;
    wire [63:0] _6749;
    wire _6740;
    wire _6738;
    wire _6741;
    wire [63:0] _6750;
    wire [63:0] _479;
    reg [63:0] _6748;
    wire _6757;
    wire _6755;
    wire _6758;
    wire [63:0] _6762;
    wire _6753;
    wire _6751;
    wire _6754;
    wire [63:0] _6763;
    wire [63:0] _480;
    reg [63:0] _6761;
    wire _6770;
    wire _6768;
    wire _6771;
    wire [63:0] _6775;
    wire _6766;
    wire _6764;
    wire _6767;
    wire [63:0] _6776;
    wire [63:0] _481;
    reg [63:0] _6774;
    wire _6783;
    wire _6781;
    wire _6784;
    wire [63:0] _6788;
    wire _6779;
    wire _6777;
    wire _6780;
    wire [63:0] _6789;
    wire [63:0] _482;
    reg [63:0] _6787;
    wire _6796;
    wire _6794;
    wire _6797;
    wire [63:0] _6801;
    wire _6792;
    wire _6790;
    wire _6793;
    wire [63:0] _6802;
    wire [63:0] _483;
    reg [63:0] _6800;
    wire _6809;
    wire _6807;
    wire _6810;
    wire [63:0] _6814;
    wire _6805;
    wire _6803;
    wire _6806;
    wire [63:0] _6815;
    wire [63:0] _484;
    reg [63:0] _6813;
    wire _6822;
    wire _6820;
    wire _6823;
    wire [63:0] _6827;
    wire _6818;
    wire _6816;
    wire _6819;
    wire [63:0] _6828;
    wire [63:0] _485;
    reg [63:0] _6826;
    wire _6835;
    wire _6833;
    wire _6836;
    wire [63:0] _6840;
    wire _6831;
    wire _6829;
    wire _6832;
    wire [63:0] _6841;
    wire [63:0] _486;
    reg [63:0] _6839;
    wire _6848;
    wire _6846;
    wire _6849;
    wire [63:0] _6853;
    wire _6844;
    wire _6842;
    wire _6845;
    wire [63:0] _6854;
    wire [63:0] _487;
    reg [63:0] _6852;
    wire _6861;
    wire _6859;
    wire _6862;
    wire [63:0] _6866;
    wire _6857;
    wire _6855;
    wire _6858;
    wire [63:0] _6867;
    wire [63:0] _488;
    reg [63:0] _6865;
    wire _6874;
    wire _6872;
    wire _6875;
    wire [63:0] _6879;
    wire _6870;
    wire _6868;
    wire _6871;
    wire [63:0] _6880;
    wire [63:0] _489;
    reg [63:0] _6878;
    wire _6887;
    wire _6885;
    wire _6888;
    wire [63:0] _6892;
    wire _6883;
    wire _6881;
    wire _6884;
    wire [63:0] _6893;
    wire [63:0] _490;
    reg [63:0] _6891;
    wire _6900;
    wire _6898;
    wire _6901;
    wire [63:0] _6905;
    wire _6896;
    wire _6894;
    wire _6897;
    wire [63:0] _6906;
    wire [63:0] _491;
    reg [63:0] _6904;
    wire _6913;
    wire _6911;
    wire _6914;
    wire [63:0] _6918;
    wire _6909;
    wire _6907;
    wire _6910;
    wire [63:0] _6919;
    wire [63:0] _492;
    reg [63:0] _6917;
    wire _6926;
    wire _6924;
    wire _6927;
    wire [63:0] _6931;
    wire _6922;
    wire _6920;
    wire _6923;
    wire [63:0] _6932;
    wire [63:0] _493;
    reg [63:0] _6930;
    wire _6939;
    wire _6937;
    wire _6940;
    wire [63:0] _6944;
    wire _6935;
    wire _6933;
    wire _6936;
    wire [63:0] _6945;
    wire [63:0] _494;
    reg [63:0] _6943;
    wire _6952;
    wire _6950;
    wire _6953;
    wire [63:0] _6957;
    wire _6948;
    wire _6946;
    wire _6949;
    wire [63:0] _6958;
    wire [63:0] _495;
    reg [63:0] _6956;
    wire _6965;
    wire _6963;
    wire _6966;
    wire [63:0] _6970;
    wire _6961;
    wire _6959;
    wire _6962;
    wire [63:0] _6971;
    wire [63:0] _496;
    reg [63:0] _6969;
    wire _6978;
    wire _6976;
    wire _6979;
    wire [63:0] _6983;
    wire _6974;
    wire _6972;
    wire _6975;
    wire [63:0] _6984;
    wire [63:0] _497;
    reg [63:0] _6982;
    wire _6991;
    wire _6989;
    wire _6992;
    wire [63:0] _6996;
    wire _6987;
    wire _6985;
    wire _6988;
    wire [63:0] _6997;
    wire [63:0] _498;
    reg [63:0] _6995;
    wire _7004;
    wire _7002;
    wire _7005;
    wire [63:0] _7009;
    wire _7000;
    wire _6998;
    wire _7001;
    wire [63:0] _7010;
    wire [63:0] _499;
    reg [63:0] _7008;
    wire _7017;
    wire _7015;
    wire _7018;
    wire [63:0] _7022;
    wire _7013;
    wire _7011;
    wire _7014;
    wire [63:0] _7023;
    wire [63:0] _500;
    reg [63:0] _7021;
    wire _7030;
    wire _7028;
    wire _7031;
    wire [63:0] _7035;
    wire _7026;
    wire _7024;
    wire _7027;
    wire [63:0] _7036;
    wire [63:0] _501;
    reg [63:0] _7034;
    wire _7043;
    wire _7041;
    wire _7044;
    wire [63:0] _7048;
    wire _7039;
    wire _7037;
    wire _7040;
    wire [63:0] _7049;
    wire [63:0] _502;
    reg [63:0] _7047;
    wire _7056;
    wire _7054;
    wire _7057;
    wire [63:0] _7061;
    wire _7052;
    wire _7050;
    wire _7053;
    wire [63:0] _7062;
    wire [63:0] _503;
    reg [63:0] _7060;
    wire _7069;
    wire _7067;
    wire _7070;
    wire [63:0] _7074;
    wire _7065;
    wire _7063;
    wire _7066;
    wire [63:0] _7075;
    wire [63:0] _504;
    reg [63:0] _7073;
    wire _7082;
    wire _7080;
    wire _7083;
    wire [63:0] _7087;
    wire _7078;
    wire _7076;
    wire _7079;
    wire [63:0] _7088;
    wire [63:0] _505;
    reg [63:0] _7086;
    wire _7095;
    wire _7093;
    wire _7096;
    wire [63:0] _7100;
    wire _7091;
    wire _7089;
    wire _7092;
    wire [63:0] _7101;
    wire [63:0] _506;
    reg [63:0] _7099;
    wire _7108;
    wire _7106;
    wire _7109;
    wire [63:0] _7113;
    wire _7104;
    wire _7102;
    wire _7105;
    wire [63:0] _7114;
    wire [63:0] _507;
    reg [63:0] _7112;
    wire _7121;
    wire _7119;
    wire _7122;
    wire [63:0] _7126;
    wire _7117;
    wire _7115;
    wire _7118;
    wire [63:0] _7127;
    wire [63:0] _508;
    reg [63:0] _7125;
    wire _7134;
    wire _7132;
    wire _7135;
    wire [63:0] _7139;
    wire _7130;
    wire _7128;
    wire _7131;
    wire [63:0] _7140;
    wire [63:0] _509;
    reg [63:0] _7138;
    wire _7147;
    wire _7145;
    wire _7148;
    wire [63:0] _7152;
    wire _7143;
    wire _7141;
    wire _7144;
    wire [63:0] _7153;
    wire [63:0] _510;
    reg [63:0] _7151;
    wire _7160;
    wire _7158;
    wire _7161;
    wire [63:0] _7165;
    wire _7156;
    wire _7154;
    wire _7157;
    wire [63:0] _7166;
    wire [63:0] _511;
    reg [63:0] _7164;
    wire _7173;
    wire _7171;
    wire _7174;
    wire [63:0] _7178;
    wire _7169;
    wire _7167;
    wire _7170;
    wire [63:0] _7179;
    wire [63:0] _512;
    reg [63:0] _7177;
    wire _7186;
    wire _7184;
    wire _7187;
    wire [63:0] _7191;
    wire _7182;
    wire _7180;
    wire _7183;
    wire [63:0] _7192;
    wire [63:0] _513;
    reg [63:0] _7190;
    wire _7199;
    wire _7197;
    wire _7200;
    wire [63:0] _7204;
    wire _7195;
    wire _7193;
    wire _7196;
    wire [63:0] _7205;
    wire [63:0] _514;
    reg [63:0] _7203;
    wire _7212;
    wire _7210;
    wire _7213;
    wire [63:0] _7217;
    wire _7208;
    wire _7206;
    wire _7209;
    wire [63:0] _7218;
    wire [63:0] _515;
    reg [63:0] _7216;
    wire _7225;
    wire _7223;
    wire _7226;
    wire [63:0] _7230;
    wire _7221;
    wire _7219;
    wire _7222;
    wire [63:0] _7231;
    wire [63:0] _516;
    reg [63:0] _7229;
    wire _7238;
    wire _7236;
    wire _7239;
    wire [63:0] _7243;
    wire _7234;
    wire _7232;
    wire _7235;
    wire [63:0] _7244;
    wire [63:0] _517;
    reg [63:0] _7242;
    wire _7251;
    wire _7249;
    wire _7252;
    wire [63:0] _7256;
    wire _7247;
    wire _7245;
    wire _7248;
    wire [63:0] _7257;
    wire [63:0] _518;
    reg [63:0] _7255;
    wire _7264;
    wire _7262;
    wire _7265;
    wire [63:0] _7269;
    wire _7260;
    wire _7258;
    wire _7261;
    wire [63:0] _7270;
    wire [63:0] _519;
    reg [63:0] _7268;
    wire [7:0] _7297;
    wire [7:0] _7298;
    wire _7271;
    wire [7:0] _7300;
    wire [7:0] _7302;
    wire [7:0] _520;
    reg [7:0] _7285;
    reg [63:0] _7286;
    wire [63:0] _522;
    wire [63:0] _7304;
    wire [63:0] _7306;
    wire [63:0] _523;
    reg [63:0] _7282;
    wire _7287;
    wire _7288;
    wire [7:0] _7308;
    wire [7:0] _615;
    wire [7:0] _7310;
    wire [7:0] _7312;
    wire [7:0] _524;
    reg [7:0] _609;
    wire _594;
    wire [63:0] _595;
    wire [63:0] _526;
    wire [63:0] _592;
    wire [63:0] _593;
    wire _589;
    wire _590;
    wire [63:0] _596;
    wire _587;
    wire _588;
    wire [63:0] _597;
    wire [63:0] _7313;
    wire [63:0] _7315;
    wire [63:0] _527;
    reg [63:0] _577;
    wire [63:0] _529;
    wire _578;
    wire _579;
    wire _572;
    wire _7316;
    wire _7317;
    wire _7319;
    wire _530;
    reg _573;
    wire _574;
    wire _580;
    wire [7:0] _616;
    wire [7:0] _7309;
    wire _7320;
    wire [7:0] _7321;
    wire [7:0] _7323;
    wire [7:0] _531;
    reg [7:0] _7275;
    wire _7277;
    wire _7278;
    wire _7272;
    wire _7279;
    wire _7289;
    wire _7295;
    wire _7325;
    wire [1:0] _552;
    wire [1:0] _557;
    wire [1:0] _555;
    wire _533;
    wire _535;
    wire _537;
    wire _539;
    wire vdd;
    wire _7328;
    wire _7329;
    wire _7331;
    wire _540;
    reg _561;
    wire _562;
    wire _563;
    wire _7303;
    wire _7335;
    wire _7337;
    wire _541;
    reg _7334;
    wire _7339;
    wire [1:0] _7340;
    wire _543;
    wire _545;
    wire _569;
    wire _570;
    wire _565;
    wire _7338;
    wire [1:0] _7341;
    wire [1:0] _7342;
    wire [1:0] _546;
    reg [1:0] _554;
    wire _558;
    wire _7324;
    wire _7326;
    wire _7349;
    wire [63:0] _7355;
    wire _548;
    wire [63:0] _7357;
    wire [63:0] _549;
    reg [63:0] _7352;
    assign _556 = _554 == _555;
    assign _567 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign _600 = _597 - _599;
    assign _601 = _586 + _600;
    assign _584 = _577 - _583;
    assign _585 = _568 + _584;
    assign _586 = _580 ? _585 : _568;
    assign _602 = _570 ? _601 : _586;
    assign _603 = _565 ? _602 : _568;
    assign _605 = _548 ? _567 : _603;
    assign _5 = _605;
    always @(posedge _539) begin
        if (_537)
            _568 <= _567;
        else
            _568 <= _5;
    end
    assign _7353 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    assign _7354 = _7352 + _7353;
    assign _7347 = _7282 < _7286;
    assign _617 = 8'b11111111;
    assign _618 = _616 == _617;
    assign _613 = _565 & _570;
    assign _619 = _613 & _618;
    assign _623 = _619 ? _599 : _622;
    assign _611 = _609 == _617;
    assign _606 = _565 & _580;
    assign _612 = _606 & _611;
    assign _624 = _612 ? _583 : _623;
    assign _7 = _624;
    always @(posedge _539) begin
        if (_537)
            _622 <= _567;
        else
            _622 <= _7;
    end
    assign _630 = 8'b11111110;
    assign _631 = _616 == _630;
    assign _629 = _565 & _570;
    assign _632 = _629 & _631;
    assign _636 = _632 ? _599 : _635;
    assign _627 = _609 == _630;
    assign _625 = _565 & _580;
    assign _628 = _625 & _627;
    assign _637 = _628 ? _583 : _636;
    assign _8 = _637;
    always @(posedge _539) begin
        if (_537)
            _635 <= _567;
        else
            _635 <= _8;
    end
    assign _643 = 8'b11111101;
    assign _644 = _616 == _643;
    assign _642 = _565 & _570;
    assign _645 = _642 & _644;
    assign _649 = _645 ? _599 : _648;
    assign _640 = _609 == _643;
    assign _638 = _565 & _580;
    assign _641 = _638 & _640;
    assign _650 = _641 ? _583 : _649;
    assign _9 = _650;
    always @(posedge _539) begin
        if (_537)
            _648 <= _567;
        else
            _648 <= _9;
    end
    assign _656 = 8'b11111100;
    assign _657 = _616 == _656;
    assign _655 = _565 & _570;
    assign _658 = _655 & _657;
    assign _662 = _658 ? _599 : _661;
    assign _653 = _609 == _656;
    assign _651 = _565 & _580;
    assign _654 = _651 & _653;
    assign _663 = _654 ? _583 : _662;
    assign _10 = _663;
    always @(posedge _539) begin
        if (_537)
            _661 <= _567;
        else
            _661 <= _10;
    end
    assign _669 = 8'b11111011;
    assign _670 = _616 == _669;
    assign _668 = _565 & _570;
    assign _671 = _668 & _670;
    assign _675 = _671 ? _599 : _674;
    assign _666 = _609 == _669;
    assign _664 = _565 & _580;
    assign _667 = _664 & _666;
    assign _676 = _667 ? _583 : _675;
    assign _11 = _676;
    always @(posedge _539) begin
        if (_537)
            _674 <= _567;
        else
            _674 <= _11;
    end
    assign _682 = 8'b11111010;
    assign _683 = _616 == _682;
    assign _681 = _565 & _570;
    assign _684 = _681 & _683;
    assign _688 = _684 ? _599 : _687;
    assign _679 = _609 == _682;
    assign _677 = _565 & _580;
    assign _680 = _677 & _679;
    assign _689 = _680 ? _583 : _688;
    assign _12 = _689;
    always @(posedge _539) begin
        if (_537)
            _687 <= _567;
        else
            _687 <= _12;
    end
    assign _695 = 8'b11111001;
    assign _696 = _616 == _695;
    assign _694 = _565 & _570;
    assign _697 = _694 & _696;
    assign _701 = _697 ? _599 : _700;
    assign _692 = _609 == _695;
    assign _690 = _565 & _580;
    assign _693 = _690 & _692;
    assign _702 = _693 ? _583 : _701;
    assign _13 = _702;
    always @(posedge _539) begin
        if (_537)
            _700 <= _567;
        else
            _700 <= _13;
    end
    assign _708 = 8'b11111000;
    assign _709 = _616 == _708;
    assign _707 = _565 & _570;
    assign _710 = _707 & _709;
    assign _714 = _710 ? _599 : _713;
    assign _705 = _609 == _708;
    assign _703 = _565 & _580;
    assign _706 = _703 & _705;
    assign _715 = _706 ? _583 : _714;
    assign _14 = _715;
    always @(posedge _539) begin
        if (_537)
            _713 <= _567;
        else
            _713 <= _14;
    end
    assign _721 = 8'b11110111;
    assign _722 = _616 == _721;
    assign _720 = _565 & _570;
    assign _723 = _720 & _722;
    assign _727 = _723 ? _599 : _726;
    assign _718 = _609 == _721;
    assign _716 = _565 & _580;
    assign _719 = _716 & _718;
    assign _728 = _719 ? _583 : _727;
    assign _15 = _728;
    always @(posedge _539) begin
        if (_537)
            _726 <= _567;
        else
            _726 <= _15;
    end
    assign _734 = 8'b11110110;
    assign _735 = _616 == _734;
    assign _733 = _565 & _570;
    assign _736 = _733 & _735;
    assign _740 = _736 ? _599 : _739;
    assign _731 = _609 == _734;
    assign _729 = _565 & _580;
    assign _732 = _729 & _731;
    assign _741 = _732 ? _583 : _740;
    assign _16 = _741;
    always @(posedge _539) begin
        if (_537)
            _739 <= _567;
        else
            _739 <= _16;
    end
    assign _747 = 8'b11110101;
    assign _748 = _616 == _747;
    assign _746 = _565 & _570;
    assign _749 = _746 & _748;
    assign _753 = _749 ? _599 : _752;
    assign _744 = _609 == _747;
    assign _742 = _565 & _580;
    assign _745 = _742 & _744;
    assign _754 = _745 ? _583 : _753;
    assign _17 = _754;
    always @(posedge _539) begin
        if (_537)
            _752 <= _567;
        else
            _752 <= _17;
    end
    assign _760 = 8'b11110100;
    assign _761 = _616 == _760;
    assign _759 = _565 & _570;
    assign _762 = _759 & _761;
    assign _766 = _762 ? _599 : _765;
    assign _757 = _609 == _760;
    assign _755 = _565 & _580;
    assign _758 = _755 & _757;
    assign _767 = _758 ? _583 : _766;
    assign _18 = _767;
    always @(posedge _539) begin
        if (_537)
            _765 <= _567;
        else
            _765 <= _18;
    end
    assign _773 = 8'b11110011;
    assign _774 = _616 == _773;
    assign _772 = _565 & _570;
    assign _775 = _772 & _774;
    assign _779 = _775 ? _599 : _778;
    assign _770 = _609 == _773;
    assign _768 = _565 & _580;
    assign _771 = _768 & _770;
    assign _780 = _771 ? _583 : _779;
    assign _19 = _780;
    always @(posedge _539) begin
        if (_537)
            _778 <= _567;
        else
            _778 <= _19;
    end
    assign _786 = 8'b11110010;
    assign _787 = _616 == _786;
    assign _785 = _565 & _570;
    assign _788 = _785 & _787;
    assign _792 = _788 ? _599 : _791;
    assign _783 = _609 == _786;
    assign _781 = _565 & _580;
    assign _784 = _781 & _783;
    assign _793 = _784 ? _583 : _792;
    assign _20 = _793;
    always @(posedge _539) begin
        if (_537)
            _791 <= _567;
        else
            _791 <= _20;
    end
    assign _799 = 8'b11110001;
    assign _800 = _616 == _799;
    assign _798 = _565 & _570;
    assign _801 = _798 & _800;
    assign _805 = _801 ? _599 : _804;
    assign _796 = _609 == _799;
    assign _794 = _565 & _580;
    assign _797 = _794 & _796;
    assign _806 = _797 ? _583 : _805;
    assign _21 = _806;
    always @(posedge _539) begin
        if (_537)
            _804 <= _567;
        else
            _804 <= _21;
    end
    assign _812 = 8'b11110000;
    assign _813 = _616 == _812;
    assign _811 = _565 & _570;
    assign _814 = _811 & _813;
    assign _818 = _814 ? _599 : _817;
    assign _809 = _609 == _812;
    assign _807 = _565 & _580;
    assign _810 = _807 & _809;
    assign _819 = _810 ? _583 : _818;
    assign _22 = _819;
    always @(posedge _539) begin
        if (_537)
            _817 <= _567;
        else
            _817 <= _22;
    end
    assign _825 = 8'b11101111;
    assign _826 = _616 == _825;
    assign _824 = _565 & _570;
    assign _827 = _824 & _826;
    assign _831 = _827 ? _599 : _830;
    assign _822 = _609 == _825;
    assign _820 = _565 & _580;
    assign _823 = _820 & _822;
    assign _832 = _823 ? _583 : _831;
    assign _23 = _832;
    always @(posedge _539) begin
        if (_537)
            _830 <= _567;
        else
            _830 <= _23;
    end
    assign _838 = 8'b11101110;
    assign _839 = _616 == _838;
    assign _837 = _565 & _570;
    assign _840 = _837 & _839;
    assign _844 = _840 ? _599 : _843;
    assign _835 = _609 == _838;
    assign _833 = _565 & _580;
    assign _836 = _833 & _835;
    assign _845 = _836 ? _583 : _844;
    assign _24 = _845;
    always @(posedge _539) begin
        if (_537)
            _843 <= _567;
        else
            _843 <= _24;
    end
    assign _851 = 8'b11101101;
    assign _852 = _616 == _851;
    assign _850 = _565 & _570;
    assign _853 = _850 & _852;
    assign _857 = _853 ? _599 : _856;
    assign _848 = _609 == _851;
    assign _846 = _565 & _580;
    assign _849 = _846 & _848;
    assign _858 = _849 ? _583 : _857;
    assign _25 = _858;
    always @(posedge _539) begin
        if (_537)
            _856 <= _567;
        else
            _856 <= _25;
    end
    assign _864 = 8'b11101100;
    assign _865 = _616 == _864;
    assign _863 = _565 & _570;
    assign _866 = _863 & _865;
    assign _870 = _866 ? _599 : _869;
    assign _861 = _609 == _864;
    assign _859 = _565 & _580;
    assign _862 = _859 & _861;
    assign _871 = _862 ? _583 : _870;
    assign _26 = _871;
    always @(posedge _539) begin
        if (_537)
            _869 <= _567;
        else
            _869 <= _26;
    end
    assign _877 = 8'b11101011;
    assign _878 = _616 == _877;
    assign _876 = _565 & _570;
    assign _879 = _876 & _878;
    assign _883 = _879 ? _599 : _882;
    assign _874 = _609 == _877;
    assign _872 = _565 & _580;
    assign _875 = _872 & _874;
    assign _884 = _875 ? _583 : _883;
    assign _27 = _884;
    always @(posedge _539) begin
        if (_537)
            _882 <= _567;
        else
            _882 <= _27;
    end
    assign _890 = 8'b11101010;
    assign _891 = _616 == _890;
    assign _889 = _565 & _570;
    assign _892 = _889 & _891;
    assign _896 = _892 ? _599 : _895;
    assign _887 = _609 == _890;
    assign _885 = _565 & _580;
    assign _888 = _885 & _887;
    assign _897 = _888 ? _583 : _896;
    assign _28 = _897;
    always @(posedge _539) begin
        if (_537)
            _895 <= _567;
        else
            _895 <= _28;
    end
    assign _903 = 8'b11101001;
    assign _904 = _616 == _903;
    assign _902 = _565 & _570;
    assign _905 = _902 & _904;
    assign _909 = _905 ? _599 : _908;
    assign _900 = _609 == _903;
    assign _898 = _565 & _580;
    assign _901 = _898 & _900;
    assign _910 = _901 ? _583 : _909;
    assign _29 = _910;
    always @(posedge _539) begin
        if (_537)
            _908 <= _567;
        else
            _908 <= _29;
    end
    assign _916 = 8'b11101000;
    assign _917 = _616 == _916;
    assign _915 = _565 & _570;
    assign _918 = _915 & _917;
    assign _922 = _918 ? _599 : _921;
    assign _913 = _609 == _916;
    assign _911 = _565 & _580;
    assign _914 = _911 & _913;
    assign _923 = _914 ? _583 : _922;
    assign _30 = _923;
    always @(posedge _539) begin
        if (_537)
            _921 <= _567;
        else
            _921 <= _30;
    end
    assign _929 = 8'b11100111;
    assign _930 = _616 == _929;
    assign _928 = _565 & _570;
    assign _931 = _928 & _930;
    assign _935 = _931 ? _599 : _934;
    assign _926 = _609 == _929;
    assign _924 = _565 & _580;
    assign _927 = _924 & _926;
    assign _936 = _927 ? _583 : _935;
    assign _31 = _936;
    always @(posedge _539) begin
        if (_537)
            _934 <= _567;
        else
            _934 <= _31;
    end
    assign _942 = 8'b11100110;
    assign _943 = _616 == _942;
    assign _941 = _565 & _570;
    assign _944 = _941 & _943;
    assign _948 = _944 ? _599 : _947;
    assign _939 = _609 == _942;
    assign _937 = _565 & _580;
    assign _940 = _937 & _939;
    assign _949 = _940 ? _583 : _948;
    assign _32 = _949;
    always @(posedge _539) begin
        if (_537)
            _947 <= _567;
        else
            _947 <= _32;
    end
    assign _955 = 8'b11100101;
    assign _956 = _616 == _955;
    assign _954 = _565 & _570;
    assign _957 = _954 & _956;
    assign _961 = _957 ? _599 : _960;
    assign _952 = _609 == _955;
    assign _950 = _565 & _580;
    assign _953 = _950 & _952;
    assign _962 = _953 ? _583 : _961;
    assign _33 = _962;
    always @(posedge _539) begin
        if (_537)
            _960 <= _567;
        else
            _960 <= _33;
    end
    assign _968 = 8'b11100100;
    assign _969 = _616 == _968;
    assign _967 = _565 & _570;
    assign _970 = _967 & _969;
    assign _974 = _970 ? _599 : _973;
    assign _965 = _609 == _968;
    assign _963 = _565 & _580;
    assign _966 = _963 & _965;
    assign _975 = _966 ? _583 : _974;
    assign _34 = _975;
    always @(posedge _539) begin
        if (_537)
            _973 <= _567;
        else
            _973 <= _34;
    end
    assign _981 = 8'b11100011;
    assign _982 = _616 == _981;
    assign _980 = _565 & _570;
    assign _983 = _980 & _982;
    assign _987 = _983 ? _599 : _986;
    assign _978 = _609 == _981;
    assign _976 = _565 & _580;
    assign _979 = _976 & _978;
    assign _988 = _979 ? _583 : _987;
    assign _35 = _988;
    always @(posedge _539) begin
        if (_537)
            _986 <= _567;
        else
            _986 <= _35;
    end
    assign _994 = 8'b11100010;
    assign _995 = _616 == _994;
    assign _993 = _565 & _570;
    assign _996 = _993 & _995;
    assign _1000 = _996 ? _599 : _999;
    assign _991 = _609 == _994;
    assign _989 = _565 & _580;
    assign _992 = _989 & _991;
    assign _1001 = _992 ? _583 : _1000;
    assign _36 = _1001;
    always @(posedge _539) begin
        if (_537)
            _999 <= _567;
        else
            _999 <= _36;
    end
    assign _1007 = 8'b11100001;
    assign _1008 = _616 == _1007;
    assign _1006 = _565 & _570;
    assign _1009 = _1006 & _1008;
    assign _1013 = _1009 ? _599 : _1012;
    assign _1004 = _609 == _1007;
    assign _1002 = _565 & _580;
    assign _1005 = _1002 & _1004;
    assign _1014 = _1005 ? _583 : _1013;
    assign _37 = _1014;
    always @(posedge _539) begin
        if (_537)
            _1012 <= _567;
        else
            _1012 <= _37;
    end
    assign _1020 = 8'b11100000;
    assign _1021 = _616 == _1020;
    assign _1019 = _565 & _570;
    assign _1022 = _1019 & _1021;
    assign _1026 = _1022 ? _599 : _1025;
    assign _1017 = _609 == _1020;
    assign _1015 = _565 & _580;
    assign _1018 = _1015 & _1017;
    assign _1027 = _1018 ? _583 : _1026;
    assign _38 = _1027;
    always @(posedge _539) begin
        if (_537)
            _1025 <= _567;
        else
            _1025 <= _38;
    end
    assign _1033 = 8'b11011111;
    assign _1034 = _616 == _1033;
    assign _1032 = _565 & _570;
    assign _1035 = _1032 & _1034;
    assign _1039 = _1035 ? _599 : _1038;
    assign _1030 = _609 == _1033;
    assign _1028 = _565 & _580;
    assign _1031 = _1028 & _1030;
    assign _1040 = _1031 ? _583 : _1039;
    assign _39 = _1040;
    always @(posedge _539) begin
        if (_537)
            _1038 <= _567;
        else
            _1038 <= _39;
    end
    assign _1046 = 8'b11011110;
    assign _1047 = _616 == _1046;
    assign _1045 = _565 & _570;
    assign _1048 = _1045 & _1047;
    assign _1052 = _1048 ? _599 : _1051;
    assign _1043 = _609 == _1046;
    assign _1041 = _565 & _580;
    assign _1044 = _1041 & _1043;
    assign _1053 = _1044 ? _583 : _1052;
    assign _40 = _1053;
    always @(posedge _539) begin
        if (_537)
            _1051 <= _567;
        else
            _1051 <= _40;
    end
    assign _1059 = 8'b11011101;
    assign _1060 = _616 == _1059;
    assign _1058 = _565 & _570;
    assign _1061 = _1058 & _1060;
    assign _1065 = _1061 ? _599 : _1064;
    assign _1056 = _609 == _1059;
    assign _1054 = _565 & _580;
    assign _1057 = _1054 & _1056;
    assign _1066 = _1057 ? _583 : _1065;
    assign _41 = _1066;
    always @(posedge _539) begin
        if (_537)
            _1064 <= _567;
        else
            _1064 <= _41;
    end
    assign _1072 = 8'b11011100;
    assign _1073 = _616 == _1072;
    assign _1071 = _565 & _570;
    assign _1074 = _1071 & _1073;
    assign _1078 = _1074 ? _599 : _1077;
    assign _1069 = _609 == _1072;
    assign _1067 = _565 & _580;
    assign _1070 = _1067 & _1069;
    assign _1079 = _1070 ? _583 : _1078;
    assign _42 = _1079;
    always @(posedge _539) begin
        if (_537)
            _1077 <= _567;
        else
            _1077 <= _42;
    end
    assign _1085 = 8'b11011011;
    assign _1086 = _616 == _1085;
    assign _1084 = _565 & _570;
    assign _1087 = _1084 & _1086;
    assign _1091 = _1087 ? _599 : _1090;
    assign _1082 = _609 == _1085;
    assign _1080 = _565 & _580;
    assign _1083 = _1080 & _1082;
    assign _1092 = _1083 ? _583 : _1091;
    assign _43 = _1092;
    always @(posedge _539) begin
        if (_537)
            _1090 <= _567;
        else
            _1090 <= _43;
    end
    assign _1098 = 8'b11011010;
    assign _1099 = _616 == _1098;
    assign _1097 = _565 & _570;
    assign _1100 = _1097 & _1099;
    assign _1104 = _1100 ? _599 : _1103;
    assign _1095 = _609 == _1098;
    assign _1093 = _565 & _580;
    assign _1096 = _1093 & _1095;
    assign _1105 = _1096 ? _583 : _1104;
    assign _44 = _1105;
    always @(posedge _539) begin
        if (_537)
            _1103 <= _567;
        else
            _1103 <= _44;
    end
    assign _1111 = 8'b11011001;
    assign _1112 = _616 == _1111;
    assign _1110 = _565 & _570;
    assign _1113 = _1110 & _1112;
    assign _1117 = _1113 ? _599 : _1116;
    assign _1108 = _609 == _1111;
    assign _1106 = _565 & _580;
    assign _1109 = _1106 & _1108;
    assign _1118 = _1109 ? _583 : _1117;
    assign _45 = _1118;
    always @(posedge _539) begin
        if (_537)
            _1116 <= _567;
        else
            _1116 <= _45;
    end
    assign _1124 = 8'b11011000;
    assign _1125 = _616 == _1124;
    assign _1123 = _565 & _570;
    assign _1126 = _1123 & _1125;
    assign _1130 = _1126 ? _599 : _1129;
    assign _1121 = _609 == _1124;
    assign _1119 = _565 & _580;
    assign _1122 = _1119 & _1121;
    assign _1131 = _1122 ? _583 : _1130;
    assign _46 = _1131;
    always @(posedge _539) begin
        if (_537)
            _1129 <= _567;
        else
            _1129 <= _46;
    end
    assign _1137 = 8'b11010111;
    assign _1138 = _616 == _1137;
    assign _1136 = _565 & _570;
    assign _1139 = _1136 & _1138;
    assign _1143 = _1139 ? _599 : _1142;
    assign _1134 = _609 == _1137;
    assign _1132 = _565 & _580;
    assign _1135 = _1132 & _1134;
    assign _1144 = _1135 ? _583 : _1143;
    assign _47 = _1144;
    always @(posedge _539) begin
        if (_537)
            _1142 <= _567;
        else
            _1142 <= _47;
    end
    assign _1150 = 8'b11010110;
    assign _1151 = _616 == _1150;
    assign _1149 = _565 & _570;
    assign _1152 = _1149 & _1151;
    assign _1156 = _1152 ? _599 : _1155;
    assign _1147 = _609 == _1150;
    assign _1145 = _565 & _580;
    assign _1148 = _1145 & _1147;
    assign _1157 = _1148 ? _583 : _1156;
    assign _48 = _1157;
    always @(posedge _539) begin
        if (_537)
            _1155 <= _567;
        else
            _1155 <= _48;
    end
    assign _1163 = 8'b11010101;
    assign _1164 = _616 == _1163;
    assign _1162 = _565 & _570;
    assign _1165 = _1162 & _1164;
    assign _1169 = _1165 ? _599 : _1168;
    assign _1160 = _609 == _1163;
    assign _1158 = _565 & _580;
    assign _1161 = _1158 & _1160;
    assign _1170 = _1161 ? _583 : _1169;
    assign _49 = _1170;
    always @(posedge _539) begin
        if (_537)
            _1168 <= _567;
        else
            _1168 <= _49;
    end
    assign _1176 = 8'b11010100;
    assign _1177 = _616 == _1176;
    assign _1175 = _565 & _570;
    assign _1178 = _1175 & _1177;
    assign _1182 = _1178 ? _599 : _1181;
    assign _1173 = _609 == _1176;
    assign _1171 = _565 & _580;
    assign _1174 = _1171 & _1173;
    assign _1183 = _1174 ? _583 : _1182;
    assign _50 = _1183;
    always @(posedge _539) begin
        if (_537)
            _1181 <= _567;
        else
            _1181 <= _50;
    end
    assign _1189 = 8'b11010011;
    assign _1190 = _616 == _1189;
    assign _1188 = _565 & _570;
    assign _1191 = _1188 & _1190;
    assign _1195 = _1191 ? _599 : _1194;
    assign _1186 = _609 == _1189;
    assign _1184 = _565 & _580;
    assign _1187 = _1184 & _1186;
    assign _1196 = _1187 ? _583 : _1195;
    assign _51 = _1196;
    always @(posedge _539) begin
        if (_537)
            _1194 <= _567;
        else
            _1194 <= _51;
    end
    assign _1202 = 8'b11010010;
    assign _1203 = _616 == _1202;
    assign _1201 = _565 & _570;
    assign _1204 = _1201 & _1203;
    assign _1208 = _1204 ? _599 : _1207;
    assign _1199 = _609 == _1202;
    assign _1197 = _565 & _580;
    assign _1200 = _1197 & _1199;
    assign _1209 = _1200 ? _583 : _1208;
    assign _52 = _1209;
    always @(posedge _539) begin
        if (_537)
            _1207 <= _567;
        else
            _1207 <= _52;
    end
    assign _1215 = 8'b11010001;
    assign _1216 = _616 == _1215;
    assign _1214 = _565 & _570;
    assign _1217 = _1214 & _1216;
    assign _1221 = _1217 ? _599 : _1220;
    assign _1212 = _609 == _1215;
    assign _1210 = _565 & _580;
    assign _1213 = _1210 & _1212;
    assign _1222 = _1213 ? _583 : _1221;
    assign _53 = _1222;
    always @(posedge _539) begin
        if (_537)
            _1220 <= _567;
        else
            _1220 <= _53;
    end
    assign _1228 = 8'b11010000;
    assign _1229 = _616 == _1228;
    assign _1227 = _565 & _570;
    assign _1230 = _1227 & _1229;
    assign _1234 = _1230 ? _599 : _1233;
    assign _1225 = _609 == _1228;
    assign _1223 = _565 & _580;
    assign _1226 = _1223 & _1225;
    assign _1235 = _1226 ? _583 : _1234;
    assign _54 = _1235;
    always @(posedge _539) begin
        if (_537)
            _1233 <= _567;
        else
            _1233 <= _54;
    end
    assign _1241 = 8'b11001111;
    assign _1242 = _616 == _1241;
    assign _1240 = _565 & _570;
    assign _1243 = _1240 & _1242;
    assign _1247 = _1243 ? _599 : _1246;
    assign _1238 = _609 == _1241;
    assign _1236 = _565 & _580;
    assign _1239 = _1236 & _1238;
    assign _1248 = _1239 ? _583 : _1247;
    assign _55 = _1248;
    always @(posedge _539) begin
        if (_537)
            _1246 <= _567;
        else
            _1246 <= _55;
    end
    assign _1254 = 8'b11001110;
    assign _1255 = _616 == _1254;
    assign _1253 = _565 & _570;
    assign _1256 = _1253 & _1255;
    assign _1260 = _1256 ? _599 : _1259;
    assign _1251 = _609 == _1254;
    assign _1249 = _565 & _580;
    assign _1252 = _1249 & _1251;
    assign _1261 = _1252 ? _583 : _1260;
    assign _56 = _1261;
    always @(posedge _539) begin
        if (_537)
            _1259 <= _567;
        else
            _1259 <= _56;
    end
    assign _1267 = 8'b11001101;
    assign _1268 = _616 == _1267;
    assign _1266 = _565 & _570;
    assign _1269 = _1266 & _1268;
    assign _1273 = _1269 ? _599 : _1272;
    assign _1264 = _609 == _1267;
    assign _1262 = _565 & _580;
    assign _1265 = _1262 & _1264;
    assign _1274 = _1265 ? _583 : _1273;
    assign _57 = _1274;
    always @(posedge _539) begin
        if (_537)
            _1272 <= _567;
        else
            _1272 <= _57;
    end
    assign _1280 = 8'b11001100;
    assign _1281 = _616 == _1280;
    assign _1279 = _565 & _570;
    assign _1282 = _1279 & _1281;
    assign _1286 = _1282 ? _599 : _1285;
    assign _1277 = _609 == _1280;
    assign _1275 = _565 & _580;
    assign _1278 = _1275 & _1277;
    assign _1287 = _1278 ? _583 : _1286;
    assign _58 = _1287;
    always @(posedge _539) begin
        if (_537)
            _1285 <= _567;
        else
            _1285 <= _58;
    end
    assign _1293 = 8'b11001011;
    assign _1294 = _616 == _1293;
    assign _1292 = _565 & _570;
    assign _1295 = _1292 & _1294;
    assign _1299 = _1295 ? _599 : _1298;
    assign _1290 = _609 == _1293;
    assign _1288 = _565 & _580;
    assign _1291 = _1288 & _1290;
    assign _1300 = _1291 ? _583 : _1299;
    assign _59 = _1300;
    always @(posedge _539) begin
        if (_537)
            _1298 <= _567;
        else
            _1298 <= _59;
    end
    assign _1306 = 8'b11001010;
    assign _1307 = _616 == _1306;
    assign _1305 = _565 & _570;
    assign _1308 = _1305 & _1307;
    assign _1312 = _1308 ? _599 : _1311;
    assign _1303 = _609 == _1306;
    assign _1301 = _565 & _580;
    assign _1304 = _1301 & _1303;
    assign _1313 = _1304 ? _583 : _1312;
    assign _60 = _1313;
    always @(posedge _539) begin
        if (_537)
            _1311 <= _567;
        else
            _1311 <= _60;
    end
    assign _1319 = 8'b11001001;
    assign _1320 = _616 == _1319;
    assign _1318 = _565 & _570;
    assign _1321 = _1318 & _1320;
    assign _1325 = _1321 ? _599 : _1324;
    assign _1316 = _609 == _1319;
    assign _1314 = _565 & _580;
    assign _1317 = _1314 & _1316;
    assign _1326 = _1317 ? _583 : _1325;
    assign _61 = _1326;
    always @(posedge _539) begin
        if (_537)
            _1324 <= _567;
        else
            _1324 <= _61;
    end
    assign _1332 = 8'b11001000;
    assign _1333 = _616 == _1332;
    assign _1331 = _565 & _570;
    assign _1334 = _1331 & _1333;
    assign _1338 = _1334 ? _599 : _1337;
    assign _1329 = _609 == _1332;
    assign _1327 = _565 & _580;
    assign _1330 = _1327 & _1329;
    assign _1339 = _1330 ? _583 : _1338;
    assign _62 = _1339;
    always @(posedge _539) begin
        if (_537)
            _1337 <= _567;
        else
            _1337 <= _62;
    end
    assign _1345 = 8'b11000111;
    assign _1346 = _616 == _1345;
    assign _1344 = _565 & _570;
    assign _1347 = _1344 & _1346;
    assign _1351 = _1347 ? _599 : _1350;
    assign _1342 = _609 == _1345;
    assign _1340 = _565 & _580;
    assign _1343 = _1340 & _1342;
    assign _1352 = _1343 ? _583 : _1351;
    assign _63 = _1352;
    always @(posedge _539) begin
        if (_537)
            _1350 <= _567;
        else
            _1350 <= _63;
    end
    assign _1358 = 8'b11000110;
    assign _1359 = _616 == _1358;
    assign _1357 = _565 & _570;
    assign _1360 = _1357 & _1359;
    assign _1364 = _1360 ? _599 : _1363;
    assign _1355 = _609 == _1358;
    assign _1353 = _565 & _580;
    assign _1356 = _1353 & _1355;
    assign _1365 = _1356 ? _583 : _1364;
    assign _64 = _1365;
    always @(posedge _539) begin
        if (_537)
            _1363 <= _567;
        else
            _1363 <= _64;
    end
    assign _1371 = 8'b11000101;
    assign _1372 = _616 == _1371;
    assign _1370 = _565 & _570;
    assign _1373 = _1370 & _1372;
    assign _1377 = _1373 ? _599 : _1376;
    assign _1368 = _609 == _1371;
    assign _1366 = _565 & _580;
    assign _1369 = _1366 & _1368;
    assign _1378 = _1369 ? _583 : _1377;
    assign _65 = _1378;
    always @(posedge _539) begin
        if (_537)
            _1376 <= _567;
        else
            _1376 <= _65;
    end
    assign _1384 = 8'b11000100;
    assign _1385 = _616 == _1384;
    assign _1383 = _565 & _570;
    assign _1386 = _1383 & _1385;
    assign _1390 = _1386 ? _599 : _1389;
    assign _1381 = _609 == _1384;
    assign _1379 = _565 & _580;
    assign _1382 = _1379 & _1381;
    assign _1391 = _1382 ? _583 : _1390;
    assign _66 = _1391;
    always @(posedge _539) begin
        if (_537)
            _1389 <= _567;
        else
            _1389 <= _66;
    end
    assign _1397 = 8'b11000011;
    assign _1398 = _616 == _1397;
    assign _1396 = _565 & _570;
    assign _1399 = _1396 & _1398;
    assign _1403 = _1399 ? _599 : _1402;
    assign _1394 = _609 == _1397;
    assign _1392 = _565 & _580;
    assign _1395 = _1392 & _1394;
    assign _1404 = _1395 ? _583 : _1403;
    assign _67 = _1404;
    always @(posedge _539) begin
        if (_537)
            _1402 <= _567;
        else
            _1402 <= _67;
    end
    assign _1410 = 8'b11000010;
    assign _1411 = _616 == _1410;
    assign _1409 = _565 & _570;
    assign _1412 = _1409 & _1411;
    assign _1416 = _1412 ? _599 : _1415;
    assign _1407 = _609 == _1410;
    assign _1405 = _565 & _580;
    assign _1408 = _1405 & _1407;
    assign _1417 = _1408 ? _583 : _1416;
    assign _68 = _1417;
    always @(posedge _539) begin
        if (_537)
            _1415 <= _567;
        else
            _1415 <= _68;
    end
    assign _1423 = 8'b11000001;
    assign _1424 = _616 == _1423;
    assign _1422 = _565 & _570;
    assign _1425 = _1422 & _1424;
    assign _1429 = _1425 ? _599 : _1428;
    assign _1420 = _609 == _1423;
    assign _1418 = _565 & _580;
    assign _1421 = _1418 & _1420;
    assign _1430 = _1421 ? _583 : _1429;
    assign _69 = _1430;
    always @(posedge _539) begin
        if (_537)
            _1428 <= _567;
        else
            _1428 <= _69;
    end
    assign _1436 = 8'b11000000;
    assign _1437 = _616 == _1436;
    assign _1435 = _565 & _570;
    assign _1438 = _1435 & _1437;
    assign _1442 = _1438 ? _599 : _1441;
    assign _1433 = _609 == _1436;
    assign _1431 = _565 & _580;
    assign _1434 = _1431 & _1433;
    assign _1443 = _1434 ? _583 : _1442;
    assign _70 = _1443;
    always @(posedge _539) begin
        if (_537)
            _1441 <= _567;
        else
            _1441 <= _70;
    end
    assign _1449 = 8'b10111111;
    assign _1450 = _616 == _1449;
    assign _1448 = _565 & _570;
    assign _1451 = _1448 & _1450;
    assign _1455 = _1451 ? _599 : _1454;
    assign _1446 = _609 == _1449;
    assign _1444 = _565 & _580;
    assign _1447 = _1444 & _1446;
    assign _1456 = _1447 ? _583 : _1455;
    assign _71 = _1456;
    always @(posedge _539) begin
        if (_537)
            _1454 <= _567;
        else
            _1454 <= _71;
    end
    assign _1462 = 8'b10111110;
    assign _1463 = _616 == _1462;
    assign _1461 = _565 & _570;
    assign _1464 = _1461 & _1463;
    assign _1468 = _1464 ? _599 : _1467;
    assign _1459 = _609 == _1462;
    assign _1457 = _565 & _580;
    assign _1460 = _1457 & _1459;
    assign _1469 = _1460 ? _583 : _1468;
    assign _72 = _1469;
    always @(posedge _539) begin
        if (_537)
            _1467 <= _567;
        else
            _1467 <= _72;
    end
    assign _1475 = 8'b10111101;
    assign _1476 = _616 == _1475;
    assign _1474 = _565 & _570;
    assign _1477 = _1474 & _1476;
    assign _1481 = _1477 ? _599 : _1480;
    assign _1472 = _609 == _1475;
    assign _1470 = _565 & _580;
    assign _1473 = _1470 & _1472;
    assign _1482 = _1473 ? _583 : _1481;
    assign _73 = _1482;
    always @(posedge _539) begin
        if (_537)
            _1480 <= _567;
        else
            _1480 <= _73;
    end
    assign _1488 = 8'b10111100;
    assign _1489 = _616 == _1488;
    assign _1487 = _565 & _570;
    assign _1490 = _1487 & _1489;
    assign _1494 = _1490 ? _599 : _1493;
    assign _1485 = _609 == _1488;
    assign _1483 = _565 & _580;
    assign _1486 = _1483 & _1485;
    assign _1495 = _1486 ? _583 : _1494;
    assign _74 = _1495;
    always @(posedge _539) begin
        if (_537)
            _1493 <= _567;
        else
            _1493 <= _74;
    end
    assign _1501 = 8'b10111011;
    assign _1502 = _616 == _1501;
    assign _1500 = _565 & _570;
    assign _1503 = _1500 & _1502;
    assign _1507 = _1503 ? _599 : _1506;
    assign _1498 = _609 == _1501;
    assign _1496 = _565 & _580;
    assign _1499 = _1496 & _1498;
    assign _1508 = _1499 ? _583 : _1507;
    assign _75 = _1508;
    always @(posedge _539) begin
        if (_537)
            _1506 <= _567;
        else
            _1506 <= _75;
    end
    assign _1514 = 8'b10111010;
    assign _1515 = _616 == _1514;
    assign _1513 = _565 & _570;
    assign _1516 = _1513 & _1515;
    assign _1520 = _1516 ? _599 : _1519;
    assign _1511 = _609 == _1514;
    assign _1509 = _565 & _580;
    assign _1512 = _1509 & _1511;
    assign _1521 = _1512 ? _583 : _1520;
    assign _76 = _1521;
    always @(posedge _539) begin
        if (_537)
            _1519 <= _567;
        else
            _1519 <= _76;
    end
    assign _1527 = 8'b10111001;
    assign _1528 = _616 == _1527;
    assign _1526 = _565 & _570;
    assign _1529 = _1526 & _1528;
    assign _1533 = _1529 ? _599 : _1532;
    assign _1524 = _609 == _1527;
    assign _1522 = _565 & _580;
    assign _1525 = _1522 & _1524;
    assign _1534 = _1525 ? _583 : _1533;
    assign _77 = _1534;
    always @(posedge _539) begin
        if (_537)
            _1532 <= _567;
        else
            _1532 <= _77;
    end
    assign _1540 = 8'b10111000;
    assign _1541 = _616 == _1540;
    assign _1539 = _565 & _570;
    assign _1542 = _1539 & _1541;
    assign _1546 = _1542 ? _599 : _1545;
    assign _1537 = _609 == _1540;
    assign _1535 = _565 & _580;
    assign _1538 = _1535 & _1537;
    assign _1547 = _1538 ? _583 : _1546;
    assign _78 = _1547;
    always @(posedge _539) begin
        if (_537)
            _1545 <= _567;
        else
            _1545 <= _78;
    end
    assign _1553 = 8'b10110111;
    assign _1554 = _616 == _1553;
    assign _1552 = _565 & _570;
    assign _1555 = _1552 & _1554;
    assign _1559 = _1555 ? _599 : _1558;
    assign _1550 = _609 == _1553;
    assign _1548 = _565 & _580;
    assign _1551 = _1548 & _1550;
    assign _1560 = _1551 ? _583 : _1559;
    assign _79 = _1560;
    always @(posedge _539) begin
        if (_537)
            _1558 <= _567;
        else
            _1558 <= _79;
    end
    assign _1566 = 8'b10110110;
    assign _1567 = _616 == _1566;
    assign _1565 = _565 & _570;
    assign _1568 = _1565 & _1567;
    assign _1572 = _1568 ? _599 : _1571;
    assign _1563 = _609 == _1566;
    assign _1561 = _565 & _580;
    assign _1564 = _1561 & _1563;
    assign _1573 = _1564 ? _583 : _1572;
    assign _80 = _1573;
    always @(posedge _539) begin
        if (_537)
            _1571 <= _567;
        else
            _1571 <= _80;
    end
    assign _1579 = 8'b10110101;
    assign _1580 = _616 == _1579;
    assign _1578 = _565 & _570;
    assign _1581 = _1578 & _1580;
    assign _1585 = _1581 ? _599 : _1584;
    assign _1576 = _609 == _1579;
    assign _1574 = _565 & _580;
    assign _1577 = _1574 & _1576;
    assign _1586 = _1577 ? _583 : _1585;
    assign _81 = _1586;
    always @(posedge _539) begin
        if (_537)
            _1584 <= _567;
        else
            _1584 <= _81;
    end
    assign _1592 = 8'b10110100;
    assign _1593 = _616 == _1592;
    assign _1591 = _565 & _570;
    assign _1594 = _1591 & _1593;
    assign _1598 = _1594 ? _599 : _1597;
    assign _1589 = _609 == _1592;
    assign _1587 = _565 & _580;
    assign _1590 = _1587 & _1589;
    assign _1599 = _1590 ? _583 : _1598;
    assign _82 = _1599;
    always @(posedge _539) begin
        if (_537)
            _1597 <= _567;
        else
            _1597 <= _82;
    end
    assign _1605 = 8'b10110011;
    assign _1606 = _616 == _1605;
    assign _1604 = _565 & _570;
    assign _1607 = _1604 & _1606;
    assign _1611 = _1607 ? _599 : _1610;
    assign _1602 = _609 == _1605;
    assign _1600 = _565 & _580;
    assign _1603 = _1600 & _1602;
    assign _1612 = _1603 ? _583 : _1611;
    assign _83 = _1612;
    always @(posedge _539) begin
        if (_537)
            _1610 <= _567;
        else
            _1610 <= _83;
    end
    assign _1618 = 8'b10110010;
    assign _1619 = _616 == _1618;
    assign _1617 = _565 & _570;
    assign _1620 = _1617 & _1619;
    assign _1624 = _1620 ? _599 : _1623;
    assign _1615 = _609 == _1618;
    assign _1613 = _565 & _580;
    assign _1616 = _1613 & _1615;
    assign _1625 = _1616 ? _583 : _1624;
    assign _84 = _1625;
    always @(posedge _539) begin
        if (_537)
            _1623 <= _567;
        else
            _1623 <= _84;
    end
    assign _1631 = 8'b10110001;
    assign _1632 = _616 == _1631;
    assign _1630 = _565 & _570;
    assign _1633 = _1630 & _1632;
    assign _1637 = _1633 ? _599 : _1636;
    assign _1628 = _609 == _1631;
    assign _1626 = _565 & _580;
    assign _1629 = _1626 & _1628;
    assign _1638 = _1629 ? _583 : _1637;
    assign _85 = _1638;
    always @(posedge _539) begin
        if (_537)
            _1636 <= _567;
        else
            _1636 <= _85;
    end
    assign _1644 = 8'b10110000;
    assign _1645 = _616 == _1644;
    assign _1643 = _565 & _570;
    assign _1646 = _1643 & _1645;
    assign _1650 = _1646 ? _599 : _1649;
    assign _1641 = _609 == _1644;
    assign _1639 = _565 & _580;
    assign _1642 = _1639 & _1641;
    assign _1651 = _1642 ? _583 : _1650;
    assign _86 = _1651;
    always @(posedge _539) begin
        if (_537)
            _1649 <= _567;
        else
            _1649 <= _86;
    end
    assign _1657 = 8'b10101111;
    assign _1658 = _616 == _1657;
    assign _1656 = _565 & _570;
    assign _1659 = _1656 & _1658;
    assign _1663 = _1659 ? _599 : _1662;
    assign _1654 = _609 == _1657;
    assign _1652 = _565 & _580;
    assign _1655 = _1652 & _1654;
    assign _1664 = _1655 ? _583 : _1663;
    assign _87 = _1664;
    always @(posedge _539) begin
        if (_537)
            _1662 <= _567;
        else
            _1662 <= _87;
    end
    assign _1670 = 8'b10101110;
    assign _1671 = _616 == _1670;
    assign _1669 = _565 & _570;
    assign _1672 = _1669 & _1671;
    assign _1676 = _1672 ? _599 : _1675;
    assign _1667 = _609 == _1670;
    assign _1665 = _565 & _580;
    assign _1668 = _1665 & _1667;
    assign _1677 = _1668 ? _583 : _1676;
    assign _88 = _1677;
    always @(posedge _539) begin
        if (_537)
            _1675 <= _567;
        else
            _1675 <= _88;
    end
    assign _1683 = 8'b10101101;
    assign _1684 = _616 == _1683;
    assign _1682 = _565 & _570;
    assign _1685 = _1682 & _1684;
    assign _1689 = _1685 ? _599 : _1688;
    assign _1680 = _609 == _1683;
    assign _1678 = _565 & _580;
    assign _1681 = _1678 & _1680;
    assign _1690 = _1681 ? _583 : _1689;
    assign _89 = _1690;
    always @(posedge _539) begin
        if (_537)
            _1688 <= _567;
        else
            _1688 <= _89;
    end
    assign _1696 = 8'b10101100;
    assign _1697 = _616 == _1696;
    assign _1695 = _565 & _570;
    assign _1698 = _1695 & _1697;
    assign _1702 = _1698 ? _599 : _1701;
    assign _1693 = _609 == _1696;
    assign _1691 = _565 & _580;
    assign _1694 = _1691 & _1693;
    assign _1703 = _1694 ? _583 : _1702;
    assign _90 = _1703;
    always @(posedge _539) begin
        if (_537)
            _1701 <= _567;
        else
            _1701 <= _90;
    end
    assign _1709 = 8'b10101011;
    assign _1710 = _616 == _1709;
    assign _1708 = _565 & _570;
    assign _1711 = _1708 & _1710;
    assign _1715 = _1711 ? _599 : _1714;
    assign _1706 = _609 == _1709;
    assign _1704 = _565 & _580;
    assign _1707 = _1704 & _1706;
    assign _1716 = _1707 ? _583 : _1715;
    assign _91 = _1716;
    always @(posedge _539) begin
        if (_537)
            _1714 <= _567;
        else
            _1714 <= _91;
    end
    assign _1722 = 8'b10101010;
    assign _1723 = _616 == _1722;
    assign _1721 = _565 & _570;
    assign _1724 = _1721 & _1723;
    assign _1728 = _1724 ? _599 : _1727;
    assign _1719 = _609 == _1722;
    assign _1717 = _565 & _580;
    assign _1720 = _1717 & _1719;
    assign _1729 = _1720 ? _583 : _1728;
    assign _92 = _1729;
    always @(posedge _539) begin
        if (_537)
            _1727 <= _567;
        else
            _1727 <= _92;
    end
    assign _1735 = 8'b10101001;
    assign _1736 = _616 == _1735;
    assign _1734 = _565 & _570;
    assign _1737 = _1734 & _1736;
    assign _1741 = _1737 ? _599 : _1740;
    assign _1732 = _609 == _1735;
    assign _1730 = _565 & _580;
    assign _1733 = _1730 & _1732;
    assign _1742 = _1733 ? _583 : _1741;
    assign _93 = _1742;
    always @(posedge _539) begin
        if (_537)
            _1740 <= _567;
        else
            _1740 <= _93;
    end
    assign _1748 = 8'b10101000;
    assign _1749 = _616 == _1748;
    assign _1747 = _565 & _570;
    assign _1750 = _1747 & _1749;
    assign _1754 = _1750 ? _599 : _1753;
    assign _1745 = _609 == _1748;
    assign _1743 = _565 & _580;
    assign _1746 = _1743 & _1745;
    assign _1755 = _1746 ? _583 : _1754;
    assign _94 = _1755;
    always @(posedge _539) begin
        if (_537)
            _1753 <= _567;
        else
            _1753 <= _94;
    end
    assign _1761 = 8'b10100111;
    assign _1762 = _616 == _1761;
    assign _1760 = _565 & _570;
    assign _1763 = _1760 & _1762;
    assign _1767 = _1763 ? _599 : _1766;
    assign _1758 = _609 == _1761;
    assign _1756 = _565 & _580;
    assign _1759 = _1756 & _1758;
    assign _1768 = _1759 ? _583 : _1767;
    assign _95 = _1768;
    always @(posedge _539) begin
        if (_537)
            _1766 <= _567;
        else
            _1766 <= _95;
    end
    assign _1774 = 8'b10100110;
    assign _1775 = _616 == _1774;
    assign _1773 = _565 & _570;
    assign _1776 = _1773 & _1775;
    assign _1780 = _1776 ? _599 : _1779;
    assign _1771 = _609 == _1774;
    assign _1769 = _565 & _580;
    assign _1772 = _1769 & _1771;
    assign _1781 = _1772 ? _583 : _1780;
    assign _96 = _1781;
    always @(posedge _539) begin
        if (_537)
            _1779 <= _567;
        else
            _1779 <= _96;
    end
    assign _1787 = 8'b10100101;
    assign _1788 = _616 == _1787;
    assign _1786 = _565 & _570;
    assign _1789 = _1786 & _1788;
    assign _1793 = _1789 ? _599 : _1792;
    assign _1784 = _609 == _1787;
    assign _1782 = _565 & _580;
    assign _1785 = _1782 & _1784;
    assign _1794 = _1785 ? _583 : _1793;
    assign _97 = _1794;
    always @(posedge _539) begin
        if (_537)
            _1792 <= _567;
        else
            _1792 <= _97;
    end
    assign _1800 = 8'b10100100;
    assign _1801 = _616 == _1800;
    assign _1799 = _565 & _570;
    assign _1802 = _1799 & _1801;
    assign _1806 = _1802 ? _599 : _1805;
    assign _1797 = _609 == _1800;
    assign _1795 = _565 & _580;
    assign _1798 = _1795 & _1797;
    assign _1807 = _1798 ? _583 : _1806;
    assign _98 = _1807;
    always @(posedge _539) begin
        if (_537)
            _1805 <= _567;
        else
            _1805 <= _98;
    end
    assign _1813 = 8'b10100011;
    assign _1814 = _616 == _1813;
    assign _1812 = _565 & _570;
    assign _1815 = _1812 & _1814;
    assign _1819 = _1815 ? _599 : _1818;
    assign _1810 = _609 == _1813;
    assign _1808 = _565 & _580;
    assign _1811 = _1808 & _1810;
    assign _1820 = _1811 ? _583 : _1819;
    assign _99 = _1820;
    always @(posedge _539) begin
        if (_537)
            _1818 <= _567;
        else
            _1818 <= _99;
    end
    assign _1826 = 8'b10100010;
    assign _1827 = _616 == _1826;
    assign _1825 = _565 & _570;
    assign _1828 = _1825 & _1827;
    assign _1832 = _1828 ? _599 : _1831;
    assign _1823 = _609 == _1826;
    assign _1821 = _565 & _580;
    assign _1824 = _1821 & _1823;
    assign _1833 = _1824 ? _583 : _1832;
    assign _100 = _1833;
    always @(posedge _539) begin
        if (_537)
            _1831 <= _567;
        else
            _1831 <= _100;
    end
    assign _1839 = 8'b10100001;
    assign _1840 = _616 == _1839;
    assign _1838 = _565 & _570;
    assign _1841 = _1838 & _1840;
    assign _1845 = _1841 ? _599 : _1844;
    assign _1836 = _609 == _1839;
    assign _1834 = _565 & _580;
    assign _1837 = _1834 & _1836;
    assign _1846 = _1837 ? _583 : _1845;
    assign _101 = _1846;
    always @(posedge _539) begin
        if (_537)
            _1844 <= _567;
        else
            _1844 <= _101;
    end
    assign _1852 = 8'b10100000;
    assign _1853 = _616 == _1852;
    assign _1851 = _565 & _570;
    assign _1854 = _1851 & _1853;
    assign _1858 = _1854 ? _599 : _1857;
    assign _1849 = _609 == _1852;
    assign _1847 = _565 & _580;
    assign _1850 = _1847 & _1849;
    assign _1859 = _1850 ? _583 : _1858;
    assign _102 = _1859;
    always @(posedge _539) begin
        if (_537)
            _1857 <= _567;
        else
            _1857 <= _102;
    end
    assign _1865 = 8'b10011111;
    assign _1866 = _616 == _1865;
    assign _1864 = _565 & _570;
    assign _1867 = _1864 & _1866;
    assign _1871 = _1867 ? _599 : _1870;
    assign _1862 = _609 == _1865;
    assign _1860 = _565 & _580;
    assign _1863 = _1860 & _1862;
    assign _1872 = _1863 ? _583 : _1871;
    assign _103 = _1872;
    always @(posedge _539) begin
        if (_537)
            _1870 <= _567;
        else
            _1870 <= _103;
    end
    assign _1878 = 8'b10011110;
    assign _1879 = _616 == _1878;
    assign _1877 = _565 & _570;
    assign _1880 = _1877 & _1879;
    assign _1884 = _1880 ? _599 : _1883;
    assign _1875 = _609 == _1878;
    assign _1873 = _565 & _580;
    assign _1876 = _1873 & _1875;
    assign _1885 = _1876 ? _583 : _1884;
    assign _104 = _1885;
    always @(posedge _539) begin
        if (_537)
            _1883 <= _567;
        else
            _1883 <= _104;
    end
    assign _1891 = 8'b10011101;
    assign _1892 = _616 == _1891;
    assign _1890 = _565 & _570;
    assign _1893 = _1890 & _1892;
    assign _1897 = _1893 ? _599 : _1896;
    assign _1888 = _609 == _1891;
    assign _1886 = _565 & _580;
    assign _1889 = _1886 & _1888;
    assign _1898 = _1889 ? _583 : _1897;
    assign _105 = _1898;
    always @(posedge _539) begin
        if (_537)
            _1896 <= _567;
        else
            _1896 <= _105;
    end
    assign _1904 = 8'b10011100;
    assign _1905 = _616 == _1904;
    assign _1903 = _565 & _570;
    assign _1906 = _1903 & _1905;
    assign _1910 = _1906 ? _599 : _1909;
    assign _1901 = _609 == _1904;
    assign _1899 = _565 & _580;
    assign _1902 = _1899 & _1901;
    assign _1911 = _1902 ? _583 : _1910;
    assign _106 = _1911;
    always @(posedge _539) begin
        if (_537)
            _1909 <= _567;
        else
            _1909 <= _106;
    end
    assign _1917 = 8'b10011011;
    assign _1918 = _616 == _1917;
    assign _1916 = _565 & _570;
    assign _1919 = _1916 & _1918;
    assign _1923 = _1919 ? _599 : _1922;
    assign _1914 = _609 == _1917;
    assign _1912 = _565 & _580;
    assign _1915 = _1912 & _1914;
    assign _1924 = _1915 ? _583 : _1923;
    assign _107 = _1924;
    always @(posedge _539) begin
        if (_537)
            _1922 <= _567;
        else
            _1922 <= _107;
    end
    assign _1930 = 8'b10011010;
    assign _1931 = _616 == _1930;
    assign _1929 = _565 & _570;
    assign _1932 = _1929 & _1931;
    assign _1936 = _1932 ? _599 : _1935;
    assign _1927 = _609 == _1930;
    assign _1925 = _565 & _580;
    assign _1928 = _1925 & _1927;
    assign _1937 = _1928 ? _583 : _1936;
    assign _108 = _1937;
    always @(posedge _539) begin
        if (_537)
            _1935 <= _567;
        else
            _1935 <= _108;
    end
    assign _1943 = 8'b10011001;
    assign _1944 = _616 == _1943;
    assign _1942 = _565 & _570;
    assign _1945 = _1942 & _1944;
    assign _1949 = _1945 ? _599 : _1948;
    assign _1940 = _609 == _1943;
    assign _1938 = _565 & _580;
    assign _1941 = _1938 & _1940;
    assign _1950 = _1941 ? _583 : _1949;
    assign _109 = _1950;
    always @(posedge _539) begin
        if (_537)
            _1948 <= _567;
        else
            _1948 <= _109;
    end
    assign _1956 = 8'b10011000;
    assign _1957 = _616 == _1956;
    assign _1955 = _565 & _570;
    assign _1958 = _1955 & _1957;
    assign _1962 = _1958 ? _599 : _1961;
    assign _1953 = _609 == _1956;
    assign _1951 = _565 & _580;
    assign _1954 = _1951 & _1953;
    assign _1963 = _1954 ? _583 : _1962;
    assign _110 = _1963;
    always @(posedge _539) begin
        if (_537)
            _1961 <= _567;
        else
            _1961 <= _110;
    end
    assign _1969 = 8'b10010111;
    assign _1970 = _616 == _1969;
    assign _1968 = _565 & _570;
    assign _1971 = _1968 & _1970;
    assign _1975 = _1971 ? _599 : _1974;
    assign _1966 = _609 == _1969;
    assign _1964 = _565 & _580;
    assign _1967 = _1964 & _1966;
    assign _1976 = _1967 ? _583 : _1975;
    assign _111 = _1976;
    always @(posedge _539) begin
        if (_537)
            _1974 <= _567;
        else
            _1974 <= _111;
    end
    assign _1982 = 8'b10010110;
    assign _1983 = _616 == _1982;
    assign _1981 = _565 & _570;
    assign _1984 = _1981 & _1983;
    assign _1988 = _1984 ? _599 : _1987;
    assign _1979 = _609 == _1982;
    assign _1977 = _565 & _580;
    assign _1980 = _1977 & _1979;
    assign _1989 = _1980 ? _583 : _1988;
    assign _112 = _1989;
    always @(posedge _539) begin
        if (_537)
            _1987 <= _567;
        else
            _1987 <= _112;
    end
    assign _1995 = 8'b10010101;
    assign _1996 = _616 == _1995;
    assign _1994 = _565 & _570;
    assign _1997 = _1994 & _1996;
    assign _2001 = _1997 ? _599 : _2000;
    assign _1992 = _609 == _1995;
    assign _1990 = _565 & _580;
    assign _1993 = _1990 & _1992;
    assign _2002 = _1993 ? _583 : _2001;
    assign _113 = _2002;
    always @(posedge _539) begin
        if (_537)
            _2000 <= _567;
        else
            _2000 <= _113;
    end
    assign _2008 = 8'b10010100;
    assign _2009 = _616 == _2008;
    assign _2007 = _565 & _570;
    assign _2010 = _2007 & _2009;
    assign _2014 = _2010 ? _599 : _2013;
    assign _2005 = _609 == _2008;
    assign _2003 = _565 & _580;
    assign _2006 = _2003 & _2005;
    assign _2015 = _2006 ? _583 : _2014;
    assign _114 = _2015;
    always @(posedge _539) begin
        if (_537)
            _2013 <= _567;
        else
            _2013 <= _114;
    end
    assign _2021 = 8'b10010011;
    assign _2022 = _616 == _2021;
    assign _2020 = _565 & _570;
    assign _2023 = _2020 & _2022;
    assign _2027 = _2023 ? _599 : _2026;
    assign _2018 = _609 == _2021;
    assign _2016 = _565 & _580;
    assign _2019 = _2016 & _2018;
    assign _2028 = _2019 ? _583 : _2027;
    assign _115 = _2028;
    always @(posedge _539) begin
        if (_537)
            _2026 <= _567;
        else
            _2026 <= _115;
    end
    assign _2034 = 8'b10010010;
    assign _2035 = _616 == _2034;
    assign _2033 = _565 & _570;
    assign _2036 = _2033 & _2035;
    assign _2040 = _2036 ? _599 : _2039;
    assign _2031 = _609 == _2034;
    assign _2029 = _565 & _580;
    assign _2032 = _2029 & _2031;
    assign _2041 = _2032 ? _583 : _2040;
    assign _116 = _2041;
    always @(posedge _539) begin
        if (_537)
            _2039 <= _567;
        else
            _2039 <= _116;
    end
    assign _2047 = 8'b10010001;
    assign _2048 = _616 == _2047;
    assign _2046 = _565 & _570;
    assign _2049 = _2046 & _2048;
    assign _2053 = _2049 ? _599 : _2052;
    assign _2044 = _609 == _2047;
    assign _2042 = _565 & _580;
    assign _2045 = _2042 & _2044;
    assign _2054 = _2045 ? _583 : _2053;
    assign _117 = _2054;
    always @(posedge _539) begin
        if (_537)
            _2052 <= _567;
        else
            _2052 <= _117;
    end
    assign _2060 = 8'b10010000;
    assign _2061 = _616 == _2060;
    assign _2059 = _565 & _570;
    assign _2062 = _2059 & _2061;
    assign _2066 = _2062 ? _599 : _2065;
    assign _2057 = _609 == _2060;
    assign _2055 = _565 & _580;
    assign _2058 = _2055 & _2057;
    assign _2067 = _2058 ? _583 : _2066;
    assign _118 = _2067;
    always @(posedge _539) begin
        if (_537)
            _2065 <= _567;
        else
            _2065 <= _118;
    end
    assign _2073 = 8'b10001111;
    assign _2074 = _616 == _2073;
    assign _2072 = _565 & _570;
    assign _2075 = _2072 & _2074;
    assign _2079 = _2075 ? _599 : _2078;
    assign _2070 = _609 == _2073;
    assign _2068 = _565 & _580;
    assign _2071 = _2068 & _2070;
    assign _2080 = _2071 ? _583 : _2079;
    assign _119 = _2080;
    always @(posedge _539) begin
        if (_537)
            _2078 <= _567;
        else
            _2078 <= _119;
    end
    assign _2086 = 8'b10001110;
    assign _2087 = _616 == _2086;
    assign _2085 = _565 & _570;
    assign _2088 = _2085 & _2087;
    assign _2092 = _2088 ? _599 : _2091;
    assign _2083 = _609 == _2086;
    assign _2081 = _565 & _580;
    assign _2084 = _2081 & _2083;
    assign _2093 = _2084 ? _583 : _2092;
    assign _120 = _2093;
    always @(posedge _539) begin
        if (_537)
            _2091 <= _567;
        else
            _2091 <= _120;
    end
    assign _2099 = 8'b10001101;
    assign _2100 = _616 == _2099;
    assign _2098 = _565 & _570;
    assign _2101 = _2098 & _2100;
    assign _2105 = _2101 ? _599 : _2104;
    assign _2096 = _609 == _2099;
    assign _2094 = _565 & _580;
    assign _2097 = _2094 & _2096;
    assign _2106 = _2097 ? _583 : _2105;
    assign _121 = _2106;
    always @(posedge _539) begin
        if (_537)
            _2104 <= _567;
        else
            _2104 <= _121;
    end
    assign _2112 = 8'b10001100;
    assign _2113 = _616 == _2112;
    assign _2111 = _565 & _570;
    assign _2114 = _2111 & _2113;
    assign _2118 = _2114 ? _599 : _2117;
    assign _2109 = _609 == _2112;
    assign _2107 = _565 & _580;
    assign _2110 = _2107 & _2109;
    assign _2119 = _2110 ? _583 : _2118;
    assign _122 = _2119;
    always @(posedge _539) begin
        if (_537)
            _2117 <= _567;
        else
            _2117 <= _122;
    end
    assign _2125 = 8'b10001011;
    assign _2126 = _616 == _2125;
    assign _2124 = _565 & _570;
    assign _2127 = _2124 & _2126;
    assign _2131 = _2127 ? _599 : _2130;
    assign _2122 = _609 == _2125;
    assign _2120 = _565 & _580;
    assign _2123 = _2120 & _2122;
    assign _2132 = _2123 ? _583 : _2131;
    assign _123 = _2132;
    always @(posedge _539) begin
        if (_537)
            _2130 <= _567;
        else
            _2130 <= _123;
    end
    assign _2138 = 8'b10001010;
    assign _2139 = _616 == _2138;
    assign _2137 = _565 & _570;
    assign _2140 = _2137 & _2139;
    assign _2144 = _2140 ? _599 : _2143;
    assign _2135 = _609 == _2138;
    assign _2133 = _565 & _580;
    assign _2136 = _2133 & _2135;
    assign _2145 = _2136 ? _583 : _2144;
    assign _124 = _2145;
    always @(posedge _539) begin
        if (_537)
            _2143 <= _567;
        else
            _2143 <= _124;
    end
    assign _2151 = 8'b10001001;
    assign _2152 = _616 == _2151;
    assign _2150 = _565 & _570;
    assign _2153 = _2150 & _2152;
    assign _2157 = _2153 ? _599 : _2156;
    assign _2148 = _609 == _2151;
    assign _2146 = _565 & _580;
    assign _2149 = _2146 & _2148;
    assign _2158 = _2149 ? _583 : _2157;
    assign _125 = _2158;
    always @(posedge _539) begin
        if (_537)
            _2156 <= _567;
        else
            _2156 <= _125;
    end
    assign _2164 = 8'b10001000;
    assign _2165 = _616 == _2164;
    assign _2163 = _565 & _570;
    assign _2166 = _2163 & _2165;
    assign _2170 = _2166 ? _599 : _2169;
    assign _2161 = _609 == _2164;
    assign _2159 = _565 & _580;
    assign _2162 = _2159 & _2161;
    assign _2171 = _2162 ? _583 : _2170;
    assign _126 = _2171;
    always @(posedge _539) begin
        if (_537)
            _2169 <= _567;
        else
            _2169 <= _126;
    end
    assign _2177 = 8'b10000111;
    assign _2178 = _616 == _2177;
    assign _2176 = _565 & _570;
    assign _2179 = _2176 & _2178;
    assign _2183 = _2179 ? _599 : _2182;
    assign _2174 = _609 == _2177;
    assign _2172 = _565 & _580;
    assign _2175 = _2172 & _2174;
    assign _2184 = _2175 ? _583 : _2183;
    assign _127 = _2184;
    always @(posedge _539) begin
        if (_537)
            _2182 <= _567;
        else
            _2182 <= _127;
    end
    assign _2190 = 8'b10000110;
    assign _2191 = _616 == _2190;
    assign _2189 = _565 & _570;
    assign _2192 = _2189 & _2191;
    assign _2196 = _2192 ? _599 : _2195;
    assign _2187 = _609 == _2190;
    assign _2185 = _565 & _580;
    assign _2188 = _2185 & _2187;
    assign _2197 = _2188 ? _583 : _2196;
    assign _128 = _2197;
    always @(posedge _539) begin
        if (_537)
            _2195 <= _567;
        else
            _2195 <= _128;
    end
    assign _2203 = 8'b10000101;
    assign _2204 = _616 == _2203;
    assign _2202 = _565 & _570;
    assign _2205 = _2202 & _2204;
    assign _2209 = _2205 ? _599 : _2208;
    assign _2200 = _609 == _2203;
    assign _2198 = _565 & _580;
    assign _2201 = _2198 & _2200;
    assign _2210 = _2201 ? _583 : _2209;
    assign _129 = _2210;
    always @(posedge _539) begin
        if (_537)
            _2208 <= _567;
        else
            _2208 <= _129;
    end
    assign _2216 = 8'b10000100;
    assign _2217 = _616 == _2216;
    assign _2215 = _565 & _570;
    assign _2218 = _2215 & _2217;
    assign _2222 = _2218 ? _599 : _2221;
    assign _2213 = _609 == _2216;
    assign _2211 = _565 & _580;
    assign _2214 = _2211 & _2213;
    assign _2223 = _2214 ? _583 : _2222;
    assign _130 = _2223;
    always @(posedge _539) begin
        if (_537)
            _2221 <= _567;
        else
            _2221 <= _130;
    end
    assign _2229 = 8'b10000011;
    assign _2230 = _616 == _2229;
    assign _2228 = _565 & _570;
    assign _2231 = _2228 & _2230;
    assign _2235 = _2231 ? _599 : _2234;
    assign _2226 = _609 == _2229;
    assign _2224 = _565 & _580;
    assign _2227 = _2224 & _2226;
    assign _2236 = _2227 ? _583 : _2235;
    assign _131 = _2236;
    always @(posedge _539) begin
        if (_537)
            _2234 <= _567;
        else
            _2234 <= _131;
    end
    assign _2242 = 8'b10000010;
    assign _2243 = _616 == _2242;
    assign _2241 = _565 & _570;
    assign _2244 = _2241 & _2243;
    assign _2248 = _2244 ? _599 : _2247;
    assign _2239 = _609 == _2242;
    assign _2237 = _565 & _580;
    assign _2240 = _2237 & _2239;
    assign _2249 = _2240 ? _583 : _2248;
    assign _132 = _2249;
    always @(posedge _539) begin
        if (_537)
            _2247 <= _567;
        else
            _2247 <= _132;
    end
    assign _2255 = 8'b10000001;
    assign _2256 = _616 == _2255;
    assign _2254 = _565 & _570;
    assign _2257 = _2254 & _2256;
    assign _2261 = _2257 ? _599 : _2260;
    assign _2252 = _609 == _2255;
    assign _2250 = _565 & _580;
    assign _2253 = _2250 & _2252;
    assign _2262 = _2253 ? _583 : _2261;
    assign _133 = _2262;
    always @(posedge _539) begin
        if (_537)
            _2260 <= _567;
        else
            _2260 <= _133;
    end
    assign _2268 = 8'b10000000;
    assign _2269 = _616 == _2268;
    assign _2267 = _565 & _570;
    assign _2270 = _2267 & _2269;
    assign _2274 = _2270 ? _599 : _2273;
    assign _2265 = _609 == _2268;
    assign _2263 = _565 & _580;
    assign _2266 = _2263 & _2265;
    assign _2275 = _2266 ? _583 : _2274;
    assign _134 = _2275;
    always @(posedge _539) begin
        if (_537)
            _2273 <= _567;
        else
            _2273 <= _134;
    end
    assign _2281 = 8'b01111111;
    assign _2282 = _616 == _2281;
    assign _2280 = _565 & _570;
    assign _2283 = _2280 & _2282;
    assign _2287 = _2283 ? _599 : _2286;
    assign _2278 = _609 == _2281;
    assign _2276 = _565 & _580;
    assign _2279 = _2276 & _2278;
    assign _2288 = _2279 ? _583 : _2287;
    assign _135 = _2288;
    always @(posedge _539) begin
        if (_537)
            _2286 <= _567;
        else
            _2286 <= _135;
    end
    assign _2294 = 8'b01111110;
    assign _2295 = _616 == _2294;
    assign _2293 = _565 & _570;
    assign _2296 = _2293 & _2295;
    assign _2300 = _2296 ? _599 : _2299;
    assign _2291 = _609 == _2294;
    assign _2289 = _565 & _580;
    assign _2292 = _2289 & _2291;
    assign _2301 = _2292 ? _583 : _2300;
    assign _136 = _2301;
    always @(posedge _539) begin
        if (_537)
            _2299 <= _567;
        else
            _2299 <= _136;
    end
    assign _2307 = 8'b01111101;
    assign _2308 = _616 == _2307;
    assign _2306 = _565 & _570;
    assign _2309 = _2306 & _2308;
    assign _2313 = _2309 ? _599 : _2312;
    assign _2304 = _609 == _2307;
    assign _2302 = _565 & _580;
    assign _2305 = _2302 & _2304;
    assign _2314 = _2305 ? _583 : _2313;
    assign _137 = _2314;
    always @(posedge _539) begin
        if (_537)
            _2312 <= _567;
        else
            _2312 <= _137;
    end
    assign _2320 = 8'b01111100;
    assign _2321 = _616 == _2320;
    assign _2319 = _565 & _570;
    assign _2322 = _2319 & _2321;
    assign _2326 = _2322 ? _599 : _2325;
    assign _2317 = _609 == _2320;
    assign _2315 = _565 & _580;
    assign _2318 = _2315 & _2317;
    assign _2327 = _2318 ? _583 : _2326;
    assign _138 = _2327;
    always @(posedge _539) begin
        if (_537)
            _2325 <= _567;
        else
            _2325 <= _138;
    end
    assign _2333 = 8'b01111011;
    assign _2334 = _616 == _2333;
    assign _2332 = _565 & _570;
    assign _2335 = _2332 & _2334;
    assign _2339 = _2335 ? _599 : _2338;
    assign _2330 = _609 == _2333;
    assign _2328 = _565 & _580;
    assign _2331 = _2328 & _2330;
    assign _2340 = _2331 ? _583 : _2339;
    assign _139 = _2340;
    always @(posedge _539) begin
        if (_537)
            _2338 <= _567;
        else
            _2338 <= _139;
    end
    assign _2346 = 8'b01111010;
    assign _2347 = _616 == _2346;
    assign _2345 = _565 & _570;
    assign _2348 = _2345 & _2347;
    assign _2352 = _2348 ? _599 : _2351;
    assign _2343 = _609 == _2346;
    assign _2341 = _565 & _580;
    assign _2344 = _2341 & _2343;
    assign _2353 = _2344 ? _583 : _2352;
    assign _140 = _2353;
    always @(posedge _539) begin
        if (_537)
            _2351 <= _567;
        else
            _2351 <= _140;
    end
    assign _2359 = 8'b01111001;
    assign _2360 = _616 == _2359;
    assign _2358 = _565 & _570;
    assign _2361 = _2358 & _2360;
    assign _2365 = _2361 ? _599 : _2364;
    assign _2356 = _609 == _2359;
    assign _2354 = _565 & _580;
    assign _2357 = _2354 & _2356;
    assign _2366 = _2357 ? _583 : _2365;
    assign _141 = _2366;
    always @(posedge _539) begin
        if (_537)
            _2364 <= _567;
        else
            _2364 <= _141;
    end
    assign _2372 = 8'b01111000;
    assign _2373 = _616 == _2372;
    assign _2371 = _565 & _570;
    assign _2374 = _2371 & _2373;
    assign _2378 = _2374 ? _599 : _2377;
    assign _2369 = _609 == _2372;
    assign _2367 = _565 & _580;
    assign _2370 = _2367 & _2369;
    assign _2379 = _2370 ? _583 : _2378;
    assign _142 = _2379;
    always @(posedge _539) begin
        if (_537)
            _2377 <= _567;
        else
            _2377 <= _142;
    end
    assign _2385 = 8'b01110111;
    assign _2386 = _616 == _2385;
    assign _2384 = _565 & _570;
    assign _2387 = _2384 & _2386;
    assign _2391 = _2387 ? _599 : _2390;
    assign _2382 = _609 == _2385;
    assign _2380 = _565 & _580;
    assign _2383 = _2380 & _2382;
    assign _2392 = _2383 ? _583 : _2391;
    assign _143 = _2392;
    always @(posedge _539) begin
        if (_537)
            _2390 <= _567;
        else
            _2390 <= _143;
    end
    assign _2398 = 8'b01110110;
    assign _2399 = _616 == _2398;
    assign _2397 = _565 & _570;
    assign _2400 = _2397 & _2399;
    assign _2404 = _2400 ? _599 : _2403;
    assign _2395 = _609 == _2398;
    assign _2393 = _565 & _580;
    assign _2396 = _2393 & _2395;
    assign _2405 = _2396 ? _583 : _2404;
    assign _144 = _2405;
    always @(posedge _539) begin
        if (_537)
            _2403 <= _567;
        else
            _2403 <= _144;
    end
    assign _2411 = 8'b01110101;
    assign _2412 = _616 == _2411;
    assign _2410 = _565 & _570;
    assign _2413 = _2410 & _2412;
    assign _2417 = _2413 ? _599 : _2416;
    assign _2408 = _609 == _2411;
    assign _2406 = _565 & _580;
    assign _2409 = _2406 & _2408;
    assign _2418 = _2409 ? _583 : _2417;
    assign _145 = _2418;
    always @(posedge _539) begin
        if (_537)
            _2416 <= _567;
        else
            _2416 <= _145;
    end
    assign _2424 = 8'b01110100;
    assign _2425 = _616 == _2424;
    assign _2423 = _565 & _570;
    assign _2426 = _2423 & _2425;
    assign _2430 = _2426 ? _599 : _2429;
    assign _2421 = _609 == _2424;
    assign _2419 = _565 & _580;
    assign _2422 = _2419 & _2421;
    assign _2431 = _2422 ? _583 : _2430;
    assign _146 = _2431;
    always @(posedge _539) begin
        if (_537)
            _2429 <= _567;
        else
            _2429 <= _146;
    end
    assign _2437 = 8'b01110011;
    assign _2438 = _616 == _2437;
    assign _2436 = _565 & _570;
    assign _2439 = _2436 & _2438;
    assign _2443 = _2439 ? _599 : _2442;
    assign _2434 = _609 == _2437;
    assign _2432 = _565 & _580;
    assign _2435 = _2432 & _2434;
    assign _2444 = _2435 ? _583 : _2443;
    assign _147 = _2444;
    always @(posedge _539) begin
        if (_537)
            _2442 <= _567;
        else
            _2442 <= _147;
    end
    assign _2450 = 8'b01110010;
    assign _2451 = _616 == _2450;
    assign _2449 = _565 & _570;
    assign _2452 = _2449 & _2451;
    assign _2456 = _2452 ? _599 : _2455;
    assign _2447 = _609 == _2450;
    assign _2445 = _565 & _580;
    assign _2448 = _2445 & _2447;
    assign _2457 = _2448 ? _583 : _2456;
    assign _148 = _2457;
    always @(posedge _539) begin
        if (_537)
            _2455 <= _567;
        else
            _2455 <= _148;
    end
    assign _2463 = 8'b01110001;
    assign _2464 = _616 == _2463;
    assign _2462 = _565 & _570;
    assign _2465 = _2462 & _2464;
    assign _2469 = _2465 ? _599 : _2468;
    assign _2460 = _609 == _2463;
    assign _2458 = _565 & _580;
    assign _2461 = _2458 & _2460;
    assign _2470 = _2461 ? _583 : _2469;
    assign _149 = _2470;
    always @(posedge _539) begin
        if (_537)
            _2468 <= _567;
        else
            _2468 <= _149;
    end
    assign _2476 = 8'b01110000;
    assign _2477 = _616 == _2476;
    assign _2475 = _565 & _570;
    assign _2478 = _2475 & _2477;
    assign _2482 = _2478 ? _599 : _2481;
    assign _2473 = _609 == _2476;
    assign _2471 = _565 & _580;
    assign _2474 = _2471 & _2473;
    assign _2483 = _2474 ? _583 : _2482;
    assign _150 = _2483;
    always @(posedge _539) begin
        if (_537)
            _2481 <= _567;
        else
            _2481 <= _150;
    end
    assign _2489 = 8'b01101111;
    assign _2490 = _616 == _2489;
    assign _2488 = _565 & _570;
    assign _2491 = _2488 & _2490;
    assign _2495 = _2491 ? _599 : _2494;
    assign _2486 = _609 == _2489;
    assign _2484 = _565 & _580;
    assign _2487 = _2484 & _2486;
    assign _2496 = _2487 ? _583 : _2495;
    assign _151 = _2496;
    always @(posedge _539) begin
        if (_537)
            _2494 <= _567;
        else
            _2494 <= _151;
    end
    assign _2502 = 8'b01101110;
    assign _2503 = _616 == _2502;
    assign _2501 = _565 & _570;
    assign _2504 = _2501 & _2503;
    assign _2508 = _2504 ? _599 : _2507;
    assign _2499 = _609 == _2502;
    assign _2497 = _565 & _580;
    assign _2500 = _2497 & _2499;
    assign _2509 = _2500 ? _583 : _2508;
    assign _152 = _2509;
    always @(posedge _539) begin
        if (_537)
            _2507 <= _567;
        else
            _2507 <= _152;
    end
    assign _2515 = 8'b01101101;
    assign _2516 = _616 == _2515;
    assign _2514 = _565 & _570;
    assign _2517 = _2514 & _2516;
    assign _2521 = _2517 ? _599 : _2520;
    assign _2512 = _609 == _2515;
    assign _2510 = _565 & _580;
    assign _2513 = _2510 & _2512;
    assign _2522 = _2513 ? _583 : _2521;
    assign _153 = _2522;
    always @(posedge _539) begin
        if (_537)
            _2520 <= _567;
        else
            _2520 <= _153;
    end
    assign _2528 = 8'b01101100;
    assign _2529 = _616 == _2528;
    assign _2527 = _565 & _570;
    assign _2530 = _2527 & _2529;
    assign _2534 = _2530 ? _599 : _2533;
    assign _2525 = _609 == _2528;
    assign _2523 = _565 & _580;
    assign _2526 = _2523 & _2525;
    assign _2535 = _2526 ? _583 : _2534;
    assign _154 = _2535;
    always @(posedge _539) begin
        if (_537)
            _2533 <= _567;
        else
            _2533 <= _154;
    end
    assign _2541 = 8'b01101011;
    assign _2542 = _616 == _2541;
    assign _2540 = _565 & _570;
    assign _2543 = _2540 & _2542;
    assign _2547 = _2543 ? _599 : _2546;
    assign _2538 = _609 == _2541;
    assign _2536 = _565 & _580;
    assign _2539 = _2536 & _2538;
    assign _2548 = _2539 ? _583 : _2547;
    assign _155 = _2548;
    always @(posedge _539) begin
        if (_537)
            _2546 <= _567;
        else
            _2546 <= _155;
    end
    assign _2554 = 8'b01101010;
    assign _2555 = _616 == _2554;
    assign _2553 = _565 & _570;
    assign _2556 = _2553 & _2555;
    assign _2560 = _2556 ? _599 : _2559;
    assign _2551 = _609 == _2554;
    assign _2549 = _565 & _580;
    assign _2552 = _2549 & _2551;
    assign _2561 = _2552 ? _583 : _2560;
    assign _156 = _2561;
    always @(posedge _539) begin
        if (_537)
            _2559 <= _567;
        else
            _2559 <= _156;
    end
    assign _2567 = 8'b01101001;
    assign _2568 = _616 == _2567;
    assign _2566 = _565 & _570;
    assign _2569 = _2566 & _2568;
    assign _2573 = _2569 ? _599 : _2572;
    assign _2564 = _609 == _2567;
    assign _2562 = _565 & _580;
    assign _2565 = _2562 & _2564;
    assign _2574 = _2565 ? _583 : _2573;
    assign _157 = _2574;
    always @(posedge _539) begin
        if (_537)
            _2572 <= _567;
        else
            _2572 <= _157;
    end
    assign _2580 = 8'b01101000;
    assign _2581 = _616 == _2580;
    assign _2579 = _565 & _570;
    assign _2582 = _2579 & _2581;
    assign _2586 = _2582 ? _599 : _2585;
    assign _2577 = _609 == _2580;
    assign _2575 = _565 & _580;
    assign _2578 = _2575 & _2577;
    assign _2587 = _2578 ? _583 : _2586;
    assign _158 = _2587;
    always @(posedge _539) begin
        if (_537)
            _2585 <= _567;
        else
            _2585 <= _158;
    end
    assign _2593 = 8'b01100111;
    assign _2594 = _616 == _2593;
    assign _2592 = _565 & _570;
    assign _2595 = _2592 & _2594;
    assign _2599 = _2595 ? _599 : _2598;
    assign _2590 = _609 == _2593;
    assign _2588 = _565 & _580;
    assign _2591 = _2588 & _2590;
    assign _2600 = _2591 ? _583 : _2599;
    assign _159 = _2600;
    always @(posedge _539) begin
        if (_537)
            _2598 <= _567;
        else
            _2598 <= _159;
    end
    assign _2606 = 8'b01100110;
    assign _2607 = _616 == _2606;
    assign _2605 = _565 & _570;
    assign _2608 = _2605 & _2607;
    assign _2612 = _2608 ? _599 : _2611;
    assign _2603 = _609 == _2606;
    assign _2601 = _565 & _580;
    assign _2604 = _2601 & _2603;
    assign _2613 = _2604 ? _583 : _2612;
    assign _160 = _2613;
    always @(posedge _539) begin
        if (_537)
            _2611 <= _567;
        else
            _2611 <= _160;
    end
    assign _2619 = 8'b01100101;
    assign _2620 = _616 == _2619;
    assign _2618 = _565 & _570;
    assign _2621 = _2618 & _2620;
    assign _2625 = _2621 ? _599 : _2624;
    assign _2616 = _609 == _2619;
    assign _2614 = _565 & _580;
    assign _2617 = _2614 & _2616;
    assign _2626 = _2617 ? _583 : _2625;
    assign _161 = _2626;
    always @(posedge _539) begin
        if (_537)
            _2624 <= _567;
        else
            _2624 <= _161;
    end
    assign _2632 = 8'b01100100;
    assign _2633 = _616 == _2632;
    assign _2631 = _565 & _570;
    assign _2634 = _2631 & _2633;
    assign _2638 = _2634 ? _599 : _2637;
    assign _2629 = _609 == _2632;
    assign _2627 = _565 & _580;
    assign _2630 = _2627 & _2629;
    assign _2639 = _2630 ? _583 : _2638;
    assign _162 = _2639;
    always @(posedge _539) begin
        if (_537)
            _2637 <= _567;
        else
            _2637 <= _162;
    end
    assign _2645 = 8'b01100011;
    assign _2646 = _616 == _2645;
    assign _2644 = _565 & _570;
    assign _2647 = _2644 & _2646;
    assign _2651 = _2647 ? _599 : _2650;
    assign _2642 = _609 == _2645;
    assign _2640 = _565 & _580;
    assign _2643 = _2640 & _2642;
    assign _2652 = _2643 ? _583 : _2651;
    assign _163 = _2652;
    always @(posedge _539) begin
        if (_537)
            _2650 <= _567;
        else
            _2650 <= _163;
    end
    assign _2658 = 8'b01100010;
    assign _2659 = _616 == _2658;
    assign _2657 = _565 & _570;
    assign _2660 = _2657 & _2659;
    assign _2664 = _2660 ? _599 : _2663;
    assign _2655 = _609 == _2658;
    assign _2653 = _565 & _580;
    assign _2656 = _2653 & _2655;
    assign _2665 = _2656 ? _583 : _2664;
    assign _164 = _2665;
    always @(posedge _539) begin
        if (_537)
            _2663 <= _567;
        else
            _2663 <= _164;
    end
    assign _2671 = 8'b01100001;
    assign _2672 = _616 == _2671;
    assign _2670 = _565 & _570;
    assign _2673 = _2670 & _2672;
    assign _2677 = _2673 ? _599 : _2676;
    assign _2668 = _609 == _2671;
    assign _2666 = _565 & _580;
    assign _2669 = _2666 & _2668;
    assign _2678 = _2669 ? _583 : _2677;
    assign _165 = _2678;
    always @(posedge _539) begin
        if (_537)
            _2676 <= _567;
        else
            _2676 <= _165;
    end
    assign _2684 = 8'b01100000;
    assign _2685 = _616 == _2684;
    assign _2683 = _565 & _570;
    assign _2686 = _2683 & _2685;
    assign _2690 = _2686 ? _599 : _2689;
    assign _2681 = _609 == _2684;
    assign _2679 = _565 & _580;
    assign _2682 = _2679 & _2681;
    assign _2691 = _2682 ? _583 : _2690;
    assign _166 = _2691;
    always @(posedge _539) begin
        if (_537)
            _2689 <= _567;
        else
            _2689 <= _166;
    end
    assign _2697 = 8'b01011111;
    assign _2698 = _616 == _2697;
    assign _2696 = _565 & _570;
    assign _2699 = _2696 & _2698;
    assign _2703 = _2699 ? _599 : _2702;
    assign _2694 = _609 == _2697;
    assign _2692 = _565 & _580;
    assign _2695 = _2692 & _2694;
    assign _2704 = _2695 ? _583 : _2703;
    assign _167 = _2704;
    always @(posedge _539) begin
        if (_537)
            _2702 <= _567;
        else
            _2702 <= _167;
    end
    assign _2710 = 8'b01011110;
    assign _2711 = _616 == _2710;
    assign _2709 = _565 & _570;
    assign _2712 = _2709 & _2711;
    assign _2716 = _2712 ? _599 : _2715;
    assign _2707 = _609 == _2710;
    assign _2705 = _565 & _580;
    assign _2708 = _2705 & _2707;
    assign _2717 = _2708 ? _583 : _2716;
    assign _168 = _2717;
    always @(posedge _539) begin
        if (_537)
            _2715 <= _567;
        else
            _2715 <= _168;
    end
    assign _2723 = 8'b01011101;
    assign _2724 = _616 == _2723;
    assign _2722 = _565 & _570;
    assign _2725 = _2722 & _2724;
    assign _2729 = _2725 ? _599 : _2728;
    assign _2720 = _609 == _2723;
    assign _2718 = _565 & _580;
    assign _2721 = _2718 & _2720;
    assign _2730 = _2721 ? _583 : _2729;
    assign _169 = _2730;
    always @(posedge _539) begin
        if (_537)
            _2728 <= _567;
        else
            _2728 <= _169;
    end
    assign _2736 = 8'b01011100;
    assign _2737 = _616 == _2736;
    assign _2735 = _565 & _570;
    assign _2738 = _2735 & _2737;
    assign _2742 = _2738 ? _599 : _2741;
    assign _2733 = _609 == _2736;
    assign _2731 = _565 & _580;
    assign _2734 = _2731 & _2733;
    assign _2743 = _2734 ? _583 : _2742;
    assign _170 = _2743;
    always @(posedge _539) begin
        if (_537)
            _2741 <= _567;
        else
            _2741 <= _170;
    end
    assign _2749 = 8'b01011011;
    assign _2750 = _616 == _2749;
    assign _2748 = _565 & _570;
    assign _2751 = _2748 & _2750;
    assign _2755 = _2751 ? _599 : _2754;
    assign _2746 = _609 == _2749;
    assign _2744 = _565 & _580;
    assign _2747 = _2744 & _2746;
    assign _2756 = _2747 ? _583 : _2755;
    assign _171 = _2756;
    always @(posedge _539) begin
        if (_537)
            _2754 <= _567;
        else
            _2754 <= _171;
    end
    assign _2762 = 8'b01011010;
    assign _2763 = _616 == _2762;
    assign _2761 = _565 & _570;
    assign _2764 = _2761 & _2763;
    assign _2768 = _2764 ? _599 : _2767;
    assign _2759 = _609 == _2762;
    assign _2757 = _565 & _580;
    assign _2760 = _2757 & _2759;
    assign _2769 = _2760 ? _583 : _2768;
    assign _172 = _2769;
    always @(posedge _539) begin
        if (_537)
            _2767 <= _567;
        else
            _2767 <= _172;
    end
    assign _2775 = 8'b01011001;
    assign _2776 = _616 == _2775;
    assign _2774 = _565 & _570;
    assign _2777 = _2774 & _2776;
    assign _2781 = _2777 ? _599 : _2780;
    assign _2772 = _609 == _2775;
    assign _2770 = _565 & _580;
    assign _2773 = _2770 & _2772;
    assign _2782 = _2773 ? _583 : _2781;
    assign _173 = _2782;
    always @(posedge _539) begin
        if (_537)
            _2780 <= _567;
        else
            _2780 <= _173;
    end
    assign _2788 = 8'b01011000;
    assign _2789 = _616 == _2788;
    assign _2787 = _565 & _570;
    assign _2790 = _2787 & _2789;
    assign _2794 = _2790 ? _599 : _2793;
    assign _2785 = _609 == _2788;
    assign _2783 = _565 & _580;
    assign _2786 = _2783 & _2785;
    assign _2795 = _2786 ? _583 : _2794;
    assign _174 = _2795;
    always @(posedge _539) begin
        if (_537)
            _2793 <= _567;
        else
            _2793 <= _174;
    end
    assign _2801 = 8'b01010111;
    assign _2802 = _616 == _2801;
    assign _2800 = _565 & _570;
    assign _2803 = _2800 & _2802;
    assign _2807 = _2803 ? _599 : _2806;
    assign _2798 = _609 == _2801;
    assign _2796 = _565 & _580;
    assign _2799 = _2796 & _2798;
    assign _2808 = _2799 ? _583 : _2807;
    assign _175 = _2808;
    always @(posedge _539) begin
        if (_537)
            _2806 <= _567;
        else
            _2806 <= _175;
    end
    assign _2814 = 8'b01010110;
    assign _2815 = _616 == _2814;
    assign _2813 = _565 & _570;
    assign _2816 = _2813 & _2815;
    assign _2820 = _2816 ? _599 : _2819;
    assign _2811 = _609 == _2814;
    assign _2809 = _565 & _580;
    assign _2812 = _2809 & _2811;
    assign _2821 = _2812 ? _583 : _2820;
    assign _176 = _2821;
    always @(posedge _539) begin
        if (_537)
            _2819 <= _567;
        else
            _2819 <= _176;
    end
    assign _2827 = 8'b01010101;
    assign _2828 = _616 == _2827;
    assign _2826 = _565 & _570;
    assign _2829 = _2826 & _2828;
    assign _2833 = _2829 ? _599 : _2832;
    assign _2824 = _609 == _2827;
    assign _2822 = _565 & _580;
    assign _2825 = _2822 & _2824;
    assign _2834 = _2825 ? _583 : _2833;
    assign _177 = _2834;
    always @(posedge _539) begin
        if (_537)
            _2832 <= _567;
        else
            _2832 <= _177;
    end
    assign _2840 = 8'b01010100;
    assign _2841 = _616 == _2840;
    assign _2839 = _565 & _570;
    assign _2842 = _2839 & _2841;
    assign _2846 = _2842 ? _599 : _2845;
    assign _2837 = _609 == _2840;
    assign _2835 = _565 & _580;
    assign _2838 = _2835 & _2837;
    assign _2847 = _2838 ? _583 : _2846;
    assign _178 = _2847;
    always @(posedge _539) begin
        if (_537)
            _2845 <= _567;
        else
            _2845 <= _178;
    end
    assign _2853 = 8'b01010011;
    assign _2854 = _616 == _2853;
    assign _2852 = _565 & _570;
    assign _2855 = _2852 & _2854;
    assign _2859 = _2855 ? _599 : _2858;
    assign _2850 = _609 == _2853;
    assign _2848 = _565 & _580;
    assign _2851 = _2848 & _2850;
    assign _2860 = _2851 ? _583 : _2859;
    assign _179 = _2860;
    always @(posedge _539) begin
        if (_537)
            _2858 <= _567;
        else
            _2858 <= _179;
    end
    assign _2866 = 8'b01010010;
    assign _2867 = _616 == _2866;
    assign _2865 = _565 & _570;
    assign _2868 = _2865 & _2867;
    assign _2872 = _2868 ? _599 : _2871;
    assign _2863 = _609 == _2866;
    assign _2861 = _565 & _580;
    assign _2864 = _2861 & _2863;
    assign _2873 = _2864 ? _583 : _2872;
    assign _180 = _2873;
    always @(posedge _539) begin
        if (_537)
            _2871 <= _567;
        else
            _2871 <= _180;
    end
    assign _2879 = 8'b01010001;
    assign _2880 = _616 == _2879;
    assign _2878 = _565 & _570;
    assign _2881 = _2878 & _2880;
    assign _2885 = _2881 ? _599 : _2884;
    assign _2876 = _609 == _2879;
    assign _2874 = _565 & _580;
    assign _2877 = _2874 & _2876;
    assign _2886 = _2877 ? _583 : _2885;
    assign _181 = _2886;
    always @(posedge _539) begin
        if (_537)
            _2884 <= _567;
        else
            _2884 <= _181;
    end
    assign _2892 = 8'b01010000;
    assign _2893 = _616 == _2892;
    assign _2891 = _565 & _570;
    assign _2894 = _2891 & _2893;
    assign _2898 = _2894 ? _599 : _2897;
    assign _2889 = _609 == _2892;
    assign _2887 = _565 & _580;
    assign _2890 = _2887 & _2889;
    assign _2899 = _2890 ? _583 : _2898;
    assign _182 = _2899;
    always @(posedge _539) begin
        if (_537)
            _2897 <= _567;
        else
            _2897 <= _182;
    end
    assign _2905 = 8'b01001111;
    assign _2906 = _616 == _2905;
    assign _2904 = _565 & _570;
    assign _2907 = _2904 & _2906;
    assign _2911 = _2907 ? _599 : _2910;
    assign _2902 = _609 == _2905;
    assign _2900 = _565 & _580;
    assign _2903 = _2900 & _2902;
    assign _2912 = _2903 ? _583 : _2911;
    assign _183 = _2912;
    always @(posedge _539) begin
        if (_537)
            _2910 <= _567;
        else
            _2910 <= _183;
    end
    assign _2918 = 8'b01001110;
    assign _2919 = _616 == _2918;
    assign _2917 = _565 & _570;
    assign _2920 = _2917 & _2919;
    assign _2924 = _2920 ? _599 : _2923;
    assign _2915 = _609 == _2918;
    assign _2913 = _565 & _580;
    assign _2916 = _2913 & _2915;
    assign _2925 = _2916 ? _583 : _2924;
    assign _184 = _2925;
    always @(posedge _539) begin
        if (_537)
            _2923 <= _567;
        else
            _2923 <= _184;
    end
    assign _2931 = 8'b01001101;
    assign _2932 = _616 == _2931;
    assign _2930 = _565 & _570;
    assign _2933 = _2930 & _2932;
    assign _2937 = _2933 ? _599 : _2936;
    assign _2928 = _609 == _2931;
    assign _2926 = _565 & _580;
    assign _2929 = _2926 & _2928;
    assign _2938 = _2929 ? _583 : _2937;
    assign _185 = _2938;
    always @(posedge _539) begin
        if (_537)
            _2936 <= _567;
        else
            _2936 <= _185;
    end
    assign _2944 = 8'b01001100;
    assign _2945 = _616 == _2944;
    assign _2943 = _565 & _570;
    assign _2946 = _2943 & _2945;
    assign _2950 = _2946 ? _599 : _2949;
    assign _2941 = _609 == _2944;
    assign _2939 = _565 & _580;
    assign _2942 = _2939 & _2941;
    assign _2951 = _2942 ? _583 : _2950;
    assign _186 = _2951;
    always @(posedge _539) begin
        if (_537)
            _2949 <= _567;
        else
            _2949 <= _186;
    end
    assign _2957 = 8'b01001011;
    assign _2958 = _616 == _2957;
    assign _2956 = _565 & _570;
    assign _2959 = _2956 & _2958;
    assign _2963 = _2959 ? _599 : _2962;
    assign _2954 = _609 == _2957;
    assign _2952 = _565 & _580;
    assign _2955 = _2952 & _2954;
    assign _2964 = _2955 ? _583 : _2963;
    assign _187 = _2964;
    always @(posedge _539) begin
        if (_537)
            _2962 <= _567;
        else
            _2962 <= _187;
    end
    assign _2970 = 8'b01001010;
    assign _2971 = _616 == _2970;
    assign _2969 = _565 & _570;
    assign _2972 = _2969 & _2971;
    assign _2976 = _2972 ? _599 : _2975;
    assign _2967 = _609 == _2970;
    assign _2965 = _565 & _580;
    assign _2968 = _2965 & _2967;
    assign _2977 = _2968 ? _583 : _2976;
    assign _188 = _2977;
    always @(posedge _539) begin
        if (_537)
            _2975 <= _567;
        else
            _2975 <= _188;
    end
    assign _2983 = 8'b01001001;
    assign _2984 = _616 == _2983;
    assign _2982 = _565 & _570;
    assign _2985 = _2982 & _2984;
    assign _2989 = _2985 ? _599 : _2988;
    assign _2980 = _609 == _2983;
    assign _2978 = _565 & _580;
    assign _2981 = _2978 & _2980;
    assign _2990 = _2981 ? _583 : _2989;
    assign _189 = _2990;
    always @(posedge _539) begin
        if (_537)
            _2988 <= _567;
        else
            _2988 <= _189;
    end
    assign _2996 = 8'b01001000;
    assign _2997 = _616 == _2996;
    assign _2995 = _565 & _570;
    assign _2998 = _2995 & _2997;
    assign _3002 = _2998 ? _599 : _3001;
    assign _2993 = _609 == _2996;
    assign _2991 = _565 & _580;
    assign _2994 = _2991 & _2993;
    assign _3003 = _2994 ? _583 : _3002;
    assign _190 = _3003;
    always @(posedge _539) begin
        if (_537)
            _3001 <= _567;
        else
            _3001 <= _190;
    end
    assign _3009 = 8'b01000111;
    assign _3010 = _616 == _3009;
    assign _3008 = _565 & _570;
    assign _3011 = _3008 & _3010;
    assign _3015 = _3011 ? _599 : _3014;
    assign _3006 = _609 == _3009;
    assign _3004 = _565 & _580;
    assign _3007 = _3004 & _3006;
    assign _3016 = _3007 ? _583 : _3015;
    assign _191 = _3016;
    always @(posedge _539) begin
        if (_537)
            _3014 <= _567;
        else
            _3014 <= _191;
    end
    assign _3022 = 8'b01000110;
    assign _3023 = _616 == _3022;
    assign _3021 = _565 & _570;
    assign _3024 = _3021 & _3023;
    assign _3028 = _3024 ? _599 : _3027;
    assign _3019 = _609 == _3022;
    assign _3017 = _565 & _580;
    assign _3020 = _3017 & _3019;
    assign _3029 = _3020 ? _583 : _3028;
    assign _192 = _3029;
    always @(posedge _539) begin
        if (_537)
            _3027 <= _567;
        else
            _3027 <= _192;
    end
    assign _3035 = 8'b01000101;
    assign _3036 = _616 == _3035;
    assign _3034 = _565 & _570;
    assign _3037 = _3034 & _3036;
    assign _3041 = _3037 ? _599 : _3040;
    assign _3032 = _609 == _3035;
    assign _3030 = _565 & _580;
    assign _3033 = _3030 & _3032;
    assign _3042 = _3033 ? _583 : _3041;
    assign _193 = _3042;
    always @(posedge _539) begin
        if (_537)
            _3040 <= _567;
        else
            _3040 <= _193;
    end
    assign _3048 = 8'b01000100;
    assign _3049 = _616 == _3048;
    assign _3047 = _565 & _570;
    assign _3050 = _3047 & _3049;
    assign _3054 = _3050 ? _599 : _3053;
    assign _3045 = _609 == _3048;
    assign _3043 = _565 & _580;
    assign _3046 = _3043 & _3045;
    assign _3055 = _3046 ? _583 : _3054;
    assign _194 = _3055;
    always @(posedge _539) begin
        if (_537)
            _3053 <= _567;
        else
            _3053 <= _194;
    end
    assign _3061 = 8'b01000011;
    assign _3062 = _616 == _3061;
    assign _3060 = _565 & _570;
    assign _3063 = _3060 & _3062;
    assign _3067 = _3063 ? _599 : _3066;
    assign _3058 = _609 == _3061;
    assign _3056 = _565 & _580;
    assign _3059 = _3056 & _3058;
    assign _3068 = _3059 ? _583 : _3067;
    assign _195 = _3068;
    always @(posedge _539) begin
        if (_537)
            _3066 <= _567;
        else
            _3066 <= _195;
    end
    assign _3074 = 8'b01000010;
    assign _3075 = _616 == _3074;
    assign _3073 = _565 & _570;
    assign _3076 = _3073 & _3075;
    assign _3080 = _3076 ? _599 : _3079;
    assign _3071 = _609 == _3074;
    assign _3069 = _565 & _580;
    assign _3072 = _3069 & _3071;
    assign _3081 = _3072 ? _583 : _3080;
    assign _196 = _3081;
    always @(posedge _539) begin
        if (_537)
            _3079 <= _567;
        else
            _3079 <= _196;
    end
    assign _3087 = 8'b01000001;
    assign _3088 = _616 == _3087;
    assign _3086 = _565 & _570;
    assign _3089 = _3086 & _3088;
    assign _3093 = _3089 ? _599 : _3092;
    assign _3084 = _609 == _3087;
    assign _3082 = _565 & _580;
    assign _3085 = _3082 & _3084;
    assign _3094 = _3085 ? _583 : _3093;
    assign _197 = _3094;
    always @(posedge _539) begin
        if (_537)
            _3092 <= _567;
        else
            _3092 <= _197;
    end
    assign _3100 = 8'b01000000;
    assign _3101 = _616 == _3100;
    assign _3099 = _565 & _570;
    assign _3102 = _3099 & _3101;
    assign _3106 = _3102 ? _599 : _3105;
    assign _3097 = _609 == _3100;
    assign _3095 = _565 & _580;
    assign _3098 = _3095 & _3097;
    assign _3107 = _3098 ? _583 : _3106;
    assign _198 = _3107;
    always @(posedge _539) begin
        if (_537)
            _3105 <= _567;
        else
            _3105 <= _198;
    end
    assign _3113 = 8'b00111111;
    assign _3114 = _616 == _3113;
    assign _3112 = _565 & _570;
    assign _3115 = _3112 & _3114;
    assign _3119 = _3115 ? _599 : _3118;
    assign _3110 = _609 == _3113;
    assign _3108 = _565 & _580;
    assign _3111 = _3108 & _3110;
    assign _3120 = _3111 ? _583 : _3119;
    assign _199 = _3120;
    always @(posedge _539) begin
        if (_537)
            _3118 <= _567;
        else
            _3118 <= _199;
    end
    assign _3126 = 8'b00111110;
    assign _3127 = _616 == _3126;
    assign _3125 = _565 & _570;
    assign _3128 = _3125 & _3127;
    assign _3132 = _3128 ? _599 : _3131;
    assign _3123 = _609 == _3126;
    assign _3121 = _565 & _580;
    assign _3124 = _3121 & _3123;
    assign _3133 = _3124 ? _583 : _3132;
    assign _200 = _3133;
    always @(posedge _539) begin
        if (_537)
            _3131 <= _567;
        else
            _3131 <= _200;
    end
    assign _3139 = 8'b00111101;
    assign _3140 = _616 == _3139;
    assign _3138 = _565 & _570;
    assign _3141 = _3138 & _3140;
    assign _3145 = _3141 ? _599 : _3144;
    assign _3136 = _609 == _3139;
    assign _3134 = _565 & _580;
    assign _3137 = _3134 & _3136;
    assign _3146 = _3137 ? _583 : _3145;
    assign _201 = _3146;
    always @(posedge _539) begin
        if (_537)
            _3144 <= _567;
        else
            _3144 <= _201;
    end
    assign _3152 = 8'b00111100;
    assign _3153 = _616 == _3152;
    assign _3151 = _565 & _570;
    assign _3154 = _3151 & _3153;
    assign _3158 = _3154 ? _599 : _3157;
    assign _3149 = _609 == _3152;
    assign _3147 = _565 & _580;
    assign _3150 = _3147 & _3149;
    assign _3159 = _3150 ? _583 : _3158;
    assign _202 = _3159;
    always @(posedge _539) begin
        if (_537)
            _3157 <= _567;
        else
            _3157 <= _202;
    end
    assign _3165 = 8'b00111011;
    assign _3166 = _616 == _3165;
    assign _3164 = _565 & _570;
    assign _3167 = _3164 & _3166;
    assign _3171 = _3167 ? _599 : _3170;
    assign _3162 = _609 == _3165;
    assign _3160 = _565 & _580;
    assign _3163 = _3160 & _3162;
    assign _3172 = _3163 ? _583 : _3171;
    assign _203 = _3172;
    always @(posedge _539) begin
        if (_537)
            _3170 <= _567;
        else
            _3170 <= _203;
    end
    assign _3178 = 8'b00111010;
    assign _3179 = _616 == _3178;
    assign _3177 = _565 & _570;
    assign _3180 = _3177 & _3179;
    assign _3184 = _3180 ? _599 : _3183;
    assign _3175 = _609 == _3178;
    assign _3173 = _565 & _580;
    assign _3176 = _3173 & _3175;
    assign _3185 = _3176 ? _583 : _3184;
    assign _204 = _3185;
    always @(posedge _539) begin
        if (_537)
            _3183 <= _567;
        else
            _3183 <= _204;
    end
    assign _3191 = 8'b00111001;
    assign _3192 = _616 == _3191;
    assign _3190 = _565 & _570;
    assign _3193 = _3190 & _3192;
    assign _3197 = _3193 ? _599 : _3196;
    assign _3188 = _609 == _3191;
    assign _3186 = _565 & _580;
    assign _3189 = _3186 & _3188;
    assign _3198 = _3189 ? _583 : _3197;
    assign _205 = _3198;
    always @(posedge _539) begin
        if (_537)
            _3196 <= _567;
        else
            _3196 <= _205;
    end
    assign _3204 = 8'b00111000;
    assign _3205 = _616 == _3204;
    assign _3203 = _565 & _570;
    assign _3206 = _3203 & _3205;
    assign _3210 = _3206 ? _599 : _3209;
    assign _3201 = _609 == _3204;
    assign _3199 = _565 & _580;
    assign _3202 = _3199 & _3201;
    assign _3211 = _3202 ? _583 : _3210;
    assign _206 = _3211;
    always @(posedge _539) begin
        if (_537)
            _3209 <= _567;
        else
            _3209 <= _206;
    end
    assign _3217 = 8'b00110111;
    assign _3218 = _616 == _3217;
    assign _3216 = _565 & _570;
    assign _3219 = _3216 & _3218;
    assign _3223 = _3219 ? _599 : _3222;
    assign _3214 = _609 == _3217;
    assign _3212 = _565 & _580;
    assign _3215 = _3212 & _3214;
    assign _3224 = _3215 ? _583 : _3223;
    assign _207 = _3224;
    always @(posedge _539) begin
        if (_537)
            _3222 <= _567;
        else
            _3222 <= _207;
    end
    assign _3230 = 8'b00110110;
    assign _3231 = _616 == _3230;
    assign _3229 = _565 & _570;
    assign _3232 = _3229 & _3231;
    assign _3236 = _3232 ? _599 : _3235;
    assign _3227 = _609 == _3230;
    assign _3225 = _565 & _580;
    assign _3228 = _3225 & _3227;
    assign _3237 = _3228 ? _583 : _3236;
    assign _208 = _3237;
    always @(posedge _539) begin
        if (_537)
            _3235 <= _567;
        else
            _3235 <= _208;
    end
    assign _3243 = 8'b00110101;
    assign _3244 = _616 == _3243;
    assign _3242 = _565 & _570;
    assign _3245 = _3242 & _3244;
    assign _3249 = _3245 ? _599 : _3248;
    assign _3240 = _609 == _3243;
    assign _3238 = _565 & _580;
    assign _3241 = _3238 & _3240;
    assign _3250 = _3241 ? _583 : _3249;
    assign _209 = _3250;
    always @(posedge _539) begin
        if (_537)
            _3248 <= _567;
        else
            _3248 <= _209;
    end
    assign _3256 = 8'b00110100;
    assign _3257 = _616 == _3256;
    assign _3255 = _565 & _570;
    assign _3258 = _3255 & _3257;
    assign _3262 = _3258 ? _599 : _3261;
    assign _3253 = _609 == _3256;
    assign _3251 = _565 & _580;
    assign _3254 = _3251 & _3253;
    assign _3263 = _3254 ? _583 : _3262;
    assign _210 = _3263;
    always @(posedge _539) begin
        if (_537)
            _3261 <= _567;
        else
            _3261 <= _210;
    end
    assign _3269 = 8'b00110011;
    assign _3270 = _616 == _3269;
    assign _3268 = _565 & _570;
    assign _3271 = _3268 & _3270;
    assign _3275 = _3271 ? _599 : _3274;
    assign _3266 = _609 == _3269;
    assign _3264 = _565 & _580;
    assign _3267 = _3264 & _3266;
    assign _3276 = _3267 ? _583 : _3275;
    assign _211 = _3276;
    always @(posedge _539) begin
        if (_537)
            _3274 <= _567;
        else
            _3274 <= _211;
    end
    assign _3282 = 8'b00110010;
    assign _3283 = _616 == _3282;
    assign _3281 = _565 & _570;
    assign _3284 = _3281 & _3283;
    assign _3288 = _3284 ? _599 : _3287;
    assign _3279 = _609 == _3282;
    assign _3277 = _565 & _580;
    assign _3280 = _3277 & _3279;
    assign _3289 = _3280 ? _583 : _3288;
    assign _212 = _3289;
    always @(posedge _539) begin
        if (_537)
            _3287 <= _567;
        else
            _3287 <= _212;
    end
    assign _3295 = 8'b00110001;
    assign _3296 = _616 == _3295;
    assign _3294 = _565 & _570;
    assign _3297 = _3294 & _3296;
    assign _3301 = _3297 ? _599 : _3300;
    assign _3292 = _609 == _3295;
    assign _3290 = _565 & _580;
    assign _3293 = _3290 & _3292;
    assign _3302 = _3293 ? _583 : _3301;
    assign _213 = _3302;
    always @(posedge _539) begin
        if (_537)
            _3300 <= _567;
        else
            _3300 <= _213;
    end
    assign _3308 = 8'b00110000;
    assign _3309 = _616 == _3308;
    assign _3307 = _565 & _570;
    assign _3310 = _3307 & _3309;
    assign _3314 = _3310 ? _599 : _3313;
    assign _3305 = _609 == _3308;
    assign _3303 = _565 & _580;
    assign _3306 = _3303 & _3305;
    assign _3315 = _3306 ? _583 : _3314;
    assign _214 = _3315;
    always @(posedge _539) begin
        if (_537)
            _3313 <= _567;
        else
            _3313 <= _214;
    end
    assign _3321 = 8'b00101111;
    assign _3322 = _616 == _3321;
    assign _3320 = _565 & _570;
    assign _3323 = _3320 & _3322;
    assign _3327 = _3323 ? _599 : _3326;
    assign _3318 = _609 == _3321;
    assign _3316 = _565 & _580;
    assign _3319 = _3316 & _3318;
    assign _3328 = _3319 ? _583 : _3327;
    assign _215 = _3328;
    always @(posedge _539) begin
        if (_537)
            _3326 <= _567;
        else
            _3326 <= _215;
    end
    assign _3334 = 8'b00101110;
    assign _3335 = _616 == _3334;
    assign _3333 = _565 & _570;
    assign _3336 = _3333 & _3335;
    assign _3340 = _3336 ? _599 : _3339;
    assign _3331 = _609 == _3334;
    assign _3329 = _565 & _580;
    assign _3332 = _3329 & _3331;
    assign _3341 = _3332 ? _583 : _3340;
    assign _216 = _3341;
    always @(posedge _539) begin
        if (_537)
            _3339 <= _567;
        else
            _3339 <= _216;
    end
    assign _3347 = 8'b00101101;
    assign _3348 = _616 == _3347;
    assign _3346 = _565 & _570;
    assign _3349 = _3346 & _3348;
    assign _3353 = _3349 ? _599 : _3352;
    assign _3344 = _609 == _3347;
    assign _3342 = _565 & _580;
    assign _3345 = _3342 & _3344;
    assign _3354 = _3345 ? _583 : _3353;
    assign _217 = _3354;
    always @(posedge _539) begin
        if (_537)
            _3352 <= _567;
        else
            _3352 <= _217;
    end
    assign _3360 = 8'b00101100;
    assign _3361 = _616 == _3360;
    assign _3359 = _565 & _570;
    assign _3362 = _3359 & _3361;
    assign _3366 = _3362 ? _599 : _3365;
    assign _3357 = _609 == _3360;
    assign _3355 = _565 & _580;
    assign _3358 = _3355 & _3357;
    assign _3367 = _3358 ? _583 : _3366;
    assign _218 = _3367;
    always @(posedge _539) begin
        if (_537)
            _3365 <= _567;
        else
            _3365 <= _218;
    end
    assign _3373 = 8'b00101011;
    assign _3374 = _616 == _3373;
    assign _3372 = _565 & _570;
    assign _3375 = _3372 & _3374;
    assign _3379 = _3375 ? _599 : _3378;
    assign _3370 = _609 == _3373;
    assign _3368 = _565 & _580;
    assign _3371 = _3368 & _3370;
    assign _3380 = _3371 ? _583 : _3379;
    assign _219 = _3380;
    always @(posedge _539) begin
        if (_537)
            _3378 <= _567;
        else
            _3378 <= _219;
    end
    assign _3386 = 8'b00101010;
    assign _3387 = _616 == _3386;
    assign _3385 = _565 & _570;
    assign _3388 = _3385 & _3387;
    assign _3392 = _3388 ? _599 : _3391;
    assign _3383 = _609 == _3386;
    assign _3381 = _565 & _580;
    assign _3384 = _3381 & _3383;
    assign _3393 = _3384 ? _583 : _3392;
    assign _220 = _3393;
    always @(posedge _539) begin
        if (_537)
            _3391 <= _567;
        else
            _3391 <= _220;
    end
    assign _3399 = 8'b00101001;
    assign _3400 = _616 == _3399;
    assign _3398 = _565 & _570;
    assign _3401 = _3398 & _3400;
    assign _3405 = _3401 ? _599 : _3404;
    assign _3396 = _609 == _3399;
    assign _3394 = _565 & _580;
    assign _3397 = _3394 & _3396;
    assign _3406 = _3397 ? _583 : _3405;
    assign _221 = _3406;
    always @(posedge _539) begin
        if (_537)
            _3404 <= _567;
        else
            _3404 <= _221;
    end
    assign _3412 = 8'b00101000;
    assign _3413 = _616 == _3412;
    assign _3411 = _565 & _570;
    assign _3414 = _3411 & _3413;
    assign _3418 = _3414 ? _599 : _3417;
    assign _3409 = _609 == _3412;
    assign _3407 = _565 & _580;
    assign _3410 = _3407 & _3409;
    assign _3419 = _3410 ? _583 : _3418;
    assign _222 = _3419;
    always @(posedge _539) begin
        if (_537)
            _3417 <= _567;
        else
            _3417 <= _222;
    end
    assign _3425 = 8'b00100111;
    assign _3426 = _616 == _3425;
    assign _3424 = _565 & _570;
    assign _3427 = _3424 & _3426;
    assign _3431 = _3427 ? _599 : _3430;
    assign _3422 = _609 == _3425;
    assign _3420 = _565 & _580;
    assign _3423 = _3420 & _3422;
    assign _3432 = _3423 ? _583 : _3431;
    assign _223 = _3432;
    always @(posedge _539) begin
        if (_537)
            _3430 <= _567;
        else
            _3430 <= _223;
    end
    assign _3438 = 8'b00100110;
    assign _3439 = _616 == _3438;
    assign _3437 = _565 & _570;
    assign _3440 = _3437 & _3439;
    assign _3444 = _3440 ? _599 : _3443;
    assign _3435 = _609 == _3438;
    assign _3433 = _565 & _580;
    assign _3436 = _3433 & _3435;
    assign _3445 = _3436 ? _583 : _3444;
    assign _224 = _3445;
    always @(posedge _539) begin
        if (_537)
            _3443 <= _567;
        else
            _3443 <= _224;
    end
    assign _3451 = 8'b00100101;
    assign _3452 = _616 == _3451;
    assign _3450 = _565 & _570;
    assign _3453 = _3450 & _3452;
    assign _3457 = _3453 ? _599 : _3456;
    assign _3448 = _609 == _3451;
    assign _3446 = _565 & _580;
    assign _3449 = _3446 & _3448;
    assign _3458 = _3449 ? _583 : _3457;
    assign _225 = _3458;
    always @(posedge _539) begin
        if (_537)
            _3456 <= _567;
        else
            _3456 <= _225;
    end
    assign _3464 = 8'b00100100;
    assign _3465 = _616 == _3464;
    assign _3463 = _565 & _570;
    assign _3466 = _3463 & _3465;
    assign _3470 = _3466 ? _599 : _3469;
    assign _3461 = _609 == _3464;
    assign _3459 = _565 & _580;
    assign _3462 = _3459 & _3461;
    assign _3471 = _3462 ? _583 : _3470;
    assign _226 = _3471;
    always @(posedge _539) begin
        if (_537)
            _3469 <= _567;
        else
            _3469 <= _226;
    end
    assign _3477 = 8'b00100011;
    assign _3478 = _616 == _3477;
    assign _3476 = _565 & _570;
    assign _3479 = _3476 & _3478;
    assign _3483 = _3479 ? _599 : _3482;
    assign _3474 = _609 == _3477;
    assign _3472 = _565 & _580;
    assign _3475 = _3472 & _3474;
    assign _3484 = _3475 ? _583 : _3483;
    assign _227 = _3484;
    always @(posedge _539) begin
        if (_537)
            _3482 <= _567;
        else
            _3482 <= _227;
    end
    assign _3490 = 8'b00100010;
    assign _3491 = _616 == _3490;
    assign _3489 = _565 & _570;
    assign _3492 = _3489 & _3491;
    assign _3496 = _3492 ? _599 : _3495;
    assign _3487 = _609 == _3490;
    assign _3485 = _565 & _580;
    assign _3488 = _3485 & _3487;
    assign _3497 = _3488 ? _583 : _3496;
    assign _228 = _3497;
    always @(posedge _539) begin
        if (_537)
            _3495 <= _567;
        else
            _3495 <= _228;
    end
    assign _3503 = 8'b00100001;
    assign _3504 = _616 == _3503;
    assign _3502 = _565 & _570;
    assign _3505 = _3502 & _3504;
    assign _3509 = _3505 ? _599 : _3508;
    assign _3500 = _609 == _3503;
    assign _3498 = _565 & _580;
    assign _3501 = _3498 & _3500;
    assign _3510 = _3501 ? _583 : _3509;
    assign _229 = _3510;
    always @(posedge _539) begin
        if (_537)
            _3508 <= _567;
        else
            _3508 <= _229;
    end
    assign _3516 = 8'b00100000;
    assign _3517 = _616 == _3516;
    assign _3515 = _565 & _570;
    assign _3518 = _3515 & _3517;
    assign _3522 = _3518 ? _599 : _3521;
    assign _3513 = _609 == _3516;
    assign _3511 = _565 & _580;
    assign _3514 = _3511 & _3513;
    assign _3523 = _3514 ? _583 : _3522;
    assign _230 = _3523;
    always @(posedge _539) begin
        if (_537)
            _3521 <= _567;
        else
            _3521 <= _230;
    end
    assign _3529 = 8'b00011111;
    assign _3530 = _616 == _3529;
    assign _3528 = _565 & _570;
    assign _3531 = _3528 & _3530;
    assign _3535 = _3531 ? _599 : _3534;
    assign _3526 = _609 == _3529;
    assign _3524 = _565 & _580;
    assign _3527 = _3524 & _3526;
    assign _3536 = _3527 ? _583 : _3535;
    assign _231 = _3536;
    always @(posedge _539) begin
        if (_537)
            _3534 <= _567;
        else
            _3534 <= _231;
    end
    assign _3542 = 8'b00011110;
    assign _3543 = _616 == _3542;
    assign _3541 = _565 & _570;
    assign _3544 = _3541 & _3543;
    assign _3548 = _3544 ? _599 : _3547;
    assign _3539 = _609 == _3542;
    assign _3537 = _565 & _580;
    assign _3540 = _3537 & _3539;
    assign _3549 = _3540 ? _583 : _3548;
    assign _232 = _3549;
    always @(posedge _539) begin
        if (_537)
            _3547 <= _567;
        else
            _3547 <= _232;
    end
    assign _3555 = 8'b00011101;
    assign _3556 = _616 == _3555;
    assign _3554 = _565 & _570;
    assign _3557 = _3554 & _3556;
    assign _3561 = _3557 ? _599 : _3560;
    assign _3552 = _609 == _3555;
    assign _3550 = _565 & _580;
    assign _3553 = _3550 & _3552;
    assign _3562 = _3553 ? _583 : _3561;
    assign _233 = _3562;
    always @(posedge _539) begin
        if (_537)
            _3560 <= _567;
        else
            _3560 <= _233;
    end
    assign _3568 = 8'b00011100;
    assign _3569 = _616 == _3568;
    assign _3567 = _565 & _570;
    assign _3570 = _3567 & _3569;
    assign _3574 = _3570 ? _599 : _3573;
    assign _3565 = _609 == _3568;
    assign _3563 = _565 & _580;
    assign _3566 = _3563 & _3565;
    assign _3575 = _3566 ? _583 : _3574;
    assign _234 = _3575;
    always @(posedge _539) begin
        if (_537)
            _3573 <= _567;
        else
            _3573 <= _234;
    end
    assign _3581 = 8'b00011011;
    assign _3582 = _616 == _3581;
    assign _3580 = _565 & _570;
    assign _3583 = _3580 & _3582;
    assign _3587 = _3583 ? _599 : _3586;
    assign _3578 = _609 == _3581;
    assign _3576 = _565 & _580;
    assign _3579 = _3576 & _3578;
    assign _3588 = _3579 ? _583 : _3587;
    assign _235 = _3588;
    always @(posedge _539) begin
        if (_537)
            _3586 <= _567;
        else
            _3586 <= _235;
    end
    assign _3594 = 8'b00011010;
    assign _3595 = _616 == _3594;
    assign _3593 = _565 & _570;
    assign _3596 = _3593 & _3595;
    assign _3600 = _3596 ? _599 : _3599;
    assign _3591 = _609 == _3594;
    assign _3589 = _565 & _580;
    assign _3592 = _3589 & _3591;
    assign _3601 = _3592 ? _583 : _3600;
    assign _236 = _3601;
    always @(posedge _539) begin
        if (_537)
            _3599 <= _567;
        else
            _3599 <= _236;
    end
    assign _3607 = 8'b00011001;
    assign _3608 = _616 == _3607;
    assign _3606 = _565 & _570;
    assign _3609 = _3606 & _3608;
    assign _3613 = _3609 ? _599 : _3612;
    assign _3604 = _609 == _3607;
    assign _3602 = _565 & _580;
    assign _3605 = _3602 & _3604;
    assign _3614 = _3605 ? _583 : _3613;
    assign _237 = _3614;
    always @(posedge _539) begin
        if (_537)
            _3612 <= _567;
        else
            _3612 <= _237;
    end
    assign _3620 = 8'b00011000;
    assign _3621 = _616 == _3620;
    assign _3619 = _565 & _570;
    assign _3622 = _3619 & _3621;
    assign _3626 = _3622 ? _599 : _3625;
    assign _3617 = _609 == _3620;
    assign _3615 = _565 & _580;
    assign _3618 = _3615 & _3617;
    assign _3627 = _3618 ? _583 : _3626;
    assign _238 = _3627;
    always @(posedge _539) begin
        if (_537)
            _3625 <= _567;
        else
            _3625 <= _238;
    end
    assign _3633 = 8'b00010111;
    assign _3634 = _616 == _3633;
    assign _3632 = _565 & _570;
    assign _3635 = _3632 & _3634;
    assign _3639 = _3635 ? _599 : _3638;
    assign _3630 = _609 == _3633;
    assign _3628 = _565 & _580;
    assign _3631 = _3628 & _3630;
    assign _3640 = _3631 ? _583 : _3639;
    assign _239 = _3640;
    always @(posedge _539) begin
        if (_537)
            _3638 <= _567;
        else
            _3638 <= _239;
    end
    assign _3646 = 8'b00010110;
    assign _3647 = _616 == _3646;
    assign _3645 = _565 & _570;
    assign _3648 = _3645 & _3647;
    assign _3652 = _3648 ? _599 : _3651;
    assign _3643 = _609 == _3646;
    assign _3641 = _565 & _580;
    assign _3644 = _3641 & _3643;
    assign _3653 = _3644 ? _583 : _3652;
    assign _240 = _3653;
    always @(posedge _539) begin
        if (_537)
            _3651 <= _567;
        else
            _3651 <= _240;
    end
    assign _3659 = 8'b00010101;
    assign _3660 = _616 == _3659;
    assign _3658 = _565 & _570;
    assign _3661 = _3658 & _3660;
    assign _3665 = _3661 ? _599 : _3664;
    assign _3656 = _609 == _3659;
    assign _3654 = _565 & _580;
    assign _3657 = _3654 & _3656;
    assign _3666 = _3657 ? _583 : _3665;
    assign _241 = _3666;
    always @(posedge _539) begin
        if (_537)
            _3664 <= _567;
        else
            _3664 <= _241;
    end
    assign _3672 = 8'b00010100;
    assign _3673 = _616 == _3672;
    assign _3671 = _565 & _570;
    assign _3674 = _3671 & _3673;
    assign _3678 = _3674 ? _599 : _3677;
    assign _3669 = _609 == _3672;
    assign _3667 = _565 & _580;
    assign _3670 = _3667 & _3669;
    assign _3679 = _3670 ? _583 : _3678;
    assign _242 = _3679;
    always @(posedge _539) begin
        if (_537)
            _3677 <= _567;
        else
            _3677 <= _242;
    end
    assign _3685 = 8'b00010011;
    assign _3686 = _616 == _3685;
    assign _3684 = _565 & _570;
    assign _3687 = _3684 & _3686;
    assign _3691 = _3687 ? _599 : _3690;
    assign _3682 = _609 == _3685;
    assign _3680 = _565 & _580;
    assign _3683 = _3680 & _3682;
    assign _3692 = _3683 ? _583 : _3691;
    assign _243 = _3692;
    always @(posedge _539) begin
        if (_537)
            _3690 <= _567;
        else
            _3690 <= _243;
    end
    assign _3698 = 8'b00010010;
    assign _3699 = _616 == _3698;
    assign _3697 = _565 & _570;
    assign _3700 = _3697 & _3699;
    assign _3704 = _3700 ? _599 : _3703;
    assign _3695 = _609 == _3698;
    assign _3693 = _565 & _580;
    assign _3696 = _3693 & _3695;
    assign _3705 = _3696 ? _583 : _3704;
    assign _244 = _3705;
    always @(posedge _539) begin
        if (_537)
            _3703 <= _567;
        else
            _3703 <= _244;
    end
    assign _3711 = 8'b00010001;
    assign _3712 = _616 == _3711;
    assign _3710 = _565 & _570;
    assign _3713 = _3710 & _3712;
    assign _3717 = _3713 ? _599 : _3716;
    assign _3708 = _609 == _3711;
    assign _3706 = _565 & _580;
    assign _3709 = _3706 & _3708;
    assign _3718 = _3709 ? _583 : _3717;
    assign _245 = _3718;
    always @(posedge _539) begin
        if (_537)
            _3716 <= _567;
        else
            _3716 <= _245;
    end
    assign _3724 = 8'b00010000;
    assign _3725 = _616 == _3724;
    assign _3723 = _565 & _570;
    assign _3726 = _3723 & _3725;
    assign _3730 = _3726 ? _599 : _3729;
    assign _3721 = _609 == _3724;
    assign _3719 = _565 & _580;
    assign _3722 = _3719 & _3721;
    assign _3731 = _3722 ? _583 : _3730;
    assign _246 = _3731;
    always @(posedge _539) begin
        if (_537)
            _3729 <= _567;
        else
            _3729 <= _246;
    end
    assign _3737 = 8'b00001111;
    assign _3738 = _616 == _3737;
    assign _3736 = _565 & _570;
    assign _3739 = _3736 & _3738;
    assign _3743 = _3739 ? _599 : _3742;
    assign _3734 = _609 == _3737;
    assign _3732 = _565 & _580;
    assign _3735 = _3732 & _3734;
    assign _3744 = _3735 ? _583 : _3743;
    assign _247 = _3744;
    always @(posedge _539) begin
        if (_537)
            _3742 <= _567;
        else
            _3742 <= _247;
    end
    assign _3750 = 8'b00001110;
    assign _3751 = _616 == _3750;
    assign _3749 = _565 & _570;
    assign _3752 = _3749 & _3751;
    assign _3756 = _3752 ? _599 : _3755;
    assign _3747 = _609 == _3750;
    assign _3745 = _565 & _580;
    assign _3748 = _3745 & _3747;
    assign _3757 = _3748 ? _583 : _3756;
    assign _248 = _3757;
    always @(posedge _539) begin
        if (_537)
            _3755 <= _567;
        else
            _3755 <= _248;
    end
    assign _3763 = 8'b00001101;
    assign _3764 = _616 == _3763;
    assign _3762 = _565 & _570;
    assign _3765 = _3762 & _3764;
    assign _3769 = _3765 ? _599 : _3768;
    assign _3760 = _609 == _3763;
    assign _3758 = _565 & _580;
    assign _3761 = _3758 & _3760;
    assign _3770 = _3761 ? _583 : _3769;
    assign _249 = _3770;
    always @(posedge _539) begin
        if (_537)
            _3768 <= _567;
        else
            _3768 <= _249;
    end
    assign _3776 = 8'b00001100;
    assign _3777 = _616 == _3776;
    assign _3775 = _565 & _570;
    assign _3778 = _3775 & _3777;
    assign _3782 = _3778 ? _599 : _3781;
    assign _3773 = _609 == _3776;
    assign _3771 = _565 & _580;
    assign _3774 = _3771 & _3773;
    assign _3783 = _3774 ? _583 : _3782;
    assign _250 = _3783;
    always @(posedge _539) begin
        if (_537)
            _3781 <= _567;
        else
            _3781 <= _250;
    end
    assign _3789 = 8'b00001011;
    assign _3790 = _616 == _3789;
    assign _3788 = _565 & _570;
    assign _3791 = _3788 & _3790;
    assign _3795 = _3791 ? _599 : _3794;
    assign _3786 = _609 == _3789;
    assign _3784 = _565 & _580;
    assign _3787 = _3784 & _3786;
    assign _3796 = _3787 ? _583 : _3795;
    assign _251 = _3796;
    always @(posedge _539) begin
        if (_537)
            _3794 <= _567;
        else
            _3794 <= _251;
    end
    assign _3802 = 8'b00001010;
    assign _3803 = _616 == _3802;
    assign _3801 = _565 & _570;
    assign _3804 = _3801 & _3803;
    assign _3808 = _3804 ? _599 : _3807;
    assign _3799 = _609 == _3802;
    assign _3797 = _565 & _580;
    assign _3800 = _3797 & _3799;
    assign _3809 = _3800 ? _583 : _3808;
    assign _252 = _3809;
    always @(posedge _539) begin
        if (_537)
            _3807 <= _567;
        else
            _3807 <= _252;
    end
    assign _3815 = 8'b00001001;
    assign _3816 = _616 == _3815;
    assign _3814 = _565 & _570;
    assign _3817 = _3814 & _3816;
    assign _3821 = _3817 ? _599 : _3820;
    assign _3812 = _609 == _3815;
    assign _3810 = _565 & _580;
    assign _3813 = _3810 & _3812;
    assign _3822 = _3813 ? _583 : _3821;
    assign _253 = _3822;
    always @(posedge _539) begin
        if (_537)
            _3820 <= _567;
        else
            _3820 <= _253;
    end
    assign _3828 = 8'b00001000;
    assign _3829 = _616 == _3828;
    assign _3827 = _565 & _570;
    assign _3830 = _3827 & _3829;
    assign _3834 = _3830 ? _599 : _3833;
    assign _3825 = _609 == _3828;
    assign _3823 = _565 & _580;
    assign _3826 = _3823 & _3825;
    assign _3835 = _3826 ? _583 : _3834;
    assign _254 = _3835;
    always @(posedge _539) begin
        if (_537)
            _3833 <= _567;
        else
            _3833 <= _254;
    end
    assign _3841 = 8'b00000111;
    assign _3842 = _616 == _3841;
    assign _3840 = _565 & _570;
    assign _3843 = _3840 & _3842;
    assign _3847 = _3843 ? _599 : _3846;
    assign _3838 = _609 == _3841;
    assign _3836 = _565 & _580;
    assign _3839 = _3836 & _3838;
    assign _3848 = _3839 ? _583 : _3847;
    assign _255 = _3848;
    always @(posedge _539) begin
        if (_537)
            _3846 <= _567;
        else
            _3846 <= _255;
    end
    assign _3854 = 8'b00000110;
    assign _3855 = _616 == _3854;
    assign _3853 = _565 & _570;
    assign _3856 = _3853 & _3855;
    assign _3860 = _3856 ? _599 : _3859;
    assign _3851 = _609 == _3854;
    assign _3849 = _565 & _580;
    assign _3852 = _3849 & _3851;
    assign _3861 = _3852 ? _583 : _3860;
    assign _256 = _3861;
    always @(posedge _539) begin
        if (_537)
            _3859 <= _567;
        else
            _3859 <= _256;
    end
    assign _3867 = 8'b00000101;
    assign _3868 = _616 == _3867;
    assign _3866 = _565 & _570;
    assign _3869 = _3866 & _3868;
    assign _3873 = _3869 ? _599 : _3872;
    assign _3864 = _609 == _3867;
    assign _3862 = _565 & _580;
    assign _3865 = _3862 & _3864;
    assign _3874 = _3865 ? _583 : _3873;
    assign _257 = _3874;
    always @(posedge _539) begin
        if (_537)
            _3872 <= _567;
        else
            _3872 <= _257;
    end
    assign _3880 = 8'b00000100;
    assign _3881 = _616 == _3880;
    assign _3879 = _565 & _570;
    assign _3882 = _3879 & _3881;
    assign _3886 = _3882 ? _599 : _3885;
    assign _3877 = _609 == _3880;
    assign _3875 = _565 & _580;
    assign _3878 = _3875 & _3877;
    assign _3887 = _3878 ? _583 : _3886;
    assign _258 = _3887;
    always @(posedge _539) begin
        if (_537)
            _3885 <= _567;
        else
            _3885 <= _258;
    end
    assign _3893 = 8'b00000011;
    assign _3894 = _616 == _3893;
    assign _3892 = _565 & _570;
    assign _3895 = _3892 & _3894;
    assign _3899 = _3895 ? _599 : _3898;
    assign _3890 = _609 == _3893;
    assign _3888 = _565 & _580;
    assign _3891 = _3888 & _3890;
    assign _3900 = _3891 ? _583 : _3899;
    assign _259 = _3900;
    always @(posedge _539) begin
        if (_537)
            _3898 <= _567;
        else
            _3898 <= _259;
    end
    assign _3906 = 8'b00000010;
    assign _3907 = _616 == _3906;
    assign _3905 = _565 & _570;
    assign _3908 = _3905 & _3907;
    assign _3912 = _3908 ? _599 : _3911;
    assign _3903 = _609 == _3906;
    assign _3901 = _565 & _580;
    assign _3904 = _3901 & _3903;
    assign _3913 = _3904 ? _583 : _3912;
    assign _260 = _3913;
    always @(posedge _539) begin
        if (_537)
            _3911 <= _567;
        else
            _3911 <= _260;
    end
    assign _3919 = 8'b00000001;
    assign _3920 = _616 == _3919;
    assign _3918 = _565 & _570;
    assign _3921 = _3918 & _3920;
    assign _3925 = _3921 ? _599 : _3924;
    assign _3916 = _609 == _3919;
    assign _3914 = _565 & _580;
    assign _3917 = _3914 & _3916;
    assign _3926 = _3917 ? _583 : _3925;
    assign _261 = _3926;
    always @(posedge _539) begin
        if (_537)
            _3924 <= _567;
        else
            _3924 <= _261;
    end
    assign _3927 = _565 ? _599 : _583;
    assign _3929 = _548 ? _567 : _3927;
    assign _262 = _3929;
    always @(posedge _539) begin
        if (_537)
            _583 <= _567;
        else
            _583 <= _262;
    end
    assign _598 = _580 ? _529 : _583;
    assign _599 = _588 ? _529 : _598;
    assign _3935 = 8'b00000000;
    assign _3936 = _616 == _3935;
    assign _3934 = _565 & _570;
    assign _3937 = _3934 & _3936;
    assign _3941 = _3937 ? _599 : _3940;
    assign _3932 = _609 == _3935;
    assign _3930 = _565 & _580;
    assign _3933 = _3930 & _3932;
    assign _3942 = _3933 ? _583 : _3941;
    assign _263 = _3942;
    always @(posedge _539) begin
        if (_537)
            _3940 <= _567;
        else
            _3940 <= _263;
    end
    always @* begin
        case (_7285)
        0:
            _7343 <= _3940;
        1:
            _7343 <= _3924;
        2:
            _7343 <= _3911;
        3:
            _7343 <= _3898;
        4:
            _7343 <= _3885;
        5:
            _7343 <= _3872;
        6:
            _7343 <= _3859;
        7:
            _7343 <= _3846;
        8:
            _7343 <= _3833;
        9:
            _7343 <= _3820;
        10:
            _7343 <= _3807;
        11:
            _7343 <= _3794;
        12:
            _7343 <= _3781;
        13:
            _7343 <= _3768;
        14:
            _7343 <= _3755;
        15:
            _7343 <= _3742;
        16:
            _7343 <= _3729;
        17:
            _7343 <= _3716;
        18:
            _7343 <= _3703;
        19:
            _7343 <= _3690;
        20:
            _7343 <= _3677;
        21:
            _7343 <= _3664;
        22:
            _7343 <= _3651;
        23:
            _7343 <= _3638;
        24:
            _7343 <= _3625;
        25:
            _7343 <= _3612;
        26:
            _7343 <= _3599;
        27:
            _7343 <= _3586;
        28:
            _7343 <= _3573;
        29:
            _7343 <= _3560;
        30:
            _7343 <= _3547;
        31:
            _7343 <= _3534;
        32:
            _7343 <= _3521;
        33:
            _7343 <= _3508;
        34:
            _7343 <= _3495;
        35:
            _7343 <= _3482;
        36:
            _7343 <= _3469;
        37:
            _7343 <= _3456;
        38:
            _7343 <= _3443;
        39:
            _7343 <= _3430;
        40:
            _7343 <= _3417;
        41:
            _7343 <= _3404;
        42:
            _7343 <= _3391;
        43:
            _7343 <= _3378;
        44:
            _7343 <= _3365;
        45:
            _7343 <= _3352;
        46:
            _7343 <= _3339;
        47:
            _7343 <= _3326;
        48:
            _7343 <= _3313;
        49:
            _7343 <= _3300;
        50:
            _7343 <= _3287;
        51:
            _7343 <= _3274;
        52:
            _7343 <= _3261;
        53:
            _7343 <= _3248;
        54:
            _7343 <= _3235;
        55:
            _7343 <= _3222;
        56:
            _7343 <= _3209;
        57:
            _7343 <= _3196;
        58:
            _7343 <= _3183;
        59:
            _7343 <= _3170;
        60:
            _7343 <= _3157;
        61:
            _7343 <= _3144;
        62:
            _7343 <= _3131;
        63:
            _7343 <= _3118;
        64:
            _7343 <= _3105;
        65:
            _7343 <= _3092;
        66:
            _7343 <= _3079;
        67:
            _7343 <= _3066;
        68:
            _7343 <= _3053;
        69:
            _7343 <= _3040;
        70:
            _7343 <= _3027;
        71:
            _7343 <= _3014;
        72:
            _7343 <= _3001;
        73:
            _7343 <= _2988;
        74:
            _7343 <= _2975;
        75:
            _7343 <= _2962;
        76:
            _7343 <= _2949;
        77:
            _7343 <= _2936;
        78:
            _7343 <= _2923;
        79:
            _7343 <= _2910;
        80:
            _7343 <= _2897;
        81:
            _7343 <= _2884;
        82:
            _7343 <= _2871;
        83:
            _7343 <= _2858;
        84:
            _7343 <= _2845;
        85:
            _7343 <= _2832;
        86:
            _7343 <= _2819;
        87:
            _7343 <= _2806;
        88:
            _7343 <= _2793;
        89:
            _7343 <= _2780;
        90:
            _7343 <= _2767;
        91:
            _7343 <= _2754;
        92:
            _7343 <= _2741;
        93:
            _7343 <= _2728;
        94:
            _7343 <= _2715;
        95:
            _7343 <= _2702;
        96:
            _7343 <= _2689;
        97:
            _7343 <= _2676;
        98:
            _7343 <= _2663;
        99:
            _7343 <= _2650;
        100:
            _7343 <= _2637;
        101:
            _7343 <= _2624;
        102:
            _7343 <= _2611;
        103:
            _7343 <= _2598;
        104:
            _7343 <= _2585;
        105:
            _7343 <= _2572;
        106:
            _7343 <= _2559;
        107:
            _7343 <= _2546;
        108:
            _7343 <= _2533;
        109:
            _7343 <= _2520;
        110:
            _7343 <= _2507;
        111:
            _7343 <= _2494;
        112:
            _7343 <= _2481;
        113:
            _7343 <= _2468;
        114:
            _7343 <= _2455;
        115:
            _7343 <= _2442;
        116:
            _7343 <= _2429;
        117:
            _7343 <= _2416;
        118:
            _7343 <= _2403;
        119:
            _7343 <= _2390;
        120:
            _7343 <= _2377;
        121:
            _7343 <= _2364;
        122:
            _7343 <= _2351;
        123:
            _7343 <= _2338;
        124:
            _7343 <= _2325;
        125:
            _7343 <= _2312;
        126:
            _7343 <= _2299;
        127:
            _7343 <= _2286;
        128:
            _7343 <= _2273;
        129:
            _7343 <= _2260;
        130:
            _7343 <= _2247;
        131:
            _7343 <= _2234;
        132:
            _7343 <= _2221;
        133:
            _7343 <= _2208;
        134:
            _7343 <= _2195;
        135:
            _7343 <= _2182;
        136:
            _7343 <= _2169;
        137:
            _7343 <= _2156;
        138:
            _7343 <= _2143;
        139:
            _7343 <= _2130;
        140:
            _7343 <= _2117;
        141:
            _7343 <= _2104;
        142:
            _7343 <= _2091;
        143:
            _7343 <= _2078;
        144:
            _7343 <= _2065;
        145:
            _7343 <= _2052;
        146:
            _7343 <= _2039;
        147:
            _7343 <= _2026;
        148:
            _7343 <= _2013;
        149:
            _7343 <= _2000;
        150:
            _7343 <= _1987;
        151:
            _7343 <= _1974;
        152:
            _7343 <= _1961;
        153:
            _7343 <= _1948;
        154:
            _7343 <= _1935;
        155:
            _7343 <= _1922;
        156:
            _7343 <= _1909;
        157:
            _7343 <= _1896;
        158:
            _7343 <= _1883;
        159:
            _7343 <= _1870;
        160:
            _7343 <= _1857;
        161:
            _7343 <= _1844;
        162:
            _7343 <= _1831;
        163:
            _7343 <= _1818;
        164:
            _7343 <= _1805;
        165:
            _7343 <= _1792;
        166:
            _7343 <= _1779;
        167:
            _7343 <= _1766;
        168:
            _7343 <= _1753;
        169:
            _7343 <= _1740;
        170:
            _7343 <= _1727;
        171:
            _7343 <= _1714;
        172:
            _7343 <= _1701;
        173:
            _7343 <= _1688;
        174:
            _7343 <= _1675;
        175:
            _7343 <= _1662;
        176:
            _7343 <= _1649;
        177:
            _7343 <= _1636;
        178:
            _7343 <= _1623;
        179:
            _7343 <= _1610;
        180:
            _7343 <= _1597;
        181:
            _7343 <= _1584;
        182:
            _7343 <= _1571;
        183:
            _7343 <= _1558;
        184:
            _7343 <= _1545;
        185:
            _7343 <= _1532;
        186:
            _7343 <= _1519;
        187:
            _7343 <= _1506;
        188:
            _7343 <= _1493;
        189:
            _7343 <= _1480;
        190:
            _7343 <= _1467;
        191:
            _7343 <= _1454;
        192:
            _7343 <= _1441;
        193:
            _7343 <= _1428;
        194:
            _7343 <= _1415;
        195:
            _7343 <= _1402;
        196:
            _7343 <= _1389;
        197:
            _7343 <= _1376;
        198:
            _7343 <= _1363;
        199:
            _7343 <= _1350;
        200:
            _7343 <= _1337;
        201:
            _7343 <= _1324;
        202:
            _7343 <= _1311;
        203:
            _7343 <= _1298;
        204:
            _7343 <= _1285;
        205:
            _7343 <= _1272;
        206:
            _7343 <= _1259;
        207:
            _7343 <= _1246;
        208:
            _7343 <= _1233;
        209:
            _7343 <= _1220;
        210:
            _7343 <= _1207;
        211:
            _7343 <= _1194;
        212:
            _7343 <= _1181;
        213:
            _7343 <= _1168;
        214:
            _7343 <= _1155;
        215:
            _7343 <= _1142;
        216:
            _7343 <= _1129;
        217:
            _7343 <= _1116;
        218:
            _7343 <= _1103;
        219:
            _7343 <= _1090;
        220:
            _7343 <= _1077;
        221:
            _7343 <= _1064;
        222:
            _7343 <= _1051;
        223:
            _7343 <= _1038;
        224:
            _7343 <= _1025;
        225:
            _7343 <= _1012;
        226:
            _7343 <= _999;
        227:
            _7343 <= _986;
        228:
            _7343 <= _973;
        229:
            _7343 <= _960;
        230:
            _7343 <= _947;
        231:
            _7343 <= _934;
        232:
            _7343 <= _921;
        233:
            _7343 <= _908;
        234:
            _7343 <= _895;
        235:
            _7343 <= _882;
        236:
            _7343 <= _869;
        237:
            _7343 <= _856;
        238:
            _7343 <= _843;
        239:
            _7343 <= _830;
        240:
            _7343 <= _817;
        241:
            _7343 <= _804;
        242:
            _7343 <= _791;
        243:
            _7343 <= _778;
        244:
            _7343 <= _765;
        245:
            _7343 <= _752;
        246:
            _7343 <= _739;
        247:
            _7343 <= _726;
        248:
            _7343 <= _713;
        249:
            _7343 <= _700;
        250:
            _7343 <= _687;
        251:
            _7343 <= _674;
        252:
            _7343 <= _661;
        253:
            _7343 <= _648;
        254:
            _7343 <= _635;
        default:
            _7343 <= _622;
        endcase
    end
    assign _7344 = _7282 < _7343;
    assign _7345 = ~ _7344;
    assign _7346 = _7278 & _7345;
    assign _7348 = _7346 & _7347;
    assign _7292 = _7275 - _3919;
    assign _7293 = _7278 ? _7292 : _3935;
    assign _7294 = _7285 < _7293;
    assign _3949 = _616 == _617;
    assign _3947 = _565 & _570;
    assign _3950 = _3947 & _3949;
    assign _3954 = _3950 ? _597 : _3953;
    assign _3945 = _609 == _617;
    assign _3943 = _565 & _580;
    assign _3946 = _3943 & _3945;
    assign _3955 = _3946 ? _577 : _3954;
    assign _264 = _3955;
    always @(posedge _539) begin
        if (_537)
            _3953 <= _567;
        else
            _3953 <= _264;
    end
    assign _3962 = _616 == _630;
    assign _3960 = _565 & _570;
    assign _3963 = _3960 & _3962;
    assign _3967 = _3963 ? _597 : _3966;
    assign _3958 = _609 == _630;
    assign _3956 = _565 & _580;
    assign _3959 = _3956 & _3958;
    assign _3968 = _3959 ? _577 : _3967;
    assign _265 = _3968;
    always @(posedge _539) begin
        if (_537)
            _3966 <= _567;
        else
            _3966 <= _265;
    end
    assign _3975 = _616 == _643;
    assign _3973 = _565 & _570;
    assign _3976 = _3973 & _3975;
    assign _3980 = _3976 ? _597 : _3979;
    assign _3971 = _609 == _643;
    assign _3969 = _565 & _580;
    assign _3972 = _3969 & _3971;
    assign _3981 = _3972 ? _577 : _3980;
    assign _266 = _3981;
    always @(posedge _539) begin
        if (_537)
            _3979 <= _567;
        else
            _3979 <= _266;
    end
    assign _3988 = _616 == _656;
    assign _3986 = _565 & _570;
    assign _3989 = _3986 & _3988;
    assign _3993 = _3989 ? _597 : _3992;
    assign _3984 = _609 == _656;
    assign _3982 = _565 & _580;
    assign _3985 = _3982 & _3984;
    assign _3994 = _3985 ? _577 : _3993;
    assign _267 = _3994;
    always @(posedge _539) begin
        if (_537)
            _3992 <= _567;
        else
            _3992 <= _267;
    end
    assign _4001 = _616 == _669;
    assign _3999 = _565 & _570;
    assign _4002 = _3999 & _4001;
    assign _4006 = _4002 ? _597 : _4005;
    assign _3997 = _609 == _669;
    assign _3995 = _565 & _580;
    assign _3998 = _3995 & _3997;
    assign _4007 = _3998 ? _577 : _4006;
    assign _268 = _4007;
    always @(posedge _539) begin
        if (_537)
            _4005 <= _567;
        else
            _4005 <= _268;
    end
    assign _4014 = _616 == _682;
    assign _4012 = _565 & _570;
    assign _4015 = _4012 & _4014;
    assign _4019 = _4015 ? _597 : _4018;
    assign _4010 = _609 == _682;
    assign _4008 = _565 & _580;
    assign _4011 = _4008 & _4010;
    assign _4020 = _4011 ? _577 : _4019;
    assign _269 = _4020;
    always @(posedge _539) begin
        if (_537)
            _4018 <= _567;
        else
            _4018 <= _269;
    end
    assign _4027 = _616 == _695;
    assign _4025 = _565 & _570;
    assign _4028 = _4025 & _4027;
    assign _4032 = _4028 ? _597 : _4031;
    assign _4023 = _609 == _695;
    assign _4021 = _565 & _580;
    assign _4024 = _4021 & _4023;
    assign _4033 = _4024 ? _577 : _4032;
    assign _270 = _4033;
    always @(posedge _539) begin
        if (_537)
            _4031 <= _567;
        else
            _4031 <= _270;
    end
    assign _4040 = _616 == _708;
    assign _4038 = _565 & _570;
    assign _4041 = _4038 & _4040;
    assign _4045 = _4041 ? _597 : _4044;
    assign _4036 = _609 == _708;
    assign _4034 = _565 & _580;
    assign _4037 = _4034 & _4036;
    assign _4046 = _4037 ? _577 : _4045;
    assign _271 = _4046;
    always @(posedge _539) begin
        if (_537)
            _4044 <= _567;
        else
            _4044 <= _271;
    end
    assign _4053 = _616 == _721;
    assign _4051 = _565 & _570;
    assign _4054 = _4051 & _4053;
    assign _4058 = _4054 ? _597 : _4057;
    assign _4049 = _609 == _721;
    assign _4047 = _565 & _580;
    assign _4050 = _4047 & _4049;
    assign _4059 = _4050 ? _577 : _4058;
    assign _272 = _4059;
    always @(posedge _539) begin
        if (_537)
            _4057 <= _567;
        else
            _4057 <= _272;
    end
    assign _4066 = _616 == _734;
    assign _4064 = _565 & _570;
    assign _4067 = _4064 & _4066;
    assign _4071 = _4067 ? _597 : _4070;
    assign _4062 = _609 == _734;
    assign _4060 = _565 & _580;
    assign _4063 = _4060 & _4062;
    assign _4072 = _4063 ? _577 : _4071;
    assign _273 = _4072;
    always @(posedge _539) begin
        if (_537)
            _4070 <= _567;
        else
            _4070 <= _273;
    end
    assign _4079 = _616 == _747;
    assign _4077 = _565 & _570;
    assign _4080 = _4077 & _4079;
    assign _4084 = _4080 ? _597 : _4083;
    assign _4075 = _609 == _747;
    assign _4073 = _565 & _580;
    assign _4076 = _4073 & _4075;
    assign _4085 = _4076 ? _577 : _4084;
    assign _274 = _4085;
    always @(posedge _539) begin
        if (_537)
            _4083 <= _567;
        else
            _4083 <= _274;
    end
    assign _4092 = _616 == _760;
    assign _4090 = _565 & _570;
    assign _4093 = _4090 & _4092;
    assign _4097 = _4093 ? _597 : _4096;
    assign _4088 = _609 == _760;
    assign _4086 = _565 & _580;
    assign _4089 = _4086 & _4088;
    assign _4098 = _4089 ? _577 : _4097;
    assign _275 = _4098;
    always @(posedge _539) begin
        if (_537)
            _4096 <= _567;
        else
            _4096 <= _275;
    end
    assign _4105 = _616 == _773;
    assign _4103 = _565 & _570;
    assign _4106 = _4103 & _4105;
    assign _4110 = _4106 ? _597 : _4109;
    assign _4101 = _609 == _773;
    assign _4099 = _565 & _580;
    assign _4102 = _4099 & _4101;
    assign _4111 = _4102 ? _577 : _4110;
    assign _276 = _4111;
    always @(posedge _539) begin
        if (_537)
            _4109 <= _567;
        else
            _4109 <= _276;
    end
    assign _4118 = _616 == _786;
    assign _4116 = _565 & _570;
    assign _4119 = _4116 & _4118;
    assign _4123 = _4119 ? _597 : _4122;
    assign _4114 = _609 == _786;
    assign _4112 = _565 & _580;
    assign _4115 = _4112 & _4114;
    assign _4124 = _4115 ? _577 : _4123;
    assign _277 = _4124;
    always @(posedge _539) begin
        if (_537)
            _4122 <= _567;
        else
            _4122 <= _277;
    end
    assign _4131 = _616 == _799;
    assign _4129 = _565 & _570;
    assign _4132 = _4129 & _4131;
    assign _4136 = _4132 ? _597 : _4135;
    assign _4127 = _609 == _799;
    assign _4125 = _565 & _580;
    assign _4128 = _4125 & _4127;
    assign _4137 = _4128 ? _577 : _4136;
    assign _278 = _4137;
    always @(posedge _539) begin
        if (_537)
            _4135 <= _567;
        else
            _4135 <= _278;
    end
    assign _4144 = _616 == _812;
    assign _4142 = _565 & _570;
    assign _4145 = _4142 & _4144;
    assign _4149 = _4145 ? _597 : _4148;
    assign _4140 = _609 == _812;
    assign _4138 = _565 & _580;
    assign _4141 = _4138 & _4140;
    assign _4150 = _4141 ? _577 : _4149;
    assign _279 = _4150;
    always @(posedge _539) begin
        if (_537)
            _4148 <= _567;
        else
            _4148 <= _279;
    end
    assign _4157 = _616 == _825;
    assign _4155 = _565 & _570;
    assign _4158 = _4155 & _4157;
    assign _4162 = _4158 ? _597 : _4161;
    assign _4153 = _609 == _825;
    assign _4151 = _565 & _580;
    assign _4154 = _4151 & _4153;
    assign _4163 = _4154 ? _577 : _4162;
    assign _280 = _4163;
    always @(posedge _539) begin
        if (_537)
            _4161 <= _567;
        else
            _4161 <= _280;
    end
    assign _4170 = _616 == _838;
    assign _4168 = _565 & _570;
    assign _4171 = _4168 & _4170;
    assign _4175 = _4171 ? _597 : _4174;
    assign _4166 = _609 == _838;
    assign _4164 = _565 & _580;
    assign _4167 = _4164 & _4166;
    assign _4176 = _4167 ? _577 : _4175;
    assign _281 = _4176;
    always @(posedge _539) begin
        if (_537)
            _4174 <= _567;
        else
            _4174 <= _281;
    end
    assign _4183 = _616 == _851;
    assign _4181 = _565 & _570;
    assign _4184 = _4181 & _4183;
    assign _4188 = _4184 ? _597 : _4187;
    assign _4179 = _609 == _851;
    assign _4177 = _565 & _580;
    assign _4180 = _4177 & _4179;
    assign _4189 = _4180 ? _577 : _4188;
    assign _282 = _4189;
    always @(posedge _539) begin
        if (_537)
            _4187 <= _567;
        else
            _4187 <= _282;
    end
    assign _4196 = _616 == _864;
    assign _4194 = _565 & _570;
    assign _4197 = _4194 & _4196;
    assign _4201 = _4197 ? _597 : _4200;
    assign _4192 = _609 == _864;
    assign _4190 = _565 & _580;
    assign _4193 = _4190 & _4192;
    assign _4202 = _4193 ? _577 : _4201;
    assign _283 = _4202;
    always @(posedge _539) begin
        if (_537)
            _4200 <= _567;
        else
            _4200 <= _283;
    end
    assign _4209 = _616 == _877;
    assign _4207 = _565 & _570;
    assign _4210 = _4207 & _4209;
    assign _4214 = _4210 ? _597 : _4213;
    assign _4205 = _609 == _877;
    assign _4203 = _565 & _580;
    assign _4206 = _4203 & _4205;
    assign _4215 = _4206 ? _577 : _4214;
    assign _284 = _4215;
    always @(posedge _539) begin
        if (_537)
            _4213 <= _567;
        else
            _4213 <= _284;
    end
    assign _4222 = _616 == _890;
    assign _4220 = _565 & _570;
    assign _4223 = _4220 & _4222;
    assign _4227 = _4223 ? _597 : _4226;
    assign _4218 = _609 == _890;
    assign _4216 = _565 & _580;
    assign _4219 = _4216 & _4218;
    assign _4228 = _4219 ? _577 : _4227;
    assign _285 = _4228;
    always @(posedge _539) begin
        if (_537)
            _4226 <= _567;
        else
            _4226 <= _285;
    end
    assign _4235 = _616 == _903;
    assign _4233 = _565 & _570;
    assign _4236 = _4233 & _4235;
    assign _4240 = _4236 ? _597 : _4239;
    assign _4231 = _609 == _903;
    assign _4229 = _565 & _580;
    assign _4232 = _4229 & _4231;
    assign _4241 = _4232 ? _577 : _4240;
    assign _286 = _4241;
    always @(posedge _539) begin
        if (_537)
            _4239 <= _567;
        else
            _4239 <= _286;
    end
    assign _4248 = _616 == _916;
    assign _4246 = _565 & _570;
    assign _4249 = _4246 & _4248;
    assign _4253 = _4249 ? _597 : _4252;
    assign _4244 = _609 == _916;
    assign _4242 = _565 & _580;
    assign _4245 = _4242 & _4244;
    assign _4254 = _4245 ? _577 : _4253;
    assign _287 = _4254;
    always @(posedge _539) begin
        if (_537)
            _4252 <= _567;
        else
            _4252 <= _287;
    end
    assign _4261 = _616 == _929;
    assign _4259 = _565 & _570;
    assign _4262 = _4259 & _4261;
    assign _4266 = _4262 ? _597 : _4265;
    assign _4257 = _609 == _929;
    assign _4255 = _565 & _580;
    assign _4258 = _4255 & _4257;
    assign _4267 = _4258 ? _577 : _4266;
    assign _288 = _4267;
    always @(posedge _539) begin
        if (_537)
            _4265 <= _567;
        else
            _4265 <= _288;
    end
    assign _4274 = _616 == _942;
    assign _4272 = _565 & _570;
    assign _4275 = _4272 & _4274;
    assign _4279 = _4275 ? _597 : _4278;
    assign _4270 = _609 == _942;
    assign _4268 = _565 & _580;
    assign _4271 = _4268 & _4270;
    assign _4280 = _4271 ? _577 : _4279;
    assign _289 = _4280;
    always @(posedge _539) begin
        if (_537)
            _4278 <= _567;
        else
            _4278 <= _289;
    end
    assign _4287 = _616 == _955;
    assign _4285 = _565 & _570;
    assign _4288 = _4285 & _4287;
    assign _4292 = _4288 ? _597 : _4291;
    assign _4283 = _609 == _955;
    assign _4281 = _565 & _580;
    assign _4284 = _4281 & _4283;
    assign _4293 = _4284 ? _577 : _4292;
    assign _290 = _4293;
    always @(posedge _539) begin
        if (_537)
            _4291 <= _567;
        else
            _4291 <= _290;
    end
    assign _4300 = _616 == _968;
    assign _4298 = _565 & _570;
    assign _4301 = _4298 & _4300;
    assign _4305 = _4301 ? _597 : _4304;
    assign _4296 = _609 == _968;
    assign _4294 = _565 & _580;
    assign _4297 = _4294 & _4296;
    assign _4306 = _4297 ? _577 : _4305;
    assign _291 = _4306;
    always @(posedge _539) begin
        if (_537)
            _4304 <= _567;
        else
            _4304 <= _291;
    end
    assign _4313 = _616 == _981;
    assign _4311 = _565 & _570;
    assign _4314 = _4311 & _4313;
    assign _4318 = _4314 ? _597 : _4317;
    assign _4309 = _609 == _981;
    assign _4307 = _565 & _580;
    assign _4310 = _4307 & _4309;
    assign _4319 = _4310 ? _577 : _4318;
    assign _292 = _4319;
    always @(posedge _539) begin
        if (_537)
            _4317 <= _567;
        else
            _4317 <= _292;
    end
    assign _4326 = _616 == _994;
    assign _4324 = _565 & _570;
    assign _4327 = _4324 & _4326;
    assign _4331 = _4327 ? _597 : _4330;
    assign _4322 = _609 == _994;
    assign _4320 = _565 & _580;
    assign _4323 = _4320 & _4322;
    assign _4332 = _4323 ? _577 : _4331;
    assign _293 = _4332;
    always @(posedge _539) begin
        if (_537)
            _4330 <= _567;
        else
            _4330 <= _293;
    end
    assign _4339 = _616 == _1007;
    assign _4337 = _565 & _570;
    assign _4340 = _4337 & _4339;
    assign _4344 = _4340 ? _597 : _4343;
    assign _4335 = _609 == _1007;
    assign _4333 = _565 & _580;
    assign _4336 = _4333 & _4335;
    assign _4345 = _4336 ? _577 : _4344;
    assign _294 = _4345;
    always @(posedge _539) begin
        if (_537)
            _4343 <= _567;
        else
            _4343 <= _294;
    end
    assign _4352 = _616 == _1020;
    assign _4350 = _565 & _570;
    assign _4353 = _4350 & _4352;
    assign _4357 = _4353 ? _597 : _4356;
    assign _4348 = _609 == _1020;
    assign _4346 = _565 & _580;
    assign _4349 = _4346 & _4348;
    assign _4358 = _4349 ? _577 : _4357;
    assign _295 = _4358;
    always @(posedge _539) begin
        if (_537)
            _4356 <= _567;
        else
            _4356 <= _295;
    end
    assign _4365 = _616 == _1033;
    assign _4363 = _565 & _570;
    assign _4366 = _4363 & _4365;
    assign _4370 = _4366 ? _597 : _4369;
    assign _4361 = _609 == _1033;
    assign _4359 = _565 & _580;
    assign _4362 = _4359 & _4361;
    assign _4371 = _4362 ? _577 : _4370;
    assign _296 = _4371;
    always @(posedge _539) begin
        if (_537)
            _4369 <= _567;
        else
            _4369 <= _296;
    end
    assign _4378 = _616 == _1046;
    assign _4376 = _565 & _570;
    assign _4379 = _4376 & _4378;
    assign _4383 = _4379 ? _597 : _4382;
    assign _4374 = _609 == _1046;
    assign _4372 = _565 & _580;
    assign _4375 = _4372 & _4374;
    assign _4384 = _4375 ? _577 : _4383;
    assign _297 = _4384;
    always @(posedge _539) begin
        if (_537)
            _4382 <= _567;
        else
            _4382 <= _297;
    end
    assign _4391 = _616 == _1059;
    assign _4389 = _565 & _570;
    assign _4392 = _4389 & _4391;
    assign _4396 = _4392 ? _597 : _4395;
    assign _4387 = _609 == _1059;
    assign _4385 = _565 & _580;
    assign _4388 = _4385 & _4387;
    assign _4397 = _4388 ? _577 : _4396;
    assign _298 = _4397;
    always @(posedge _539) begin
        if (_537)
            _4395 <= _567;
        else
            _4395 <= _298;
    end
    assign _4404 = _616 == _1072;
    assign _4402 = _565 & _570;
    assign _4405 = _4402 & _4404;
    assign _4409 = _4405 ? _597 : _4408;
    assign _4400 = _609 == _1072;
    assign _4398 = _565 & _580;
    assign _4401 = _4398 & _4400;
    assign _4410 = _4401 ? _577 : _4409;
    assign _299 = _4410;
    always @(posedge _539) begin
        if (_537)
            _4408 <= _567;
        else
            _4408 <= _299;
    end
    assign _4417 = _616 == _1085;
    assign _4415 = _565 & _570;
    assign _4418 = _4415 & _4417;
    assign _4422 = _4418 ? _597 : _4421;
    assign _4413 = _609 == _1085;
    assign _4411 = _565 & _580;
    assign _4414 = _4411 & _4413;
    assign _4423 = _4414 ? _577 : _4422;
    assign _300 = _4423;
    always @(posedge _539) begin
        if (_537)
            _4421 <= _567;
        else
            _4421 <= _300;
    end
    assign _4430 = _616 == _1098;
    assign _4428 = _565 & _570;
    assign _4431 = _4428 & _4430;
    assign _4435 = _4431 ? _597 : _4434;
    assign _4426 = _609 == _1098;
    assign _4424 = _565 & _580;
    assign _4427 = _4424 & _4426;
    assign _4436 = _4427 ? _577 : _4435;
    assign _301 = _4436;
    always @(posedge _539) begin
        if (_537)
            _4434 <= _567;
        else
            _4434 <= _301;
    end
    assign _4443 = _616 == _1111;
    assign _4441 = _565 & _570;
    assign _4444 = _4441 & _4443;
    assign _4448 = _4444 ? _597 : _4447;
    assign _4439 = _609 == _1111;
    assign _4437 = _565 & _580;
    assign _4440 = _4437 & _4439;
    assign _4449 = _4440 ? _577 : _4448;
    assign _302 = _4449;
    always @(posedge _539) begin
        if (_537)
            _4447 <= _567;
        else
            _4447 <= _302;
    end
    assign _4456 = _616 == _1124;
    assign _4454 = _565 & _570;
    assign _4457 = _4454 & _4456;
    assign _4461 = _4457 ? _597 : _4460;
    assign _4452 = _609 == _1124;
    assign _4450 = _565 & _580;
    assign _4453 = _4450 & _4452;
    assign _4462 = _4453 ? _577 : _4461;
    assign _303 = _4462;
    always @(posedge _539) begin
        if (_537)
            _4460 <= _567;
        else
            _4460 <= _303;
    end
    assign _4469 = _616 == _1137;
    assign _4467 = _565 & _570;
    assign _4470 = _4467 & _4469;
    assign _4474 = _4470 ? _597 : _4473;
    assign _4465 = _609 == _1137;
    assign _4463 = _565 & _580;
    assign _4466 = _4463 & _4465;
    assign _4475 = _4466 ? _577 : _4474;
    assign _304 = _4475;
    always @(posedge _539) begin
        if (_537)
            _4473 <= _567;
        else
            _4473 <= _304;
    end
    assign _4482 = _616 == _1150;
    assign _4480 = _565 & _570;
    assign _4483 = _4480 & _4482;
    assign _4487 = _4483 ? _597 : _4486;
    assign _4478 = _609 == _1150;
    assign _4476 = _565 & _580;
    assign _4479 = _4476 & _4478;
    assign _4488 = _4479 ? _577 : _4487;
    assign _305 = _4488;
    always @(posedge _539) begin
        if (_537)
            _4486 <= _567;
        else
            _4486 <= _305;
    end
    assign _4495 = _616 == _1163;
    assign _4493 = _565 & _570;
    assign _4496 = _4493 & _4495;
    assign _4500 = _4496 ? _597 : _4499;
    assign _4491 = _609 == _1163;
    assign _4489 = _565 & _580;
    assign _4492 = _4489 & _4491;
    assign _4501 = _4492 ? _577 : _4500;
    assign _306 = _4501;
    always @(posedge _539) begin
        if (_537)
            _4499 <= _567;
        else
            _4499 <= _306;
    end
    assign _4508 = _616 == _1176;
    assign _4506 = _565 & _570;
    assign _4509 = _4506 & _4508;
    assign _4513 = _4509 ? _597 : _4512;
    assign _4504 = _609 == _1176;
    assign _4502 = _565 & _580;
    assign _4505 = _4502 & _4504;
    assign _4514 = _4505 ? _577 : _4513;
    assign _307 = _4514;
    always @(posedge _539) begin
        if (_537)
            _4512 <= _567;
        else
            _4512 <= _307;
    end
    assign _4521 = _616 == _1189;
    assign _4519 = _565 & _570;
    assign _4522 = _4519 & _4521;
    assign _4526 = _4522 ? _597 : _4525;
    assign _4517 = _609 == _1189;
    assign _4515 = _565 & _580;
    assign _4518 = _4515 & _4517;
    assign _4527 = _4518 ? _577 : _4526;
    assign _308 = _4527;
    always @(posedge _539) begin
        if (_537)
            _4525 <= _567;
        else
            _4525 <= _308;
    end
    assign _4534 = _616 == _1202;
    assign _4532 = _565 & _570;
    assign _4535 = _4532 & _4534;
    assign _4539 = _4535 ? _597 : _4538;
    assign _4530 = _609 == _1202;
    assign _4528 = _565 & _580;
    assign _4531 = _4528 & _4530;
    assign _4540 = _4531 ? _577 : _4539;
    assign _309 = _4540;
    always @(posedge _539) begin
        if (_537)
            _4538 <= _567;
        else
            _4538 <= _309;
    end
    assign _4547 = _616 == _1215;
    assign _4545 = _565 & _570;
    assign _4548 = _4545 & _4547;
    assign _4552 = _4548 ? _597 : _4551;
    assign _4543 = _609 == _1215;
    assign _4541 = _565 & _580;
    assign _4544 = _4541 & _4543;
    assign _4553 = _4544 ? _577 : _4552;
    assign _310 = _4553;
    always @(posedge _539) begin
        if (_537)
            _4551 <= _567;
        else
            _4551 <= _310;
    end
    assign _4560 = _616 == _1228;
    assign _4558 = _565 & _570;
    assign _4561 = _4558 & _4560;
    assign _4565 = _4561 ? _597 : _4564;
    assign _4556 = _609 == _1228;
    assign _4554 = _565 & _580;
    assign _4557 = _4554 & _4556;
    assign _4566 = _4557 ? _577 : _4565;
    assign _311 = _4566;
    always @(posedge _539) begin
        if (_537)
            _4564 <= _567;
        else
            _4564 <= _311;
    end
    assign _4573 = _616 == _1241;
    assign _4571 = _565 & _570;
    assign _4574 = _4571 & _4573;
    assign _4578 = _4574 ? _597 : _4577;
    assign _4569 = _609 == _1241;
    assign _4567 = _565 & _580;
    assign _4570 = _4567 & _4569;
    assign _4579 = _4570 ? _577 : _4578;
    assign _312 = _4579;
    always @(posedge _539) begin
        if (_537)
            _4577 <= _567;
        else
            _4577 <= _312;
    end
    assign _4586 = _616 == _1254;
    assign _4584 = _565 & _570;
    assign _4587 = _4584 & _4586;
    assign _4591 = _4587 ? _597 : _4590;
    assign _4582 = _609 == _1254;
    assign _4580 = _565 & _580;
    assign _4583 = _4580 & _4582;
    assign _4592 = _4583 ? _577 : _4591;
    assign _313 = _4592;
    always @(posedge _539) begin
        if (_537)
            _4590 <= _567;
        else
            _4590 <= _313;
    end
    assign _4599 = _616 == _1267;
    assign _4597 = _565 & _570;
    assign _4600 = _4597 & _4599;
    assign _4604 = _4600 ? _597 : _4603;
    assign _4595 = _609 == _1267;
    assign _4593 = _565 & _580;
    assign _4596 = _4593 & _4595;
    assign _4605 = _4596 ? _577 : _4604;
    assign _314 = _4605;
    always @(posedge _539) begin
        if (_537)
            _4603 <= _567;
        else
            _4603 <= _314;
    end
    assign _4612 = _616 == _1280;
    assign _4610 = _565 & _570;
    assign _4613 = _4610 & _4612;
    assign _4617 = _4613 ? _597 : _4616;
    assign _4608 = _609 == _1280;
    assign _4606 = _565 & _580;
    assign _4609 = _4606 & _4608;
    assign _4618 = _4609 ? _577 : _4617;
    assign _315 = _4618;
    always @(posedge _539) begin
        if (_537)
            _4616 <= _567;
        else
            _4616 <= _315;
    end
    assign _4625 = _616 == _1293;
    assign _4623 = _565 & _570;
    assign _4626 = _4623 & _4625;
    assign _4630 = _4626 ? _597 : _4629;
    assign _4621 = _609 == _1293;
    assign _4619 = _565 & _580;
    assign _4622 = _4619 & _4621;
    assign _4631 = _4622 ? _577 : _4630;
    assign _316 = _4631;
    always @(posedge _539) begin
        if (_537)
            _4629 <= _567;
        else
            _4629 <= _316;
    end
    assign _4638 = _616 == _1306;
    assign _4636 = _565 & _570;
    assign _4639 = _4636 & _4638;
    assign _4643 = _4639 ? _597 : _4642;
    assign _4634 = _609 == _1306;
    assign _4632 = _565 & _580;
    assign _4635 = _4632 & _4634;
    assign _4644 = _4635 ? _577 : _4643;
    assign _317 = _4644;
    always @(posedge _539) begin
        if (_537)
            _4642 <= _567;
        else
            _4642 <= _317;
    end
    assign _4651 = _616 == _1319;
    assign _4649 = _565 & _570;
    assign _4652 = _4649 & _4651;
    assign _4656 = _4652 ? _597 : _4655;
    assign _4647 = _609 == _1319;
    assign _4645 = _565 & _580;
    assign _4648 = _4645 & _4647;
    assign _4657 = _4648 ? _577 : _4656;
    assign _318 = _4657;
    always @(posedge _539) begin
        if (_537)
            _4655 <= _567;
        else
            _4655 <= _318;
    end
    assign _4664 = _616 == _1332;
    assign _4662 = _565 & _570;
    assign _4665 = _4662 & _4664;
    assign _4669 = _4665 ? _597 : _4668;
    assign _4660 = _609 == _1332;
    assign _4658 = _565 & _580;
    assign _4661 = _4658 & _4660;
    assign _4670 = _4661 ? _577 : _4669;
    assign _319 = _4670;
    always @(posedge _539) begin
        if (_537)
            _4668 <= _567;
        else
            _4668 <= _319;
    end
    assign _4677 = _616 == _1345;
    assign _4675 = _565 & _570;
    assign _4678 = _4675 & _4677;
    assign _4682 = _4678 ? _597 : _4681;
    assign _4673 = _609 == _1345;
    assign _4671 = _565 & _580;
    assign _4674 = _4671 & _4673;
    assign _4683 = _4674 ? _577 : _4682;
    assign _320 = _4683;
    always @(posedge _539) begin
        if (_537)
            _4681 <= _567;
        else
            _4681 <= _320;
    end
    assign _4690 = _616 == _1358;
    assign _4688 = _565 & _570;
    assign _4691 = _4688 & _4690;
    assign _4695 = _4691 ? _597 : _4694;
    assign _4686 = _609 == _1358;
    assign _4684 = _565 & _580;
    assign _4687 = _4684 & _4686;
    assign _4696 = _4687 ? _577 : _4695;
    assign _321 = _4696;
    always @(posedge _539) begin
        if (_537)
            _4694 <= _567;
        else
            _4694 <= _321;
    end
    assign _4703 = _616 == _1371;
    assign _4701 = _565 & _570;
    assign _4704 = _4701 & _4703;
    assign _4708 = _4704 ? _597 : _4707;
    assign _4699 = _609 == _1371;
    assign _4697 = _565 & _580;
    assign _4700 = _4697 & _4699;
    assign _4709 = _4700 ? _577 : _4708;
    assign _322 = _4709;
    always @(posedge _539) begin
        if (_537)
            _4707 <= _567;
        else
            _4707 <= _322;
    end
    assign _4716 = _616 == _1384;
    assign _4714 = _565 & _570;
    assign _4717 = _4714 & _4716;
    assign _4721 = _4717 ? _597 : _4720;
    assign _4712 = _609 == _1384;
    assign _4710 = _565 & _580;
    assign _4713 = _4710 & _4712;
    assign _4722 = _4713 ? _577 : _4721;
    assign _323 = _4722;
    always @(posedge _539) begin
        if (_537)
            _4720 <= _567;
        else
            _4720 <= _323;
    end
    assign _4729 = _616 == _1397;
    assign _4727 = _565 & _570;
    assign _4730 = _4727 & _4729;
    assign _4734 = _4730 ? _597 : _4733;
    assign _4725 = _609 == _1397;
    assign _4723 = _565 & _580;
    assign _4726 = _4723 & _4725;
    assign _4735 = _4726 ? _577 : _4734;
    assign _324 = _4735;
    always @(posedge _539) begin
        if (_537)
            _4733 <= _567;
        else
            _4733 <= _324;
    end
    assign _4742 = _616 == _1410;
    assign _4740 = _565 & _570;
    assign _4743 = _4740 & _4742;
    assign _4747 = _4743 ? _597 : _4746;
    assign _4738 = _609 == _1410;
    assign _4736 = _565 & _580;
    assign _4739 = _4736 & _4738;
    assign _4748 = _4739 ? _577 : _4747;
    assign _325 = _4748;
    always @(posedge _539) begin
        if (_537)
            _4746 <= _567;
        else
            _4746 <= _325;
    end
    assign _4755 = _616 == _1423;
    assign _4753 = _565 & _570;
    assign _4756 = _4753 & _4755;
    assign _4760 = _4756 ? _597 : _4759;
    assign _4751 = _609 == _1423;
    assign _4749 = _565 & _580;
    assign _4752 = _4749 & _4751;
    assign _4761 = _4752 ? _577 : _4760;
    assign _326 = _4761;
    always @(posedge _539) begin
        if (_537)
            _4759 <= _567;
        else
            _4759 <= _326;
    end
    assign _4768 = _616 == _1436;
    assign _4766 = _565 & _570;
    assign _4769 = _4766 & _4768;
    assign _4773 = _4769 ? _597 : _4772;
    assign _4764 = _609 == _1436;
    assign _4762 = _565 & _580;
    assign _4765 = _4762 & _4764;
    assign _4774 = _4765 ? _577 : _4773;
    assign _327 = _4774;
    always @(posedge _539) begin
        if (_537)
            _4772 <= _567;
        else
            _4772 <= _327;
    end
    assign _4781 = _616 == _1449;
    assign _4779 = _565 & _570;
    assign _4782 = _4779 & _4781;
    assign _4786 = _4782 ? _597 : _4785;
    assign _4777 = _609 == _1449;
    assign _4775 = _565 & _580;
    assign _4778 = _4775 & _4777;
    assign _4787 = _4778 ? _577 : _4786;
    assign _328 = _4787;
    always @(posedge _539) begin
        if (_537)
            _4785 <= _567;
        else
            _4785 <= _328;
    end
    assign _4794 = _616 == _1462;
    assign _4792 = _565 & _570;
    assign _4795 = _4792 & _4794;
    assign _4799 = _4795 ? _597 : _4798;
    assign _4790 = _609 == _1462;
    assign _4788 = _565 & _580;
    assign _4791 = _4788 & _4790;
    assign _4800 = _4791 ? _577 : _4799;
    assign _329 = _4800;
    always @(posedge _539) begin
        if (_537)
            _4798 <= _567;
        else
            _4798 <= _329;
    end
    assign _4807 = _616 == _1475;
    assign _4805 = _565 & _570;
    assign _4808 = _4805 & _4807;
    assign _4812 = _4808 ? _597 : _4811;
    assign _4803 = _609 == _1475;
    assign _4801 = _565 & _580;
    assign _4804 = _4801 & _4803;
    assign _4813 = _4804 ? _577 : _4812;
    assign _330 = _4813;
    always @(posedge _539) begin
        if (_537)
            _4811 <= _567;
        else
            _4811 <= _330;
    end
    assign _4820 = _616 == _1488;
    assign _4818 = _565 & _570;
    assign _4821 = _4818 & _4820;
    assign _4825 = _4821 ? _597 : _4824;
    assign _4816 = _609 == _1488;
    assign _4814 = _565 & _580;
    assign _4817 = _4814 & _4816;
    assign _4826 = _4817 ? _577 : _4825;
    assign _331 = _4826;
    always @(posedge _539) begin
        if (_537)
            _4824 <= _567;
        else
            _4824 <= _331;
    end
    assign _4833 = _616 == _1501;
    assign _4831 = _565 & _570;
    assign _4834 = _4831 & _4833;
    assign _4838 = _4834 ? _597 : _4837;
    assign _4829 = _609 == _1501;
    assign _4827 = _565 & _580;
    assign _4830 = _4827 & _4829;
    assign _4839 = _4830 ? _577 : _4838;
    assign _332 = _4839;
    always @(posedge _539) begin
        if (_537)
            _4837 <= _567;
        else
            _4837 <= _332;
    end
    assign _4846 = _616 == _1514;
    assign _4844 = _565 & _570;
    assign _4847 = _4844 & _4846;
    assign _4851 = _4847 ? _597 : _4850;
    assign _4842 = _609 == _1514;
    assign _4840 = _565 & _580;
    assign _4843 = _4840 & _4842;
    assign _4852 = _4843 ? _577 : _4851;
    assign _333 = _4852;
    always @(posedge _539) begin
        if (_537)
            _4850 <= _567;
        else
            _4850 <= _333;
    end
    assign _4859 = _616 == _1527;
    assign _4857 = _565 & _570;
    assign _4860 = _4857 & _4859;
    assign _4864 = _4860 ? _597 : _4863;
    assign _4855 = _609 == _1527;
    assign _4853 = _565 & _580;
    assign _4856 = _4853 & _4855;
    assign _4865 = _4856 ? _577 : _4864;
    assign _334 = _4865;
    always @(posedge _539) begin
        if (_537)
            _4863 <= _567;
        else
            _4863 <= _334;
    end
    assign _4872 = _616 == _1540;
    assign _4870 = _565 & _570;
    assign _4873 = _4870 & _4872;
    assign _4877 = _4873 ? _597 : _4876;
    assign _4868 = _609 == _1540;
    assign _4866 = _565 & _580;
    assign _4869 = _4866 & _4868;
    assign _4878 = _4869 ? _577 : _4877;
    assign _335 = _4878;
    always @(posedge _539) begin
        if (_537)
            _4876 <= _567;
        else
            _4876 <= _335;
    end
    assign _4885 = _616 == _1553;
    assign _4883 = _565 & _570;
    assign _4886 = _4883 & _4885;
    assign _4890 = _4886 ? _597 : _4889;
    assign _4881 = _609 == _1553;
    assign _4879 = _565 & _580;
    assign _4882 = _4879 & _4881;
    assign _4891 = _4882 ? _577 : _4890;
    assign _336 = _4891;
    always @(posedge _539) begin
        if (_537)
            _4889 <= _567;
        else
            _4889 <= _336;
    end
    assign _4898 = _616 == _1566;
    assign _4896 = _565 & _570;
    assign _4899 = _4896 & _4898;
    assign _4903 = _4899 ? _597 : _4902;
    assign _4894 = _609 == _1566;
    assign _4892 = _565 & _580;
    assign _4895 = _4892 & _4894;
    assign _4904 = _4895 ? _577 : _4903;
    assign _337 = _4904;
    always @(posedge _539) begin
        if (_537)
            _4902 <= _567;
        else
            _4902 <= _337;
    end
    assign _4911 = _616 == _1579;
    assign _4909 = _565 & _570;
    assign _4912 = _4909 & _4911;
    assign _4916 = _4912 ? _597 : _4915;
    assign _4907 = _609 == _1579;
    assign _4905 = _565 & _580;
    assign _4908 = _4905 & _4907;
    assign _4917 = _4908 ? _577 : _4916;
    assign _338 = _4917;
    always @(posedge _539) begin
        if (_537)
            _4915 <= _567;
        else
            _4915 <= _338;
    end
    assign _4924 = _616 == _1592;
    assign _4922 = _565 & _570;
    assign _4925 = _4922 & _4924;
    assign _4929 = _4925 ? _597 : _4928;
    assign _4920 = _609 == _1592;
    assign _4918 = _565 & _580;
    assign _4921 = _4918 & _4920;
    assign _4930 = _4921 ? _577 : _4929;
    assign _339 = _4930;
    always @(posedge _539) begin
        if (_537)
            _4928 <= _567;
        else
            _4928 <= _339;
    end
    assign _4937 = _616 == _1605;
    assign _4935 = _565 & _570;
    assign _4938 = _4935 & _4937;
    assign _4942 = _4938 ? _597 : _4941;
    assign _4933 = _609 == _1605;
    assign _4931 = _565 & _580;
    assign _4934 = _4931 & _4933;
    assign _4943 = _4934 ? _577 : _4942;
    assign _340 = _4943;
    always @(posedge _539) begin
        if (_537)
            _4941 <= _567;
        else
            _4941 <= _340;
    end
    assign _4950 = _616 == _1618;
    assign _4948 = _565 & _570;
    assign _4951 = _4948 & _4950;
    assign _4955 = _4951 ? _597 : _4954;
    assign _4946 = _609 == _1618;
    assign _4944 = _565 & _580;
    assign _4947 = _4944 & _4946;
    assign _4956 = _4947 ? _577 : _4955;
    assign _341 = _4956;
    always @(posedge _539) begin
        if (_537)
            _4954 <= _567;
        else
            _4954 <= _341;
    end
    assign _4963 = _616 == _1631;
    assign _4961 = _565 & _570;
    assign _4964 = _4961 & _4963;
    assign _4968 = _4964 ? _597 : _4967;
    assign _4959 = _609 == _1631;
    assign _4957 = _565 & _580;
    assign _4960 = _4957 & _4959;
    assign _4969 = _4960 ? _577 : _4968;
    assign _342 = _4969;
    always @(posedge _539) begin
        if (_537)
            _4967 <= _567;
        else
            _4967 <= _342;
    end
    assign _4976 = _616 == _1644;
    assign _4974 = _565 & _570;
    assign _4977 = _4974 & _4976;
    assign _4981 = _4977 ? _597 : _4980;
    assign _4972 = _609 == _1644;
    assign _4970 = _565 & _580;
    assign _4973 = _4970 & _4972;
    assign _4982 = _4973 ? _577 : _4981;
    assign _343 = _4982;
    always @(posedge _539) begin
        if (_537)
            _4980 <= _567;
        else
            _4980 <= _343;
    end
    assign _4989 = _616 == _1657;
    assign _4987 = _565 & _570;
    assign _4990 = _4987 & _4989;
    assign _4994 = _4990 ? _597 : _4993;
    assign _4985 = _609 == _1657;
    assign _4983 = _565 & _580;
    assign _4986 = _4983 & _4985;
    assign _4995 = _4986 ? _577 : _4994;
    assign _344 = _4995;
    always @(posedge _539) begin
        if (_537)
            _4993 <= _567;
        else
            _4993 <= _344;
    end
    assign _5002 = _616 == _1670;
    assign _5000 = _565 & _570;
    assign _5003 = _5000 & _5002;
    assign _5007 = _5003 ? _597 : _5006;
    assign _4998 = _609 == _1670;
    assign _4996 = _565 & _580;
    assign _4999 = _4996 & _4998;
    assign _5008 = _4999 ? _577 : _5007;
    assign _345 = _5008;
    always @(posedge _539) begin
        if (_537)
            _5006 <= _567;
        else
            _5006 <= _345;
    end
    assign _5015 = _616 == _1683;
    assign _5013 = _565 & _570;
    assign _5016 = _5013 & _5015;
    assign _5020 = _5016 ? _597 : _5019;
    assign _5011 = _609 == _1683;
    assign _5009 = _565 & _580;
    assign _5012 = _5009 & _5011;
    assign _5021 = _5012 ? _577 : _5020;
    assign _346 = _5021;
    always @(posedge _539) begin
        if (_537)
            _5019 <= _567;
        else
            _5019 <= _346;
    end
    assign _5028 = _616 == _1696;
    assign _5026 = _565 & _570;
    assign _5029 = _5026 & _5028;
    assign _5033 = _5029 ? _597 : _5032;
    assign _5024 = _609 == _1696;
    assign _5022 = _565 & _580;
    assign _5025 = _5022 & _5024;
    assign _5034 = _5025 ? _577 : _5033;
    assign _347 = _5034;
    always @(posedge _539) begin
        if (_537)
            _5032 <= _567;
        else
            _5032 <= _347;
    end
    assign _5041 = _616 == _1709;
    assign _5039 = _565 & _570;
    assign _5042 = _5039 & _5041;
    assign _5046 = _5042 ? _597 : _5045;
    assign _5037 = _609 == _1709;
    assign _5035 = _565 & _580;
    assign _5038 = _5035 & _5037;
    assign _5047 = _5038 ? _577 : _5046;
    assign _348 = _5047;
    always @(posedge _539) begin
        if (_537)
            _5045 <= _567;
        else
            _5045 <= _348;
    end
    assign _5054 = _616 == _1722;
    assign _5052 = _565 & _570;
    assign _5055 = _5052 & _5054;
    assign _5059 = _5055 ? _597 : _5058;
    assign _5050 = _609 == _1722;
    assign _5048 = _565 & _580;
    assign _5051 = _5048 & _5050;
    assign _5060 = _5051 ? _577 : _5059;
    assign _349 = _5060;
    always @(posedge _539) begin
        if (_537)
            _5058 <= _567;
        else
            _5058 <= _349;
    end
    assign _5067 = _616 == _1735;
    assign _5065 = _565 & _570;
    assign _5068 = _5065 & _5067;
    assign _5072 = _5068 ? _597 : _5071;
    assign _5063 = _609 == _1735;
    assign _5061 = _565 & _580;
    assign _5064 = _5061 & _5063;
    assign _5073 = _5064 ? _577 : _5072;
    assign _350 = _5073;
    always @(posedge _539) begin
        if (_537)
            _5071 <= _567;
        else
            _5071 <= _350;
    end
    assign _5080 = _616 == _1748;
    assign _5078 = _565 & _570;
    assign _5081 = _5078 & _5080;
    assign _5085 = _5081 ? _597 : _5084;
    assign _5076 = _609 == _1748;
    assign _5074 = _565 & _580;
    assign _5077 = _5074 & _5076;
    assign _5086 = _5077 ? _577 : _5085;
    assign _351 = _5086;
    always @(posedge _539) begin
        if (_537)
            _5084 <= _567;
        else
            _5084 <= _351;
    end
    assign _5093 = _616 == _1761;
    assign _5091 = _565 & _570;
    assign _5094 = _5091 & _5093;
    assign _5098 = _5094 ? _597 : _5097;
    assign _5089 = _609 == _1761;
    assign _5087 = _565 & _580;
    assign _5090 = _5087 & _5089;
    assign _5099 = _5090 ? _577 : _5098;
    assign _352 = _5099;
    always @(posedge _539) begin
        if (_537)
            _5097 <= _567;
        else
            _5097 <= _352;
    end
    assign _5106 = _616 == _1774;
    assign _5104 = _565 & _570;
    assign _5107 = _5104 & _5106;
    assign _5111 = _5107 ? _597 : _5110;
    assign _5102 = _609 == _1774;
    assign _5100 = _565 & _580;
    assign _5103 = _5100 & _5102;
    assign _5112 = _5103 ? _577 : _5111;
    assign _353 = _5112;
    always @(posedge _539) begin
        if (_537)
            _5110 <= _567;
        else
            _5110 <= _353;
    end
    assign _5119 = _616 == _1787;
    assign _5117 = _565 & _570;
    assign _5120 = _5117 & _5119;
    assign _5124 = _5120 ? _597 : _5123;
    assign _5115 = _609 == _1787;
    assign _5113 = _565 & _580;
    assign _5116 = _5113 & _5115;
    assign _5125 = _5116 ? _577 : _5124;
    assign _354 = _5125;
    always @(posedge _539) begin
        if (_537)
            _5123 <= _567;
        else
            _5123 <= _354;
    end
    assign _5132 = _616 == _1800;
    assign _5130 = _565 & _570;
    assign _5133 = _5130 & _5132;
    assign _5137 = _5133 ? _597 : _5136;
    assign _5128 = _609 == _1800;
    assign _5126 = _565 & _580;
    assign _5129 = _5126 & _5128;
    assign _5138 = _5129 ? _577 : _5137;
    assign _355 = _5138;
    always @(posedge _539) begin
        if (_537)
            _5136 <= _567;
        else
            _5136 <= _355;
    end
    assign _5145 = _616 == _1813;
    assign _5143 = _565 & _570;
    assign _5146 = _5143 & _5145;
    assign _5150 = _5146 ? _597 : _5149;
    assign _5141 = _609 == _1813;
    assign _5139 = _565 & _580;
    assign _5142 = _5139 & _5141;
    assign _5151 = _5142 ? _577 : _5150;
    assign _356 = _5151;
    always @(posedge _539) begin
        if (_537)
            _5149 <= _567;
        else
            _5149 <= _356;
    end
    assign _5158 = _616 == _1826;
    assign _5156 = _565 & _570;
    assign _5159 = _5156 & _5158;
    assign _5163 = _5159 ? _597 : _5162;
    assign _5154 = _609 == _1826;
    assign _5152 = _565 & _580;
    assign _5155 = _5152 & _5154;
    assign _5164 = _5155 ? _577 : _5163;
    assign _357 = _5164;
    always @(posedge _539) begin
        if (_537)
            _5162 <= _567;
        else
            _5162 <= _357;
    end
    assign _5171 = _616 == _1839;
    assign _5169 = _565 & _570;
    assign _5172 = _5169 & _5171;
    assign _5176 = _5172 ? _597 : _5175;
    assign _5167 = _609 == _1839;
    assign _5165 = _565 & _580;
    assign _5168 = _5165 & _5167;
    assign _5177 = _5168 ? _577 : _5176;
    assign _358 = _5177;
    always @(posedge _539) begin
        if (_537)
            _5175 <= _567;
        else
            _5175 <= _358;
    end
    assign _5184 = _616 == _1852;
    assign _5182 = _565 & _570;
    assign _5185 = _5182 & _5184;
    assign _5189 = _5185 ? _597 : _5188;
    assign _5180 = _609 == _1852;
    assign _5178 = _565 & _580;
    assign _5181 = _5178 & _5180;
    assign _5190 = _5181 ? _577 : _5189;
    assign _359 = _5190;
    always @(posedge _539) begin
        if (_537)
            _5188 <= _567;
        else
            _5188 <= _359;
    end
    assign _5197 = _616 == _1865;
    assign _5195 = _565 & _570;
    assign _5198 = _5195 & _5197;
    assign _5202 = _5198 ? _597 : _5201;
    assign _5193 = _609 == _1865;
    assign _5191 = _565 & _580;
    assign _5194 = _5191 & _5193;
    assign _5203 = _5194 ? _577 : _5202;
    assign _360 = _5203;
    always @(posedge _539) begin
        if (_537)
            _5201 <= _567;
        else
            _5201 <= _360;
    end
    assign _5210 = _616 == _1878;
    assign _5208 = _565 & _570;
    assign _5211 = _5208 & _5210;
    assign _5215 = _5211 ? _597 : _5214;
    assign _5206 = _609 == _1878;
    assign _5204 = _565 & _580;
    assign _5207 = _5204 & _5206;
    assign _5216 = _5207 ? _577 : _5215;
    assign _361 = _5216;
    always @(posedge _539) begin
        if (_537)
            _5214 <= _567;
        else
            _5214 <= _361;
    end
    assign _5223 = _616 == _1891;
    assign _5221 = _565 & _570;
    assign _5224 = _5221 & _5223;
    assign _5228 = _5224 ? _597 : _5227;
    assign _5219 = _609 == _1891;
    assign _5217 = _565 & _580;
    assign _5220 = _5217 & _5219;
    assign _5229 = _5220 ? _577 : _5228;
    assign _362 = _5229;
    always @(posedge _539) begin
        if (_537)
            _5227 <= _567;
        else
            _5227 <= _362;
    end
    assign _5236 = _616 == _1904;
    assign _5234 = _565 & _570;
    assign _5237 = _5234 & _5236;
    assign _5241 = _5237 ? _597 : _5240;
    assign _5232 = _609 == _1904;
    assign _5230 = _565 & _580;
    assign _5233 = _5230 & _5232;
    assign _5242 = _5233 ? _577 : _5241;
    assign _363 = _5242;
    always @(posedge _539) begin
        if (_537)
            _5240 <= _567;
        else
            _5240 <= _363;
    end
    assign _5249 = _616 == _1917;
    assign _5247 = _565 & _570;
    assign _5250 = _5247 & _5249;
    assign _5254 = _5250 ? _597 : _5253;
    assign _5245 = _609 == _1917;
    assign _5243 = _565 & _580;
    assign _5246 = _5243 & _5245;
    assign _5255 = _5246 ? _577 : _5254;
    assign _364 = _5255;
    always @(posedge _539) begin
        if (_537)
            _5253 <= _567;
        else
            _5253 <= _364;
    end
    assign _5262 = _616 == _1930;
    assign _5260 = _565 & _570;
    assign _5263 = _5260 & _5262;
    assign _5267 = _5263 ? _597 : _5266;
    assign _5258 = _609 == _1930;
    assign _5256 = _565 & _580;
    assign _5259 = _5256 & _5258;
    assign _5268 = _5259 ? _577 : _5267;
    assign _365 = _5268;
    always @(posedge _539) begin
        if (_537)
            _5266 <= _567;
        else
            _5266 <= _365;
    end
    assign _5275 = _616 == _1943;
    assign _5273 = _565 & _570;
    assign _5276 = _5273 & _5275;
    assign _5280 = _5276 ? _597 : _5279;
    assign _5271 = _609 == _1943;
    assign _5269 = _565 & _580;
    assign _5272 = _5269 & _5271;
    assign _5281 = _5272 ? _577 : _5280;
    assign _366 = _5281;
    always @(posedge _539) begin
        if (_537)
            _5279 <= _567;
        else
            _5279 <= _366;
    end
    assign _5288 = _616 == _1956;
    assign _5286 = _565 & _570;
    assign _5289 = _5286 & _5288;
    assign _5293 = _5289 ? _597 : _5292;
    assign _5284 = _609 == _1956;
    assign _5282 = _565 & _580;
    assign _5285 = _5282 & _5284;
    assign _5294 = _5285 ? _577 : _5293;
    assign _367 = _5294;
    always @(posedge _539) begin
        if (_537)
            _5292 <= _567;
        else
            _5292 <= _367;
    end
    assign _5301 = _616 == _1969;
    assign _5299 = _565 & _570;
    assign _5302 = _5299 & _5301;
    assign _5306 = _5302 ? _597 : _5305;
    assign _5297 = _609 == _1969;
    assign _5295 = _565 & _580;
    assign _5298 = _5295 & _5297;
    assign _5307 = _5298 ? _577 : _5306;
    assign _368 = _5307;
    always @(posedge _539) begin
        if (_537)
            _5305 <= _567;
        else
            _5305 <= _368;
    end
    assign _5314 = _616 == _1982;
    assign _5312 = _565 & _570;
    assign _5315 = _5312 & _5314;
    assign _5319 = _5315 ? _597 : _5318;
    assign _5310 = _609 == _1982;
    assign _5308 = _565 & _580;
    assign _5311 = _5308 & _5310;
    assign _5320 = _5311 ? _577 : _5319;
    assign _369 = _5320;
    always @(posedge _539) begin
        if (_537)
            _5318 <= _567;
        else
            _5318 <= _369;
    end
    assign _5327 = _616 == _1995;
    assign _5325 = _565 & _570;
    assign _5328 = _5325 & _5327;
    assign _5332 = _5328 ? _597 : _5331;
    assign _5323 = _609 == _1995;
    assign _5321 = _565 & _580;
    assign _5324 = _5321 & _5323;
    assign _5333 = _5324 ? _577 : _5332;
    assign _370 = _5333;
    always @(posedge _539) begin
        if (_537)
            _5331 <= _567;
        else
            _5331 <= _370;
    end
    assign _5340 = _616 == _2008;
    assign _5338 = _565 & _570;
    assign _5341 = _5338 & _5340;
    assign _5345 = _5341 ? _597 : _5344;
    assign _5336 = _609 == _2008;
    assign _5334 = _565 & _580;
    assign _5337 = _5334 & _5336;
    assign _5346 = _5337 ? _577 : _5345;
    assign _371 = _5346;
    always @(posedge _539) begin
        if (_537)
            _5344 <= _567;
        else
            _5344 <= _371;
    end
    assign _5353 = _616 == _2021;
    assign _5351 = _565 & _570;
    assign _5354 = _5351 & _5353;
    assign _5358 = _5354 ? _597 : _5357;
    assign _5349 = _609 == _2021;
    assign _5347 = _565 & _580;
    assign _5350 = _5347 & _5349;
    assign _5359 = _5350 ? _577 : _5358;
    assign _372 = _5359;
    always @(posedge _539) begin
        if (_537)
            _5357 <= _567;
        else
            _5357 <= _372;
    end
    assign _5366 = _616 == _2034;
    assign _5364 = _565 & _570;
    assign _5367 = _5364 & _5366;
    assign _5371 = _5367 ? _597 : _5370;
    assign _5362 = _609 == _2034;
    assign _5360 = _565 & _580;
    assign _5363 = _5360 & _5362;
    assign _5372 = _5363 ? _577 : _5371;
    assign _373 = _5372;
    always @(posedge _539) begin
        if (_537)
            _5370 <= _567;
        else
            _5370 <= _373;
    end
    assign _5379 = _616 == _2047;
    assign _5377 = _565 & _570;
    assign _5380 = _5377 & _5379;
    assign _5384 = _5380 ? _597 : _5383;
    assign _5375 = _609 == _2047;
    assign _5373 = _565 & _580;
    assign _5376 = _5373 & _5375;
    assign _5385 = _5376 ? _577 : _5384;
    assign _374 = _5385;
    always @(posedge _539) begin
        if (_537)
            _5383 <= _567;
        else
            _5383 <= _374;
    end
    assign _5392 = _616 == _2060;
    assign _5390 = _565 & _570;
    assign _5393 = _5390 & _5392;
    assign _5397 = _5393 ? _597 : _5396;
    assign _5388 = _609 == _2060;
    assign _5386 = _565 & _580;
    assign _5389 = _5386 & _5388;
    assign _5398 = _5389 ? _577 : _5397;
    assign _375 = _5398;
    always @(posedge _539) begin
        if (_537)
            _5396 <= _567;
        else
            _5396 <= _375;
    end
    assign _5405 = _616 == _2073;
    assign _5403 = _565 & _570;
    assign _5406 = _5403 & _5405;
    assign _5410 = _5406 ? _597 : _5409;
    assign _5401 = _609 == _2073;
    assign _5399 = _565 & _580;
    assign _5402 = _5399 & _5401;
    assign _5411 = _5402 ? _577 : _5410;
    assign _376 = _5411;
    always @(posedge _539) begin
        if (_537)
            _5409 <= _567;
        else
            _5409 <= _376;
    end
    assign _5418 = _616 == _2086;
    assign _5416 = _565 & _570;
    assign _5419 = _5416 & _5418;
    assign _5423 = _5419 ? _597 : _5422;
    assign _5414 = _609 == _2086;
    assign _5412 = _565 & _580;
    assign _5415 = _5412 & _5414;
    assign _5424 = _5415 ? _577 : _5423;
    assign _377 = _5424;
    always @(posedge _539) begin
        if (_537)
            _5422 <= _567;
        else
            _5422 <= _377;
    end
    assign _5431 = _616 == _2099;
    assign _5429 = _565 & _570;
    assign _5432 = _5429 & _5431;
    assign _5436 = _5432 ? _597 : _5435;
    assign _5427 = _609 == _2099;
    assign _5425 = _565 & _580;
    assign _5428 = _5425 & _5427;
    assign _5437 = _5428 ? _577 : _5436;
    assign _378 = _5437;
    always @(posedge _539) begin
        if (_537)
            _5435 <= _567;
        else
            _5435 <= _378;
    end
    assign _5444 = _616 == _2112;
    assign _5442 = _565 & _570;
    assign _5445 = _5442 & _5444;
    assign _5449 = _5445 ? _597 : _5448;
    assign _5440 = _609 == _2112;
    assign _5438 = _565 & _580;
    assign _5441 = _5438 & _5440;
    assign _5450 = _5441 ? _577 : _5449;
    assign _379 = _5450;
    always @(posedge _539) begin
        if (_537)
            _5448 <= _567;
        else
            _5448 <= _379;
    end
    assign _5457 = _616 == _2125;
    assign _5455 = _565 & _570;
    assign _5458 = _5455 & _5457;
    assign _5462 = _5458 ? _597 : _5461;
    assign _5453 = _609 == _2125;
    assign _5451 = _565 & _580;
    assign _5454 = _5451 & _5453;
    assign _5463 = _5454 ? _577 : _5462;
    assign _380 = _5463;
    always @(posedge _539) begin
        if (_537)
            _5461 <= _567;
        else
            _5461 <= _380;
    end
    assign _5470 = _616 == _2138;
    assign _5468 = _565 & _570;
    assign _5471 = _5468 & _5470;
    assign _5475 = _5471 ? _597 : _5474;
    assign _5466 = _609 == _2138;
    assign _5464 = _565 & _580;
    assign _5467 = _5464 & _5466;
    assign _5476 = _5467 ? _577 : _5475;
    assign _381 = _5476;
    always @(posedge _539) begin
        if (_537)
            _5474 <= _567;
        else
            _5474 <= _381;
    end
    assign _5483 = _616 == _2151;
    assign _5481 = _565 & _570;
    assign _5484 = _5481 & _5483;
    assign _5488 = _5484 ? _597 : _5487;
    assign _5479 = _609 == _2151;
    assign _5477 = _565 & _580;
    assign _5480 = _5477 & _5479;
    assign _5489 = _5480 ? _577 : _5488;
    assign _382 = _5489;
    always @(posedge _539) begin
        if (_537)
            _5487 <= _567;
        else
            _5487 <= _382;
    end
    assign _5496 = _616 == _2164;
    assign _5494 = _565 & _570;
    assign _5497 = _5494 & _5496;
    assign _5501 = _5497 ? _597 : _5500;
    assign _5492 = _609 == _2164;
    assign _5490 = _565 & _580;
    assign _5493 = _5490 & _5492;
    assign _5502 = _5493 ? _577 : _5501;
    assign _383 = _5502;
    always @(posedge _539) begin
        if (_537)
            _5500 <= _567;
        else
            _5500 <= _383;
    end
    assign _5509 = _616 == _2177;
    assign _5507 = _565 & _570;
    assign _5510 = _5507 & _5509;
    assign _5514 = _5510 ? _597 : _5513;
    assign _5505 = _609 == _2177;
    assign _5503 = _565 & _580;
    assign _5506 = _5503 & _5505;
    assign _5515 = _5506 ? _577 : _5514;
    assign _384 = _5515;
    always @(posedge _539) begin
        if (_537)
            _5513 <= _567;
        else
            _5513 <= _384;
    end
    assign _5522 = _616 == _2190;
    assign _5520 = _565 & _570;
    assign _5523 = _5520 & _5522;
    assign _5527 = _5523 ? _597 : _5526;
    assign _5518 = _609 == _2190;
    assign _5516 = _565 & _580;
    assign _5519 = _5516 & _5518;
    assign _5528 = _5519 ? _577 : _5527;
    assign _385 = _5528;
    always @(posedge _539) begin
        if (_537)
            _5526 <= _567;
        else
            _5526 <= _385;
    end
    assign _5535 = _616 == _2203;
    assign _5533 = _565 & _570;
    assign _5536 = _5533 & _5535;
    assign _5540 = _5536 ? _597 : _5539;
    assign _5531 = _609 == _2203;
    assign _5529 = _565 & _580;
    assign _5532 = _5529 & _5531;
    assign _5541 = _5532 ? _577 : _5540;
    assign _386 = _5541;
    always @(posedge _539) begin
        if (_537)
            _5539 <= _567;
        else
            _5539 <= _386;
    end
    assign _5548 = _616 == _2216;
    assign _5546 = _565 & _570;
    assign _5549 = _5546 & _5548;
    assign _5553 = _5549 ? _597 : _5552;
    assign _5544 = _609 == _2216;
    assign _5542 = _565 & _580;
    assign _5545 = _5542 & _5544;
    assign _5554 = _5545 ? _577 : _5553;
    assign _387 = _5554;
    always @(posedge _539) begin
        if (_537)
            _5552 <= _567;
        else
            _5552 <= _387;
    end
    assign _5561 = _616 == _2229;
    assign _5559 = _565 & _570;
    assign _5562 = _5559 & _5561;
    assign _5566 = _5562 ? _597 : _5565;
    assign _5557 = _609 == _2229;
    assign _5555 = _565 & _580;
    assign _5558 = _5555 & _5557;
    assign _5567 = _5558 ? _577 : _5566;
    assign _388 = _5567;
    always @(posedge _539) begin
        if (_537)
            _5565 <= _567;
        else
            _5565 <= _388;
    end
    assign _5574 = _616 == _2242;
    assign _5572 = _565 & _570;
    assign _5575 = _5572 & _5574;
    assign _5579 = _5575 ? _597 : _5578;
    assign _5570 = _609 == _2242;
    assign _5568 = _565 & _580;
    assign _5571 = _5568 & _5570;
    assign _5580 = _5571 ? _577 : _5579;
    assign _389 = _5580;
    always @(posedge _539) begin
        if (_537)
            _5578 <= _567;
        else
            _5578 <= _389;
    end
    assign _5587 = _616 == _2255;
    assign _5585 = _565 & _570;
    assign _5588 = _5585 & _5587;
    assign _5592 = _5588 ? _597 : _5591;
    assign _5583 = _609 == _2255;
    assign _5581 = _565 & _580;
    assign _5584 = _5581 & _5583;
    assign _5593 = _5584 ? _577 : _5592;
    assign _390 = _5593;
    always @(posedge _539) begin
        if (_537)
            _5591 <= _567;
        else
            _5591 <= _390;
    end
    assign _5600 = _616 == _2268;
    assign _5598 = _565 & _570;
    assign _5601 = _5598 & _5600;
    assign _5605 = _5601 ? _597 : _5604;
    assign _5596 = _609 == _2268;
    assign _5594 = _565 & _580;
    assign _5597 = _5594 & _5596;
    assign _5606 = _5597 ? _577 : _5605;
    assign _391 = _5606;
    always @(posedge _539) begin
        if (_537)
            _5604 <= _567;
        else
            _5604 <= _391;
    end
    assign _5613 = _616 == _2281;
    assign _5611 = _565 & _570;
    assign _5614 = _5611 & _5613;
    assign _5618 = _5614 ? _597 : _5617;
    assign _5609 = _609 == _2281;
    assign _5607 = _565 & _580;
    assign _5610 = _5607 & _5609;
    assign _5619 = _5610 ? _577 : _5618;
    assign _392 = _5619;
    always @(posedge _539) begin
        if (_537)
            _5617 <= _567;
        else
            _5617 <= _392;
    end
    assign _5626 = _616 == _2294;
    assign _5624 = _565 & _570;
    assign _5627 = _5624 & _5626;
    assign _5631 = _5627 ? _597 : _5630;
    assign _5622 = _609 == _2294;
    assign _5620 = _565 & _580;
    assign _5623 = _5620 & _5622;
    assign _5632 = _5623 ? _577 : _5631;
    assign _393 = _5632;
    always @(posedge _539) begin
        if (_537)
            _5630 <= _567;
        else
            _5630 <= _393;
    end
    assign _5639 = _616 == _2307;
    assign _5637 = _565 & _570;
    assign _5640 = _5637 & _5639;
    assign _5644 = _5640 ? _597 : _5643;
    assign _5635 = _609 == _2307;
    assign _5633 = _565 & _580;
    assign _5636 = _5633 & _5635;
    assign _5645 = _5636 ? _577 : _5644;
    assign _394 = _5645;
    always @(posedge _539) begin
        if (_537)
            _5643 <= _567;
        else
            _5643 <= _394;
    end
    assign _5652 = _616 == _2320;
    assign _5650 = _565 & _570;
    assign _5653 = _5650 & _5652;
    assign _5657 = _5653 ? _597 : _5656;
    assign _5648 = _609 == _2320;
    assign _5646 = _565 & _580;
    assign _5649 = _5646 & _5648;
    assign _5658 = _5649 ? _577 : _5657;
    assign _395 = _5658;
    always @(posedge _539) begin
        if (_537)
            _5656 <= _567;
        else
            _5656 <= _395;
    end
    assign _5665 = _616 == _2333;
    assign _5663 = _565 & _570;
    assign _5666 = _5663 & _5665;
    assign _5670 = _5666 ? _597 : _5669;
    assign _5661 = _609 == _2333;
    assign _5659 = _565 & _580;
    assign _5662 = _5659 & _5661;
    assign _5671 = _5662 ? _577 : _5670;
    assign _396 = _5671;
    always @(posedge _539) begin
        if (_537)
            _5669 <= _567;
        else
            _5669 <= _396;
    end
    assign _5678 = _616 == _2346;
    assign _5676 = _565 & _570;
    assign _5679 = _5676 & _5678;
    assign _5683 = _5679 ? _597 : _5682;
    assign _5674 = _609 == _2346;
    assign _5672 = _565 & _580;
    assign _5675 = _5672 & _5674;
    assign _5684 = _5675 ? _577 : _5683;
    assign _397 = _5684;
    always @(posedge _539) begin
        if (_537)
            _5682 <= _567;
        else
            _5682 <= _397;
    end
    assign _5691 = _616 == _2359;
    assign _5689 = _565 & _570;
    assign _5692 = _5689 & _5691;
    assign _5696 = _5692 ? _597 : _5695;
    assign _5687 = _609 == _2359;
    assign _5685 = _565 & _580;
    assign _5688 = _5685 & _5687;
    assign _5697 = _5688 ? _577 : _5696;
    assign _398 = _5697;
    always @(posedge _539) begin
        if (_537)
            _5695 <= _567;
        else
            _5695 <= _398;
    end
    assign _5704 = _616 == _2372;
    assign _5702 = _565 & _570;
    assign _5705 = _5702 & _5704;
    assign _5709 = _5705 ? _597 : _5708;
    assign _5700 = _609 == _2372;
    assign _5698 = _565 & _580;
    assign _5701 = _5698 & _5700;
    assign _5710 = _5701 ? _577 : _5709;
    assign _399 = _5710;
    always @(posedge _539) begin
        if (_537)
            _5708 <= _567;
        else
            _5708 <= _399;
    end
    assign _5717 = _616 == _2385;
    assign _5715 = _565 & _570;
    assign _5718 = _5715 & _5717;
    assign _5722 = _5718 ? _597 : _5721;
    assign _5713 = _609 == _2385;
    assign _5711 = _565 & _580;
    assign _5714 = _5711 & _5713;
    assign _5723 = _5714 ? _577 : _5722;
    assign _400 = _5723;
    always @(posedge _539) begin
        if (_537)
            _5721 <= _567;
        else
            _5721 <= _400;
    end
    assign _5730 = _616 == _2398;
    assign _5728 = _565 & _570;
    assign _5731 = _5728 & _5730;
    assign _5735 = _5731 ? _597 : _5734;
    assign _5726 = _609 == _2398;
    assign _5724 = _565 & _580;
    assign _5727 = _5724 & _5726;
    assign _5736 = _5727 ? _577 : _5735;
    assign _401 = _5736;
    always @(posedge _539) begin
        if (_537)
            _5734 <= _567;
        else
            _5734 <= _401;
    end
    assign _5743 = _616 == _2411;
    assign _5741 = _565 & _570;
    assign _5744 = _5741 & _5743;
    assign _5748 = _5744 ? _597 : _5747;
    assign _5739 = _609 == _2411;
    assign _5737 = _565 & _580;
    assign _5740 = _5737 & _5739;
    assign _5749 = _5740 ? _577 : _5748;
    assign _402 = _5749;
    always @(posedge _539) begin
        if (_537)
            _5747 <= _567;
        else
            _5747 <= _402;
    end
    assign _5756 = _616 == _2424;
    assign _5754 = _565 & _570;
    assign _5757 = _5754 & _5756;
    assign _5761 = _5757 ? _597 : _5760;
    assign _5752 = _609 == _2424;
    assign _5750 = _565 & _580;
    assign _5753 = _5750 & _5752;
    assign _5762 = _5753 ? _577 : _5761;
    assign _403 = _5762;
    always @(posedge _539) begin
        if (_537)
            _5760 <= _567;
        else
            _5760 <= _403;
    end
    assign _5769 = _616 == _2437;
    assign _5767 = _565 & _570;
    assign _5770 = _5767 & _5769;
    assign _5774 = _5770 ? _597 : _5773;
    assign _5765 = _609 == _2437;
    assign _5763 = _565 & _580;
    assign _5766 = _5763 & _5765;
    assign _5775 = _5766 ? _577 : _5774;
    assign _404 = _5775;
    always @(posedge _539) begin
        if (_537)
            _5773 <= _567;
        else
            _5773 <= _404;
    end
    assign _5782 = _616 == _2450;
    assign _5780 = _565 & _570;
    assign _5783 = _5780 & _5782;
    assign _5787 = _5783 ? _597 : _5786;
    assign _5778 = _609 == _2450;
    assign _5776 = _565 & _580;
    assign _5779 = _5776 & _5778;
    assign _5788 = _5779 ? _577 : _5787;
    assign _405 = _5788;
    always @(posedge _539) begin
        if (_537)
            _5786 <= _567;
        else
            _5786 <= _405;
    end
    assign _5795 = _616 == _2463;
    assign _5793 = _565 & _570;
    assign _5796 = _5793 & _5795;
    assign _5800 = _5796 ? _597 : _5799;
    assign _5791 = _609 == _2463;
    assign _5789 = _565 & _580;
    assign _5792 = _5789 & _5791;
    assign _5801 = _5792 ? _577 : _5800;
    assign _406 = _5801;
    always @(posedge _539) begin
        if (_537)
            _5799 <= _567;
        else
            _5799 <= _406;
    end
    assign _5808 = _616 == _2476;
    assign _5806 = _565 & _570;
    assign _5809 = _5806 & _5808;
    assign _5813 = _5809 ? _597 : _5812;
    assign _5804 = _609 == _2476;
    assign _5802 = _565 & _580;
    assign _5805 = _5802 & _5804;
    assign _5814 = _5805 ? _577 : _5813;
    assign _407 = _5814;
    always @(posedge _539) begin
        if (_537)
            _5812 <= _567;
        else
            _5812 <= _407;
    end
    assign _5821 = _616 == _2489;
    assign _5819 = _565 & _570;
    assign _5822 = _5819 & _5821;
    assign _5826 = _5822 ? _597 : _5825;
    assign _5817 = _609 == _2489;
    assign _5815 = _565 & _580;
    assign _5818 = _5815 & _5817;
    assign _5827 = _5818 ? _577 : _5826;
    assign _408 = _5827;
    always @(posedge _539) begin
        if (_537)
            _5825 <= _567;
        else
            _5825 <= _408;
    end
    assign _5834 = _616 == _2502;
    assign _5832 = _565 & _570;
    assign _5835 = _5832 & _5834;
    assign _5839 = _5835 ? _597 : _5838;
    assign _5830 = _609 == _2502;
    assign _5828 = _565 & _580;
    assign _5831 = _5828 & _5830;
    assign _5840 = _5831 ? _577 : _5839;
    assign _409 = _5840;
    always @(posedge _539) begin
        if (_537)
            _5838 <= _567;
        else
            _5838 <= _409;
    end
    assign _5847 = _616 == _2515;
    assign _5845 = _565 & _570;
    assign _5848 = _5845 & _5847;
    assign _5852 = _5848 ? _597 : _5851;
    assign _5843 = _609 == _2515;
    assign _5841 = _565 & _580;
    assign _5844 = _5841 & _5843;
    assign _5853 = _5844 ? _577 : _5852;
    assign _410 = _5853;
    always @(posedge _539) begin
        if (_537)
            _5851 <= _567;
        else
            _5851 <= _410;
    end
    assign _5860 = _616 == _2528;
    assign _5858 = _565 & _570;
    assign _5861 = _5858 & _5860;
    assign _5865 = _5861 ? _597 : _5864;
    assign _5856 = _609 == _2528;
    assign _5854 = _565 & _580;
    assign _5857 = _5854 & _5856;
    assign _5866 = _5857 ? _577 : _5865;
    assign _411 = _5866;
    always @(posedge _539) begin
        if (_537)
            _5864 <= _567;
        else
            _5864 <= _411;
    end
    assign _5873 = _616 == _2541;
    assign _5871 = _565 & _570;
    assign _5874 = _5871 & _5873;
    assign _5878 = _5874 ? _597 : _5877;
    assign _5869 = _609 == _2541;
    assign _5867 = _565 & _580;
    assign _5870 = _5867 & _5869;
    assign _5879 = _5870 ? _577 : _5878;
    assign _412 = _5879;
    always @(posedge _539) begin
        if (_537)
            _5877 <= _567;
        else
            _5877 <= _412;
    end
    assign _5886 = _616 == _2554;
    assign _5884 = _565 & _570;
    assign _5887 = _5884 & _5886;
    assign _5891 = _5887 ? _597 : _5890;
    assign _5882 = _609 == _2554;
    assign _5880 = _565 & _580;
    assign _5883 = _5880 & _5882;
    assign _5892 = _5883 ? _577 : _5891;
    assign _413 = _5892;
    always @(posedge _539) begin
        if (_537)
            _5890 <= _567;
        else
            _5890 <= _413;
    end
    assign _5899 = _616 == _2567;
    assign _5897 = _565 & _570;
    assign _5900 = _5897 & _5899;
    assign _5904 = _5900 ? _597 : _5903;
    assign _5895 = _609 == _2567;
    assign _5893 = _565 & _580;
    assign _5896 = _5893 & _5895;
    assign _5905 = _5896 ? _577 : _5904;
    assign _414 = _5905;
    always @(posedge _539) begin
        if (_537)
            _5903 <= _567;
        else
            _5903 <= _414;
    end
    assign _5912 = _616 == _2580;
    assign _5910 = _565 & _570;
    assign _5913 = _5910 & _5912;
    assign _5917 = _5913 ? _597 : _5916;
    assign _5908 = _609 == _2580;
    assign _5906 = _565 & _580;
    assign _5909 = _5906 & _5908;
    assign _5918 = _5909 ? _577 : _5917;
    assign _415 = _5918;
    always @(posedge _539) begin
        if (_537)
            _5916 <= _567;
        else
            _5916 <= _415;
    end
    assign _5925 = _616 == _2593;
    assign _5923 = _565 & _570;
    assign _5926 = _5923 & _5925;
    assign _5930 = _5926 ? _597 : _5929;
    assign _5921 = _609 == _2593;
    assign _5919 = _565 & _580;
    assign _5922 = _5919 & _5921;
    assign _5931 = _5922 ? _577 : _5930;
    assign _416 = _5931;
    always @(posedge _539) begin
        if (_537)
            _5929 <= _567;
        else
            _5929 <= _416;
    end
    assign _5938 = _616 == _2606;
    assign _5936 = _565 & _570;
    assign _5939 = _5936 & _5938;
    assign _5943 = _5939 ? _597 : _5942;
    assign _5934 = _609 == _2606;
    assign _5932 = _565 & _580;
    assign _5935 = _5932 & _5934;
    assign _5944 = _5935 ? _577 : _5943;
    assign _417 = _5944;
    always @(posedge _539) begin
        if (_537)
            _5942 <= _567;
        else
            _5942 <= _417;
    end
    assign _5951 = _616 == _2619;
    assign _5949 = _565 & _570;
    assign _5952 = _5949 & _5951;
    assign _5956 = _5952 ? _597 : _5955;
    assign _5947 = _609 == _2619;
    assign _5945 = _565 & _580;
    assign _5948 = _5945 & _5947;
    assign _5957 = _5948 ? _577 : _5956;
    assign _418 = _5957;
    always @(posedge _539) begin
        if (_537)
            _5955 <= _567;
        else
            _5955 <= _418;
    end
    assign _5964 = _616 == _2632;
    assign _5962 = _565 & _570;
    assign _5965 = _5962 & _5964;
    assign _5969 = _5965 ? _597 : _5968;
    assign _5960 = _609 == _2632;
    assign _5958 = _565 & _580;
    assign _5961 = _5958 & _5960;
    assign _5970 = _5961 ? _577 : _5969;
    assign _419 = _5970;
    always @(posedge _539) begin
        if (_537)
            _5968 <= _567;
        else
            _5968 <= _419;
    end
    assign _5977 = _616 == _2645;
    assign _5975 = _565 & _570;
    assign _5978 = _5975 & _5977;
    assign _5982 = _5978 ? _597 : _5981;
    assign _5973 = _609 == _2645;
    assign _5971 = _565 & _580;
    assign _5974 = _5971 & _5973;
    assign _5983 = _5974 ? _577 : _5982;
    assign _420 = _5983;
    always @(posedge _539) begin
        if (_537)
            _5981 <= _567;
        else
            _5981 <= _420;
    end
    assign _5990 = _616 == _2658;
    assign _5988 = _565 & _570;
    assign _5991 = _5988 & _5990;
    assign _5995 = _5991 ? _597 : _5994;
    assign _5986 = _609 == _2658;
    assign _5984 = _565 & _580;
    assign _5987 = _5984 & _5986;
    assign _5996 = _5987 ? _577 : _5995;
    assign _421 = _5996;
    always @(posedge _539) begin
        if (_537)
            _5994 <= _567;
        else
            _5994 <= _421;
    end
    assign _6003 = _616 == _2671;
    assign _6001 = _565 & _570;
    assign _6004 = _6001 & _6003;
    assign _6008 = _6004 ? _597 : _6007;
    assign _5999 = _609 == _2671;
    assign _5997 = _565 & _580;
    assign _6000 = _5997 & _5999;
    assign _6009 = _6000 ? _577 : _6008;
    assign _422 = _6009;
    always @(posedge _539) begin
        if (_537)
            _6007 <= _567;
        else
            _6007 <= _422;
    end
    assign _6016 = _616 == _2684;
    assign _6014 = _565 & _570;
    assign _6017 = _6014 & _6016;
    assign _6021 = _6017 ? _597 : _6020;
    assign _6012 = _609 == _2684;
    assign _6010 = _565 & _580;
    assign _6013 = _6010 & _6012;
    assign _6022 = _6013 ? _577 : _6021;
    assign _423 = _6022;
    always @(posedge _539) begin
        if (_537)
            _6020 <= _567;
        else
            _6020 <= _423;
    end
    assign _6029 = _616 == _2697;
    assign _6027 = _565 & _570;
    assign _6030 = _6027 & _6029;
    assign _6034 = _6030 ? _597 : _6033;
    assign _6025 = _609 == _2697;
    assign _6023 = _565 & _580;
    assign _6026 = _6023 & _6025;
    assign _6035 = _6026 ? _577 : _6034;
    assign _424 = _6035;
    always @(posedge _539) begin
        if (_537)
            _6033 <= _567;
        else
            _6033 <= _424;
    end
    assign _6042 = _616 == _2710;
    assign _6040 = _565 & _570;
    assign _6043 = _6040 & _6042;
    assign _6047 = _6043 ? _597 : _6046;
    assign _6038 = _609 == _2710;
    assign _6036 = _565 & _580;
    assign _6039 = _6036 & _6038;
    assign _6048 = _6039 ? _577 : _6047;
    assign _425 = _6048;
    always @(posedge _539) begin
        if (_537)
            _6046 <= _567;
        else
            _6046 <= _425;
    end
    assign _6055 = _616 == _2723;
    assign _6053 = _565 & _570;
    assign _6056 = _6053 & _6055;
    assign _6060 = _6056 ? _597 : _6059;
    assign _6051 = _609 == _2723;
    assign _6049 = _565 & _580;
    assign _6052 = _6049 & _6051;
    assign _6061 = _6052 ? _577 : _6060;
    assign _426 = _6061;
    always @(posedge _539) begin
        if (_537)
            _6059 <= _567;
        else
            _6059 <= _426;
    end
    assign _6068 = _616 == _2736;
    assign _6066 = _565 & _570;
    assign _6069 = _6066 & _6068;
    assign _6073 = _6069 ? _597 : _6072;
    assign _6064 = _609 == _2736;
    assign _6062 = _565 & _580;
    assign _6065 = _6062 & _6064;
    assign _6074 = _6065 ? _577 : _6073;
    assign _427 = _6074;
    always @(posedge _539) begin
        if (_537)
            _6072 <= _567;
        else
            _6072 <= _427;
    end
    assign _6081 = _616 == _2749;
    assign _6079 = _565 & _570;
    assign _6082 = _6079 & _6081;
    assign _6086 = _6082 ? _597 : _6085;
    assign _6077 = _609 == _2749;
    assign _6075 = _565 & _580;
    assign _6078 = _6075 & _6077;
    assign _6087 = _6078 ? _577 : _6086;
    assign _428 = _6087;
    always @(posedge _539) begin
        if (_537)
            _6085 <= _567;
        else
            _6085 <= _428;
    end
    assign _6094 = _616 == _2762;
    assign _6092 = _565 & _570;
    assign _6095 = _6092 & _6094;
    assign _6099 = _6095 ? _597 : _6098;
    assign _6090 = _609 == _2762;
    assign _6088 = _565 & _580;
    assign _6091 = _6088 & _6090;
    assign _6100 = _6091 ? _577 : _6099;
    assign _429 = _6100;
    always @(posedge _539) begin
        if (_537)
            _6098 <= _567;
        else
            _6098 <= _429;
    end
    assign _6107 = _616 == _2775;
    assign _6105 = _565 & _570;
    assign _6108 = _6105 & _6107;
    assign _6112 = _6108 ? _597 : _6111;
    assign _6103 = _609 == _2775;
    assign _6101 = _565 & _580;
    assign _6104 = _6101 & _6103;
    assign _6113 = _6104 ? _577 : _6112;
    assign _430 = _6113;
    always @(posedge _539) begin
        if (_537)
            _6111 <= _567;
        else
            _6111 <= _430;
    end
    assign _6120 = _616 == _2788;
    assign _6118 = _565 & _570;
    assign _6121 = _6118 & _6120;
    assign _6125 = _6121 ? _597 : _6124;
    assign _6116 = _609 == _2788;
    assign _6114 = _565 & _580;
    assign _6117 = _6114 & _6116;
    assign _6126 = _6117 ? _577 : _6125;
    assign _431 = _6126;
    always @(posedge _539) begin
        if (_537)
            _6124 <= _567;
        else
            _6124 <= _431;
    end
    assign _6133 = _616 == _2801;
    assign _6131 = _565 & _570;
    assign _6134 = _6131 & _6133;
    assign _6138 = _6134 ? _597 : _6137;
    assign _6129 = _609 == _2801;
    assign _6127 = _565 & _580;
    assign _6130 = _6127 & _6129;
    assign _6139 = _6130 ? _577 : _6138;
    assign _432 = _6139;
    always @(posedge _539) begin
        if (_537)
            _6137 <= _567;
        else
            _6137 <= _432;
    end
    assign _6146 = _616 == _2814;
    assign _6144 = _565 & _570;
    assign _6147 = _6144 & _6146;
    assign _6151 = _6147 ? _597 : _6150;
    assign _6142 = _609 == _2814;
    assign _6140 = _565 & _580;
    assign _6143 = _6140 & _6142;
    assign _6152 = _6143 ? _577 : _6151;
    assign _433 = _6152;
    always @(posedge _539) begin
        if (_537)
            _6150 <= _567;
        else
            _6150 <= _433;
    end
    assign _6159 = _616 == _2827;
    assign _6157 = _565 & _570;
    assign _6160 = _6157 & _6159;
    assign _6164 = _6160 ? _597 : _6163;
    assign _6155 = _609 == _2827;
    assign _6153 = _565 & _580;
    assign _6156 = _6153 & _6155;
    assign _6165 = _6156 ? _577 : _6164;
    assign _434 = _6165;
    always @(posedge _539) begin
        if (_537)
            _6163 <= _567;
        else
            _6163 <= _434;
    end
    assign _6172 = _616 == _2840;
    assign _6170 = _565 & _570;
    assign _6173 = _6170 & _6172;
    assign _6177 = _6173 ? _597 : _6176;
    assign _6168 = _609 == _2840;
    assign _6166 = _565 & _580;
    assign _6169 = _6166 & _6168;
    assign _6178 = _6169 ? _577 : _6177;
    assign _435 = _6178;
    always @(posedge _539) begin
        if (_537)
            _6176 <= _567;
        else
            _6176 <= _435;
    end
    assign _6185 = _616 == _2853;
    assign _6183 = _565 & _570;
    assign _6186 = _6183 & _6185;
    assign _6190 = _6186 ? _597 : _6189;
    assign _6181 = _609 == _2853;
    assign _6179 = _565 & _580;
    assign _6182 = _6179 & _6181;
    assign _6191 = _6182 ? _577 : _6190;
    assign _436 = _6191;
    always @(posedge _539) begin
        if (_537)
            _6189 <= _567;
        else
            _6189 <= _436;
    end
    assign _6198 = _616 == _2866;
    assign _6196 = _565 & _570;
    assign _6199 = _6196 & _6198;
    assign _6203 = _6199 ? _597 : _6202;
    assign _6194 = _609 == _2866;
    assign _6192 = _565 & _580;
    assign _6195 = _6192 & _6194;
    assign _6204 = _6195 ? _577 : _6203;
    assign _437 = _6204;
    always @(posedge _539) begin
        if (_537)
            _6202 <= _567;
        else
            _6202 <= _437;
    end
    assign _6211 = _616 == _2879;
    assign _6209 = _565 & _570;
    assign _6212 = _6209 & _6211;
    assign _6216 = _6212 ? _597 : _6215;
    assign _6207 = _609 == _2879;
    assign _6205 = _565 & _580;
    assign _6208 = _6205 & _6207;
    assign _6217 = _6208 ? _577 : _6216;
    assign _438 = _6217;
    always @(posedge _539) begin
        if (_537)
            _6215 <= _567;
        else
            _6215 <= _438;
    end
    assign _6224 = _616 == _2892;
    assign _6222 = _565 & _570;
    assign _6225 = _6222 & _6224;
    assign _6229 = _6225 ? _597 : _6228;
    assign _6220 = _609 == _2892;
    assign _6218 = _565 & _580;
    assign _6221 = _6218 & _6220;
    assign _6230 = _6221 ? _577 : _6229;
    assign _439 = _6230;
    always @(posedge _539) begin
        if (_537)
            _6228 <= _567;
        else
            _6228 <= _439;
    end
    assign _6237 = _616 == _2905;
    assign _6235 = _565 & _570;
    assign _6238 = _6235 & _6237;
    assign _6242 = _6238 ? _597 : _6241;
    assign _6233 = _609 == _2905;
    assign _6231 = _565 & _580;
    assign _6234 = _6231 & _6233;
    assign _6243 = _6234 ? _577 : _6242;
    assign _440 = _6243;
    always @(posedge _539) begin
        if (_537)
            _6241 <= _567;
        else
            _6241 <= _440;
    end
    assign _6250 = _616 == _2918;
    assign _6248 = _565 & _570;
    assign _6251 = _6248 & _6250;
    assign _6255 = _6251 ? _597 : _6254;
    assign _6246 = _609 == _2918;
    assign _6244 = _565 & _580;
    assign _6247 = _6244 & _6246;
    assign _6256 = _6247 ? _577 : _6255;
    assign _441 = _6256;
    always @(posedge _539) begin
        if (_537)
            _6254 <= _567;
        else
            _6254 <= _441;
    end
    assign _6263 = _616 == _2931;
    assign _6261 = _565 & _570;
    assign _6264 = _6261 & _6263;
    assign _6268 = _6264 ? _597 : _6267;
    assign _6259 = _609 == _2931;
    assign _6257 = _565 & _580;
    assign _6260 = _6257 & _6259;
    assign _6269 = _6260 ? _577 : _6268;
    assign _442 = _6269;
    always @(posedge _539) begin
        if (_537)
            _6267 <= _567;
        else
            _6267 <= _442;
    end
    assign _6276 = _616 == _2944;
    assign _6274 = _565 & _570;
    assign _6277 = _6274 & _6276;
    assign _6281 = _6277 ? _597 : _6280;
    assign _6272 = _609 == _2944;
    assign _6270 = _565 & _580;
    assign _6273 = _6270 & _6272;
    assign _6282 = _6273 ? _577 : _6281;
    assign _443 = _6282;
    always @(posedge _539) begin
        if (_537)
            _6280 <= _567;
        else
            _6280 <= _443;
    end
    assign _6289 = _616 == _2957;
    assign _6287 = _565 & _570;
    assign _6290 = _6287 & _6289;
    assign _6294 = _6290 ? _597 : _6293;
    assign _6285 = _609 == _2957;
    assign _6283 = _565 & _580;
    assign _6286 = _6283 & _6285;
    assign _6295 = _6286 ? _577 : _6294;
    assign _444 = _6295;
    always @(posedge _539) begin
        if (_537)
            _6293 <= _567;
        else
            _6293 <= _444;
    end
    assign _6302 = _616 == _2970;
    assign _6300 = _565 & _570;
    assign _6303 = _6300 & _6302;
    assign _6307 = _6303 ? _597 : _6306;
    assign _6298 = _609 == _2970;
    assign _6296 = _565 & _580;
    assign _6299 = _6296 & _6298;
    assign _6308 = _6299 ? _577 : _6307;
    assign _445 = _6308;
    always @(posedge _539) begin
        if (_537)
            _6306 <= _567;
        else
            _6306 <= _445;
    end
    assign _6315 = _616 == _2983;
    assign _6313 = _565 & _570;
    assign _6316 = _6313 & _6315;
    assign _6320 = _6316 ? _597 : _6319;
    assign _6311 = _609 == _2983;
    assign _6309 = _565 & _580;
    assign _6312 = _6309 & _6311;
    assign _6321 = _6312 ? _577 : _6320;
    assign _446 = _6321;
    always @(posedge _539) begin
        if (_537)
            _6319 <= _567;
        else
            _6319 <= _446;
    end
    assign _6328 = _616 == _2996;
    assign _6326 = _565 & _570;
    assign _6329 = _6326 & _6328;
    assign _6333 = _6329 ? _597 : _6332;
    assign _6324 = _609 == _2996;
    assign _6322 = _565 & _580;
    assign _6325 = _6322 & _6324;
    assign _6334 = _6325 ? _577 : _6333;
    assign _447 = _6334;
    always @(posedge _539) begin
        if (_537)
            _6332 <= _567;
        else
            _6332 <= _447;
    end
    assign _6341 = _616 == _3009;
    assign _6339 = _565 & _570;
    assign _6342 = _6339 & _6341;
    assign _6346 = _6342 ? _597 : _6345;
    assign _6337 = _609 == _3009;
    assign _6335 = _565 & _580;
    assign _6338 = _6335 & _6337;
    assign _6347 = _6338 ? _577 : _6346;
    assign _448 = _6347;
    always @(posedge _539) begin
        if (_537)
            _6345 <= _567;
        else
            _6345 <= _448;
    end
    assign _6354 = _616 == _3022;
    assign _6352 = _565 & _570;
    assign _6355 = _6352 & _6354;
    assign _6359 = _6355 ? _597 : _6358;
    assign _6350 = _609 == _3022;
    assign _6348 = _565 & _580;
    assign _6351 = _6348 & _6350;
    assign _6360 = _6351 ? _577 : _6359;
    assign _449 = _6360;
    always @(posedge _539) begin
        if (_537)
            _6358 <= _567;
        else
            _6358 <= _449;
    end
    assign _6367 = _616 == _3035;
    assign _6365 = _565 & _570;
    assign _6368 = _6365 & _6367;
    assign _6372 = _6368 ? _597 : _6371;
    assign _6363 = _609 == _3035;
    assign _6361 = _565 & _580;
    assign _6364 = _6361 & _6363;
    assign _6373 = _6364 ? _577 : _6372;
    assign _450 = _6373;
    always @(posedge _539) begin
        if (_537)
            _6371 <= _567;
        else
            _6371 <= _450;
    end
    assign _6380 = _616 == _3048;
    assign _6378 = _565 & _570;
    assign _6381 = _6378 & _6380;
    assign _6385 = _6381 ? _597 : _6384;
    assign _6376 = _609 == _3048;
    assign _6374 = _565 & _580;
    assign _6377 = _6374 & _6376;
    assign _6386 = _6377 ? _577 : _6385;
    assign _451 = _6386;
    always @(posedge _539) begin
        if (_537)
            _6384 <= _567;
        else
            _6384 <= _451;
    end
    assign _6393 = _616 == _3061;
    assign _6391 = _565 & _570;
    assign _6394 = _6391 & _6393;
    assign _6398 = _6394 ? _597 : _6397;
    assign _6389 = _609 == _3061;
    assign _6387 = _565 & _580;
    assign _6390 = _6387 & _6389;
    assign _6399 = _6390 ? _577 : _6398;
    assign _452 = _6399;
    always @(posedge _539) begin
        if (_537)
            _6397 <= _567;
        else
            _6397 <= _452;
    end
    assign _6406 = _616 == _3074;
    assign _6404 = _565 & _570;
    assign _6407 = _6404 & _6406;
    assign _6411 = _6407 ? _597 : _6410;
    assign _6402 = _609 == _3074;
    assign _6400 = _565 & _580;
    assign _6403 = _6400 & _6402;
    assign _6412 = _6403 ? _577 : _6411;
    assign _453 = _6412;
    always @(posedge _539) begin
        if (_537)
            _6410 <= _567;
        else
            _6410 <= _453;
    end
    assign _6419 = _616 == _3087;
    assign _6417 = _565 & _570;
    assign _6420 = _6417 & _6419;
    assign _6424 = _6420 ? _597 : _6423;
    assign _6415 = _609 == _3087;
    assign _6413 = _565 & _580;
    assign _6416 = _6413 & _6415;
    assign _6425 = _6416 ? _577 : _6424;
    assign _454 = _6425;
    always @(posedge _539) begin
        if (_537)
            _6423 <= _567;
        else
            _6423 <= _454;
    end
    assign _6432 = _616 == _3100;
    assign _6430 = _565 & _570;
    assign _6433 = _6430 & _6432;
    assign _6437 = _6433 ? _597 : _6436;
    assign _6428 = _609 == _3100;
    assign _6426 = _565 & _580;
    assign _6429 = _6426 & _6428;
    assign _6438 = _6429 ? _577 : _6437;
    assign _455 = _6438;
    always @(posedge _539) begin
        if (_537)
            _6436 <= _567;
        else
            _6436 <= _455;
    end
    assign _6445 = _616 == _3113;
    assign _6443 = _565 & _570;
    assign _6446 = _6443 & _6445;
    assign _6450 = _6446 ? _597 : _6449;
    assign _6441 = _609 == _3113;
    assign _6439 = _565 & _580;
    assign _6442 = _6439 & _6441;
    assign _6451 = _6442 ? _577 : _6450;
    assign _456 = _6451;
    always @(posedge _539) begin
        if (_537)
            _6449 <= _567;
        else
            _6449 <= _456;
    end
    assign _6458 = _616 == _3126;
    assign _6456 = _565 & _570;
    assign _6459 = _6456 & _6458;
    assign _6463 = _6459 ? _597 : _6462;
    assign _6454 = _609 == _3126;
    assign _6452 = _565 & _580;
    assign _6455 = _6452 & _6454;
    assign _6464 = _6455 ? _577 : _6463;
    assign _457 = _6464;
    always @(posedge _539) begin
        if (_537)
            _6462 <= _567;
        else
            _6462 <= _457;
    end
    assign _6471 = _616 == _3139;
    assign _6469 = _565 & _570;
    assign _6472 = _6469 & _6471;
    assign _6476 = _6472 ? _597 : _6475;
    assign _6467 = _609 == _3139;
    assign _6465 = _565 & _580;
    assign _6468 = _6465 & _6467;
    assign _6477 = _6468 ? _577 : _6476;
    assign _458 = _6477;
    always @(posedge _539) begin
        if (_537)
            _6475 <= _567;
        else
            _6475 <= _458;
    end
    assign _6484 = _616 == _3152;
    assign _6482 = _565 & _570;
    assign _6485 = _6482 & _6484;
    assign _6489 = _6485 ? _597 : _6488;
    assign _6480 = _609 == _3152;
    assign _6478 = _565 & _580;
    assign _6481 = _6478 & _6480;
    assign _6490 = _6481 ? _577 : _6489;
    assign _459 = _6490;
    always @(posedge _539) begin
        if (_537)
            _6488 <= _567;
        else
            _6488 <= _459;
    end
    assign _6497 = _616 == _3165;
    assign _6495 = _565 & _570;
    assign _6498 = _6495 & _6497;
    assign _6502 = _6498 ? _597 : _6501;
    assign _6493 = _609 == _3165;
    assign _6491 = _565 & _580;
    assign _6494 = _6491 & _6493;
    assign _6503 = _6494 ? _577 : _6502;
    assign _460 = _6503;
    always @(posedge _539) begin
        if (_537)
            _6501 <= _567;
        else
            _6501 <= _460;
    end
    assign _6510 = _616 == _3178;
    assign _6508 = _565 & _570;
    assign _6511 = _6508 & _6510;
    assign _6515 = _6511 ? _597 : _6514;
    assign _6506 = _609 == _3178;
    assign _6504 = _565 & _580;
    assign _6507 = _6504 & _6506;
    assign _6516 = _6507 ? _577 : _6515;
    assign _461 = _6516;
    always @(posedge _539) begin
        if (_537)
            _6514 <= _567;
        else
            _6514 <= _461;
    end
    assign _6523 = _616 == _3191;
    assign _6521 = _565 & _570;
    assign _6524 = _6521 & _6523;
    assign _6528 = _6524 ? _597 : _6527;
    assign _6519 = _609 == _3191;
    assign _6517 = _565 & _580;
    assign _6520 = _6517 & _6519;
    assign _6529 = _6520 ? _577 : _6528;
    assign _462 = _6529;
    always @(posedge _539) begin
        if (_537)
            _6527 <= _567;
        else
            _6527 <= _462;
    end
    assign _6536 = _616 == _3204;
    assign _6534 = _565 & _570;
    assign _6537 = _6534 & _6536;
    assign _6541 = _6537 ? _597 : _6540;
    assign _6532 = _609 == _3204;
    assign _6530 = _565 & _580;
    assign _6533 = _6530 & _6532;
    assign _6542 = _6533 ? _577 : _6541;
    assign _463 = _6542;
    always @(posedge _539) begin
        if (_537)
            _6540 <= _567;
        else
            _6540 <= _463;
    end
    assign _6549 = _616 == _3217;
    assign _6547 = _565 & _570;
    assign _6550 = _6547 & _6549;
    assign _6554 = _6550 ? _597 : _6553;
    assign _6545 = _609 == _3217;
    assign _6543 = _565 & _580;
    assign _6546 = _6543 & _6545;
    assign _6555 = _6546 ? _577 : _6554;
    assign _464 = _6555;
    always @(posedge _539) begin
        if (_537)
            _6553 <= _567;
        else
            _6553 <= _464;
    end
    assign _6562 = _616 == _3230;
    assign _6560 = _565 & _570;
    assign _6563 = _6560 & _6562;
    assign _6567 = _6563 ? _597 : _6566;
    assign _6558 = _609 == _3230;
    assign _6556 = _565 & _580;
    assign _6559 = _6556 & _6558;
    assign _6568 = _6559 ? _577 : _6567;
    assign _465 = _6568;
    always @(posedge _539) begin
        if (_537)
            _6566 <= _567;
        else
            _6566 <= _465;
    end
    assign _6575 = _616 == _3243;
    assign _6573 = _565 & _570;
    assign _6576 = _6573 & _6575;
    assign _6580 = _6576 ? _597 : _6579;
    assign _6571 = _609 == _3243;
    assign _6569 = _565 & _580;
    assign _6572 = _6569 & _6571;
    assign _6581 = _6572 ? _577 : _6580;
    assign _466 = _6581;
    always @(posedge _539) begin
        if (_537)
            _6579 <= _567;
        else
            _6579 <= _466;
    end
    assign _6588 = _616 == _3256;
    assign _6586 = _565 & _570;
    assign _6589 = _6586 & _6588;
    assign _6593 = _6589 ? _597 : _6592;
    assign _6584 = _609 == _3256;
    assign _6582 = _565 & _580;
    assign _6585 = _6582 & _6584;
    assign _6594 = _6585 ? _577 : _6593;
    assign _467 = _6594;
    always @(posedge _539) begin
        if (_537)
            _6592 <= _567;
        else
            _6592 <= _467;
    end
    assign _6601 = _616 == _3269;
    assign _6599 = _565 & _570;
    assign _6602 = _6599 & _6601;
    assign _6606 = _6602 ? _597 : _6605;
    assign _6597 = _609 == _3269;
    assign _6595 = _565 & _580;
    assign _6598 = _6595 & _6597;
    assign _6607 = _6598 ? _577 : _6606;
    assign _468 = _6607;
    always @(posedge _539) begin
        if (_537)
            _6605 <= _567;
        else
            _6605 <= _468;
    end
    assign _6614 = _616 == _3282;
    assign _6612 = _565 & _570;
    assign _6615 = _6612 & _6614;
    assign _6619 = _6615 ? _597 : _6618;
    assign _6610 = _609 == _3282;
    assign _6608 = _565 & _580;
    assign _6611 = _6608 & _6610;
    assign _6620 = _6611 ? _577 : _6619;
    assign _469 = _6620;
    always @(posedge _539) begin
        if (_537)
            _6618 <= _567;
        else
            _6618 <= _469;
    end
    assign _6627 = _616 == _3295;
    assign _6625 = _565 & _570;
    assign _6628 = _6625 & _6627;
    assign _6632 = _6628 ? _597 : _6631;
    assign _6623 = _609 == _3295;
    assign _6621 = _565 & _580;
    assign _6624 = _6621 & _6623;
    assign _6633 = _6624 ? _577 : _6632;
    assign _470 = _6633;
    always @(posedge _539) begin
        if (_537)
            _6631 <= _567;
        else
            _6631 <= _470;
    end
    assign _6640 = _616 == _3308;
    assign _6638 = _565 & _570;
    assign _6641 = _6638 & _6640;
    assign _6645 = _6641 ? _597 : _6644;
    assign _6636 = _609 == _3308;
    assign _6634 = _565 & _580;
    assign _6637 = _6634 & _6636;
    assign _6646 = _6637 ? _577 : _6645;
    assign _471 = _6646;
    always @(posedge _539) begin
        if (_537)
            _6644 <= _567;
        else
            _6644 <= _471;
    end
    assign _6653 = _616 == _3321;
    assign _6651 = _565 & _570;
    assign _6654 = _6651 & _6653;
    assign _6658 = _6654 ? _597 : _6657;
    assign _6649 = _609 == _3321;
    assign _6647 = _565 & _580;
    assign _6650 = _6647 & _6649;
    assign _6659 = _6650 ? _577 : _6658;
    assign _472 = _6659;
    always @(posedge _539) begin
        if (_537)
            _6657 <= _567;
        else
            _6657 <= _472;
    end
    assign _6666 = _616 == _3334;
    assign _6664 = _565 & _570;
    assign _6667 = _6664 & _6666;
    assign _6671 = _6667 ? _597 : _6670;
    assign _6662 = _609 == _3334;
    assign _6660 = _565 & _580;
    assign _6663 = _6660 & _6662;
    assign _6672 = _6663 ? _577 : _6671;
    assign _473 = _6672;
    always @(posedge _539) begin
        if (_537)
            _6670 <= _567;
        else
            _6670 <= _473;
    end
    assign _6679 = _616 == _3347;
    assign _6677 = _565 & _570;
    assign _6680 = _6677 & _6679;
    assign _6684 = _6680 ? _597 : _6683;
    assign _6675 = _609 == _3347;
    assign _6673 = _565 & _580;
    assign _6676 = _6673 & _6675;
    assign _6685 = _6676 ? _577 : _6684;
    assign _474 = _6685;
    always @(posedge _539) begin
        if (_537)
            _6683 <= _567;
        else
            _6683 <= _474;
    end
    assign _6692 = _616 == _3360;
    assign _6690 = _565 & _570;
    assign _6693 = _6690 & _6692;
    assign _6697 = _6693 ? _597 : _6696;
    assign _6688 = _609 == _3360;
    assign _6686 = _565 & _580;
    assign _6689 = _6686 & _6688;
    assign _6698 = _6689 ? _577 : _6697;
    assign _475 = _6698;
    always @(posedge _539) begin
        if (_537)
            _6696 <= _567;
        else
            _6696 <= _475;
    end
    assign _6705 = _616 == _3373;
    assign _6703 = _565 & _570;
    assign _6706 = _6703 & _6705;
    assign _6710 = _6706 ? _597 : _6709;
    assign _6701 = _609 == _3373;
    assign _6699 = _565 & _580;
    assign _6702 = _6699 & _6701;
    assign _6711 = _6702 ? _577 : _6710;
    assign _476 = _6711;
    always @(posedge _539) begin
        if (_537)
            _6709 <= _567;
        else
            _6709 <= _476;
    end
    assign _6718 = _616 == _3386;
    assign _6716 = _565 & _570;
    assign _6719 = _6716 & _6718;
    assign _6723 = _6719 ? _597 : _6722;
    assign _6714 = _609 == _3386;
    assign _6712 = _565 & _580;
    assign _6715 = _6712 & _6714;
    assign _6724 = _6715 ? _577 : _6723;
    assign _477 = _6724;
    always @(posedge _539) begin
        if (_537)
            _6722 <= _567;
        else
            _6722 <= _477;
    end
    assign _6731 = _616 == _3399;
    assign _6729 = _565 & _570;
    assign _6732 = _6729 & _6731;
    assign _6736 = _6732 ? _597 : _6735;
    assign _6727 = _609 == _3399;
    assign _6725 = _565 & _580;
    assign _6728 = _6725 & _6727;
    assign _6737 = _6728 ? _577 : _6736;
    assign _478 = _6737;
    always @(posedge _539) begin
        if (_537)
            _6735 <= _567;
        else
            _6735 <= _478;
    end
    assign _6744 = _616 == _3412;
    assign _6742 = _565 & _570;
    assign _6745 = _6742 & _6744;
    assign _6749 = _6745 ? _597 : _6748;
    assign _6740 = _609 == _3412;
    assign _6738 = _565 & _580;
    assign _6741 = _6738 & _6740;
    assign _6750 = _6741 ? _577 : _6749;
    assign _479 = _6750;
    always @(posedge _539) begin
        if (_537)
            _6748 <= _567;
        else
            _6748 <= _479;
    end
    assign _6757 = _616 == _3425;
    assign _6755 = _565 & _570;
    assign _6758 = _6755 & _6757;
    assign _6762 = _6758 ? _597 : _6761;
    assign _6753 = _609 == _3425;
    assign _6751 = _565 & _580;
    assign _6754 = _6751 & _6753;
    assign _6763 = _6754 ? _577 : _6762;
    assign _480 = _6763;
    always @(posedge _539) begin
        if (_537)
            _6761 <= _567;
        else
            _6761 <= _480;
    end
    assign _6770 = _616 == _3438;
    assign _6768 = _565 & _570;
    assign _6771 = _6768 & _6770;
    assign _6775 = _6771 ? _597 : _6774;
    assign _6766 = _609 == _3438;
    assign _6764 = _565 & _580;
    assign _6767 = _6764 & _6766;
    assign _6776 = _6767 ? _577 : _6775;
    assign _481 = _6776;
    always @(posedge _539) begin
        if (_537)
            _6774 <= _567;
        else
            _6774 <= _481;
    end
    assign _6783 = _616 == _3451;
    assign _6781 = _565 & _570;
    assign _6784 = _6781 & _6783;
    assign _6788 = _6784 ? _597 : _6787;
    assign _6779 = _609 == _3451;
    assign _6777 = _565 & _580;
    assign _6780 = _6777 & _6779;
    assign _6789 = _6780 ? _577 : _6788;
    assign _482 = _6789;
    always @(posedge _539) begin
        if (_537)
            _6787 <= _567;
        else
            _6787 <= _482;
    end
    assign _6796 = _616 == _3464;
    assign _6794 = _565 & _570;
    assign _6797 = _6794 & _6796;
    assign _6801 = _6797 ? _597 : _6800;
    assign _6792 = _609 == _3464;
    assign _6790 = _565 & _580;
    assign _6793 = _6790 & _6792;
    assign _6802 = _6793 ? _577 : _6801;
    assign _483 = _6802;
    always @(posedge _539) begin
        if (_537)
            _6800 <= _567;
        else
            _6800 <= _483;
    end
    assign _6809 = _616 == _3477;
    assign _6807 = _565 & _570;
    assign _6810 = _6807 & _6809;
    assign _6814 = _6810 ? _597 : _6813;
    assign _6805 = _609 == _3477;
    assign _6803 = _565 & _580;
    assign _6806 = _6803 & _6805;
    assign _6815 = _6806 ? _577 : _6814;
    assign _484 = _6815;
    always @(posedge _539) begin
        if (_537)
            _6813 <= _567;
        else
            _6813 <= _484;
    end
    assign _6822 = _616 == _3490;
    assign _6820 = _565 & _570;
    assign _6823 = _6820 & _6822;
    assign _6827 = _6823 ? _597 : _6826;
    assign _6818 = _609 == _3490;
    assign _6816 = _565 & _580;
    assign _6819 = _6816 & _6818;
    assign _6828 = _6819 ? _577 : _6827;
    assign _485 = _6828;
    always @(posedge _539) begin
        if (_537)
            _6826 <= _567;
        else
            _6826 <= _485;
    end
    assign _6835 = _616 == _3503;
    assign _6833 = _565 & _570;
    assign _6836 = _6833 & _6835;
    assign _6840 = _6836 ? _597 : _6839;
    assign _6831 = _609 == _3503;
    assign _6829 = _565 & _580;
    assign _6832 = _6829 & _6831;
    assign _6841 = _6832 ? _577 : _6840;
    assign _486 = _6841;
    always @(posedge _539) begin
        if (_537)
            _6839 <= _567;
        else
            _6839 <= _486;
    end
    assign _6848 = _616 == _3516;
    assign _6846 = _565 & _570;
    assign _6849 = _6846 & _6848;
    assign _6853 = _6849 ? _597 : _6852;
    assign _6844 = _609 == _3516;
    assign _6842 = _565 & _580;
    assign _6845 = _6842 & _6844;
    assign _6854 = _6845 ? _577 : _6853;
    assign _487 = _6854;
    always @(posedge _539) begin
        if (_537)
            _6852 <= _567;
        else
            _6852 <= _487;
    end
    assign _6861 = _616 == _3529;
    assign _6859 = _565 & _570;
    assign _6862 = _6859 & _6861;
    assign _6866 = _6862 ? _597 : _6865;
    assign _6857 = _609 == _3529;
    assign _6855 = _565 & _580;
    assign _6858 = _6855 & _6857;
    assign _6867 = _6858 ? _577 : _6866;
    assign _488 = _6867;
    always @(posedge _539) begin
        if (_537)
            _6865 <= _567;
        else
            _6865 <= _488;
    end
    assign _6874 = _616 == _3542;
    assign _6872 = _565 & _570;
    assign _6875 = _6872 & _6874;
    assign _6879 = _6875 ? _597 : _6878;
    assign _6870 = _609 == _3542;
    assign _6868 = _565 & _580;
    assign _6871 = _6868 & _6870;
    assign _6880 = _6871 ? _577 : _6879;
    assign _489 = _6880;
    always @(posedge _539) begin
        if (_537)
            _6878 <= _567;
        else
            _6878 <= _489;
    end
    assign _6887 = _616 == _3555;
    assign _6885 = _565 & _570;
    assign _6888 = _6885 & _6887;
    assign _6892 = _6888 ? _597 : _6891;
    assign _6883 = _609 == _3555;
    assign _6881 = _565 & _580;
    assign _6884 = _6881 & _6883;
    assign _6893 = _6884 ? _577 : _6892;
    assign _490 = _6893;
    always @(posedge _539) begin
        if (_537)
            _6891 <= _567;
        else
            _6891 <= _490;
    end
    assign _6900 = _616 == _3568;
    assign _6898 = _565 & _570;
    assign _6901 = _6898 & _6900;
    assign _6905 = _6901 ? _597 : _6904;
    assign _6896 = _609 == _3568;
    assign _6894 = _565 & _580;
    assign _6897 = _6894 & _6896;
    assign _6906 = _6897 ? _577 : _6905;
    assign _491 = _6906;
    always @(posedge _539) begin
        if (_537)
            _6904 <= _567;
        else
            _6904 <= _491;
    end
    assign _6913 = _616 == _3581;
    assign _6911 = _565 & _570;
    assign _6914 = _6911 & _6913;
    assign _6918 = _6914 ? _597 : _6917;
    assign _6909 = _609 == _3581;
    assign _6907 = _565 & _580;
    assign _6910 = _6907 & _6909;
    assign _6919 = _6910 ? _577 : _6918;
    assign _492 = _6919;
    always @(posedge _539) begin
        if (_537)
            _6917 <= _567;
        else
            _6917 <= _492;
    end
    assign _6926 = _616 == _3594;
    assign _6924 = _565 & _570;
    assign _6927 = _6924 & _6926;
    assign _6931 = _6927 ? _597 : _6930;
    assign _6922 = _609 == _3594;
    assign _6920 = _565 & _580;
    assign _6923 = _6920 & _6922;
    assign _6932 = _6923 ? _577 : _6931;
    assign _493 = _6932;
    always @(posedge _539) begin
        if (_537)
            _6930 <= _567;
        else
            _6930 <= _493;
    end
    assign _6939 = _616 == _3607;
    assign _6937 = _565 & _570;
    assign _6940 = _6937 & _6939;
    assign _6944 = _6940 ? _597 : _6943;
    assign _6935 = _609 == _3607;
    assign _6933 = _565 & _580;
    assign _6936 = _6933 & _6935;
    assign _6945 = _6936 ? _577 : _6944;
    assign _494 = _6945;
    always @(posedge _539) begin
        if (_537)
            _6943 <= _567;
        else
            _6943 <= _494;
    end
    assign _6952 = _616 == _3620;
    assign _6950 = _565 & _570;
    assign _6953 = _6950 & _6952;
    assign _6957 = _6953 ? _597 : _6956;
    assign _6948 = _609 == _3620;
    assign _6946 = _565 & _580;
    assign _6949 = _6946 & _6948;
    assign _6958 = _6949 ? _577 : _6957;
    assign _495 = _6958;
    always @(posedge _539) begin
        if (_537)
            _6956 <= _567;
        else
            _6956 <= _495;
    end
    assign _6965 = _616 == _3633;
    assign _6963 = _565 & _570;
    assign _6966 = _6963 & _6965;
    assign _6970 = _6966 ? _597 : _6969;
    assign _6961 = _609 == _3633;
    assign _6959 = _565 & _580;
    assign _6962 = _6959 & _6961;
    assign _6971 = _6962 ? _577 : _6970;
    assign _496 = _6971;
    always @(posedge _539) begin
        if (_537)
            _6969 <= _567;
        else
            _6969 <= _496;
    end
    assign _6978 = _616 == _3646;
    assign _6976 = _565 & _570;
    assign _6979 = _6976 & _6978;
    assign _6983 = _6979 ? _597 : _6982;
    assign _6974 = _609 == _3646;
    assign _6972 = _565 & _580;
    assign _6975 = _6972 & _6974;
    assign _6984 = _6975 ? _577 : _6983;
    assign _497 = _6984;
    always @(posedge _539) begin
        if (_537)
            _6982 <= _567;
        else
            _6982 <= _497;
    end
    assign _6991 = _616 == _3659;
    assign _6989 = _565 & _570;
    assign _6992 = _6989 & _6991;
    assign _6996 = _6992 ? _597 : _6995;
    assign _6987 = _609 == _3659;
    assign _6985 = _565 & _580;
    assign _6988 = _6985 & _6987;
    assign _6997 = _6988 ? _577 : _6996;
    assign _498 = _6997;
    always @(posedge _539) begin
        if (_537)
            _6995 <= _567;
        else
            _6995 <= _498;
    end
    assign _7004 = _616 == _3672;
    assign _7002 = _565 & _570;
    assign _7005 = _7002 & _7004;
    assign _7009 = _7005 ? _597 : _7008;
    assign _7000 = _609 == _3672;
    assign _6998 = _565 & _580;
    assign _7001 = _6998 & _7000;
    assign _7010 = _7001 ? _577 : _7009;
    assign _499 = _7010;
    always @(posedge _539) begin
        if (_537)
            _7008 <= _567;
        else
            _7008 <= _499;
    end
    assign _7017 = _616 == _3685;
    assign _7015 = _565 & _570;
    assign _7018 = _7015 & _7017;
    assign _7022 = _7018 ? _597 : _7021;
    assign _7013 = _609 == _3685;
    assign _7011 = _565 & _580;
    assign _7014 = _7011 & _7013;
    assign _7023 = _7014 ? _577 : _7022;
    assign _500 = _7023;
    always @(posedge _539) begin
        if (_537)
            _7021 <= _567;
        else
            _7021 <= _500;
    end
    assign _7030 = _616 == _3698;
    assign _7028 = _565 & _570;
    assign _7031 = _7028 & _7030;
    assign _7035 = _7031 ? _597 : _7034;
    assign _7026 = _609 == _3698;
    assign _7024 = _565 & _580;
    assign _7027 = _7024 & _7026;
    assign _7036 = _7027 ? _577 : _7035;
    assign _501 = _7036;
    always @(posedge _539) begin
        if (_537)
            _7034 <= _567;
        else
            _7034 <= _501;
    end
    assign _7043 = _616 == _3711;
    assign _7041 = _565 & _570;
    assign _7044 = _7041 & _7043;
    assign _7048 = _7044 ? _597 : _7047;
    assign _7039 = _609 == _3711;
    assign _7037 = _565 & _580;
    assign _7040 = _7037 & _7039;
    assign _7049 = _7040 ? _577 : _7048;
    assign _502 = _7049;
    always @(posedge _539) begin
        if (_537)
            _7047 <= _567;
        else
            _7047 <= _502;
    end
    assign _7056 = _616 == _3724;
    assign _7054 = _565 & _570;
    assign _7057 = _7054 & _7056;
    assign _7061 = _7057 ? _597 : _7060;
    assign _7052 = _609 == _3724;
    assign _7050 = _565 & _580;
    assign _7053 = _7050 & _7052;
    assign _7062 = _7053 ? _577 : _7061;
    assign _503 = _7062;
    always @(posedge _539) begin
        if (_537)
            _7060 <= _567;
        else
            _7060 <= _503;
    end
    assign _7069 = _616 == _3737;
    assign _7067 = _565 & _570;
    assign _7070 = _7067 & _7069;
    assign _7074 = _7070 ? _597 : _7073;
    assign _7065 = _609 == _3737;
    assign _7063 = _565 & _580;
    assign _7066 = _7063 & _7065;
    assign _7075 = _7066 ? _577 : _7074;
    assign _504 = _7075;
    always @(posedge _539) begin
        if (_537)
            _7073 <= _567;
        else
            _7073 <= _504;
    end
    assign _7082 = _616 == _3750;
    assign _7080 = _565 & _570;
    assign _7083 = _7080 & _7082;
    assign _7087 = _7083 ? _597 : _7086;
    assign _7078 = _609 == _3750;
    assign _7076 = _565 & _580;
    assign _7079 = _7076 & _7078;
    assign _7088 = _7079 ? _577 : _7087;
    assign _505 = _7088;
    always @(posedge _539) begin
        if (_537)
            _7086 <= _567;
        else
            _7086 <= _505;
    end
    assign _7095 = _616 == _3763;
    assign _7093 = _565 & _570;
    assign _7096 = _7093 & _7095;
    assign _7100 = _7096 ? _597 : _7099;
    assign _7091 = _609 == _3763;
    assign _7089 = _565 & _580;
    assign _7092 = _7089 & _7091;
    assign _7101 = _7092 ? _577 : _7100;
    assign _506 = _7101;
    always @(posedge _539) begin
        if (_537)
            _7099 <= _567;
        else
            _7099 <= _506;
    end
    assign _7108 = _616 == _3776;
    assign _7106 = _565 & _570;
    assign _7109 = _7106 & _7108;
    assign _7113 = _7109 ? _597 : _7112;
    assign _7104 = _609 == _3776;
    assign _7102 = _565 & _580;
    assign _7105 = _7102 & _7104;
    assign _7114 = _7105 ? _577 : _7113;
    assign _507 = _7114;
    always @(posedge _539) begin
        if (_537)
            _7112 <= _567;
        else
            _7112 <= _507;
    end
    assign _7121 = _616 == _3789;
    assign _7119 = _565 & _570;
    assign _7122 = _7119 & _7121;
    assign _7126 = _7122 ? _597 : _7125;
    assign _7117 = _609 == _3789;
    assign _7115 = _565 & _580;
    assign _7118 = _7115 & _7117;
    assign _7127 = _7118 ? _577 : _7126;
    assign _508 = _7127;
    always @(posedge _539) begin
        if (_537)
            _7125 <= _567;
        else
            _7125 <= _508;
    end
    assign _7134 = _616 == _3802;
    assign _7132 = _565 & _570;
    assign _7135 = _7132 & _7134;
    assign _7139 = _7135 ? _597 : _7138;
    assign _7130 = _609 == _3802;
    assign _7128 = _565 & _580;
    assign _7131 = _7128 & _7130;
    assign _7140 = _7131 ? _577 : _7139;
    assign _509 = _7140;
    always @(posedge _539) begin
        if (_537)
            _7138 <= _567;
        else
            _7138 <= _509;
    end
    assign _7147 = _616 == _3815;
    assign _7145 = _565 & _570;
    assign _7148 = _7145 & _7147;
    assign _7152 = _7148 ? _597 : _7151;
    assign _7143 = _609 == _3815;
    assign _7141 = _565 & _580;
    assign _7144 = _7141 & _7143;
    assign _7153 = _7144 ? _577 : _7152;
    assign _510 = _7153;
    always @(posedge _539) begin
        if (_537)
            _7151 <= _567;
        else
            _7151 <= _510;
    end
    assign _7160 = _616 == _3828;
    assign _7158 = _565 & _570;
    assign _7161 = _7158 & _7160;
    assign _7165 = _7161 ? _597 : _7164;
    assign _7156 = _609 == _3828;
    assign _7154 = _565 & _580;
    assign _7157 = _7154 & _7156;
    assign _7166 = _7157 ? _577 : _7165;
    assign _511 = _7166;
    always @(posedge _539) begin
        if (_537)
            _7164 <= _567;
        else
            _7164 <= _511;
    end
    assign _7173 = _616 == _3841;
    assign _7171 = _565 & _570;
    assign _7174 = _7171 & _7173;
    assign _7178 = _7174 ? _597 : _7177;
    assign _7169 = _609 == _3841;
    assign _7167 = _565 & _580;
    assign _7170 = _7167 & _7169;
    assign _7179 = _7170 ? _577 : _7178;
    assign _512 = _7179;
    always @(posedge _539) begin
        if (_537)
            _7177 <= _567;
        else
            _7177 <= _512;
    end
    assign _7186 = _616 == _3854;
    assign _7184 = _565 & _570;
    assign _7187 = _7184 & _7186;
    assign _7191 = _7187 ? _597 : _7190;
    assign _7182 = _609 == _3854;
    assign _7180 = _565 & _580;
    assign _7183 = _7180 & _7182;
    assign _7192 = _7183 ? _577 : _7191;
    assign _513 = _7192;
    always @(posedge _539) begin
        if (_537)
            _7190 <= _567;
        else
            _7190 <= _513;
    end
    assign _7199 = _616 == _3867;
    assign _7197 = _565 & _570;
    assign _7200 = _7197 & _7199;
    assign _7204 = _7200 ? _597 : _7203;
    assign _7195 = _609 == _3867;
    assign _7193 = _565 & _580;
    assign _7196 = _7193 & _7195;
    assign _7205 = _7196 ? _577 : _7204;
    assign _514 = _7205;
    always @(posedge _539) begin
        if (_537)
            _7203 <= _567;
        else
            _7203 <= _514;
    end
    assign _7212 = _616 == _3880;
    assign _7210 = _565 & _570;
    assign _7213 = _7210 & _7212;
    assign _7217 = _7213 ? _597 : _7216;
    assign _7208 = _609 == _3880;
    assign _7206 = _565 & _580;
    assign _7209 = _7206 & _7208;
    assign _7218 = _7209 ? _577 : _7217;
    assign _515 = _7218;
    always @(posedge _539) begin
        if (_537)
            _7216 <= _567;
        else
            _7216 <= _515;
    end
    assign _7225 = _616 == _3893;
    assign _7223 = _565 & _570;
    assign _7226 = _7223 & _7225;
    assign _7230 = _7226 ? _597 : _7229;
    assign _7221 = _609 == _3893;
    assign _7219 = _565 & _580;
    assign _7222 = _7219 & _7221;
    assign _7231 = _7222 ? _577 : _7230;
    assign _516 = _7231;
    always @(posedge _539) begin
        if (_537)
            _7229 <= _567;
        else
            _7229 <= _516;
    end
    assign _7238 = _616 == _3906;
    assign _7236 = _565 & _570;
    assign _7239 = _7236 & _7238;
    assign _7243 = _7239 ? _597 : _7242;
    assign _7234 = _609 == _3906;
    assign _7232 = _565 & _580;
    assign _7235 = _7232 & _7234;
    assign _7244 = _7235 ? _577 : _7243;
    assign _517 = _7244;
    always @(posedge _539) begin
        if (_537)
            _7242 <= _567;
        else
            _7242 <= _517;
    end
    assign _7251 = _616 == _3919;
    assign _7249 = _565 & _570;
    assign _7252 = _7249 & _7251;
    assign _7256 = _7252 ? _597 : _7255;
    assign _7247 = _609 == _3919;
    assign _7245 = _565 & _580;
    assign _7248 = _7245 & _7247;
    assign _7257 = _7248 ? _577 : _7256;
    assign _518 = _7257;
    always @(posedge _539) begin
        if (_537)
            _7255 <= _567;
        else
            _7255 <= _518;
    end
    assign _7264 = _616 == _3935;
    assign _7262 = _565 & _570;
    assign _7265 = _7262 & _7264;
    assign _7269 = _7265 ? _597 : _7268;
    assign _7260 = _609 == _3935;
    assign _7258 = _565 & _580;
    assign _7261 = _7258 & _7260;
    assign _7270 = _7261 ? _577 : _7269;
    assign _519 = _7270;
    always @(posedge _539) begin
        if (_537)
            _7268 <= _567;
        else
            _7268 <= _519;
    end
    assign _7297 = _7285 + _3919;
    assign _7298 = _7295 ? _7297 : _7285;
    assign _7271 = _565 & _570;
    assign _7300 = _7271 ? _3935 : _7298;
    assign _7302 = _548 ? _3935 : _7300;
    assign _520 = _7302;
    always @(posedge _539) begin
        if (_537)
            _7285 <= _3935;
        else
            _7285 <= _520;
    end
    always @* begin
        case (_7285)
        0:
            _7286 <= _7268;
        1:
            _7286 <= _7255;
        2:
            _7286 <= _7242;
        3:
            _7286 <= _7229;
        4:
            _7286 <= _7216;
        5:
            _7286 <= _7203;
        6:
            _7286 <= _7190;
        7:
            _7286 <= _7177;
        8:
            _7286 <= _7164;
        9:
            _7286 <= _7151;
        10:
            _7286 <= _7138;
        11:
            _7286 <= _7125;
        12:
            _7286 <= _7112;
        13:
            _7286 <= _7099;
        14:
            _7286 <= _7086;
        15:
            _7286 <= _7073;
        16:
            _7286 <= _7060;
        17:
            _7286 <= _7047;
        18:
            _7286 <= _7034;
        19:
            _7286 <= _7021;
        20:
            _7286 <= _7008;
        21:
            _7286 <= _6995;
        22:
            _7286 <= _6982;
        23:
            _7286 <= _6969;
        24:
            _7286 <= _6956;
        25:
            _7286 <= _6943;
        26:
            _7286 <= _6930;
        27:
            _7286 <= _6917;
        28:
            _7286 <= _6904;
        29:
            _7286 <= _6891;
        30:
            _7286 <= _6878;
        31:
            _7286 <= _6865;
        32:
            _7286 <= _6852;
        33:
            _7286 <= _6839;
        34:
            _7286 <= _6826;
        35:
            _7286 <= _6813;
        36:
            _7286 <= _6800;
        37:
            _7286 <= _6787;
        38:
            _7286 <= _6774;
        39:
            _7286 <= _6761;
        40:
            _7286 <= _6748;
        41:
            _7286 <= _6735;
        42:
            _7286 <= _6722;
        43:
            _7286 <= _6709;
        44:
            _7286 <= _6696;
        45:
            _7286 <= _6683;
        46:
            _7286 <= _6670;
        47:
            _7286 <= _6657;
        48:
            _7286 <= _6644;
        49:
            _7286 <= _6631;
        50:
            _7286 <= _6618;
        51:
            _7286 <= _6605;
        52:
            _7286 <= _6592;
        53:
            _7286 <= _6579;
        54:
            _7286 <= _6566;
        55:
            _7286 <= _6553;
        56:
            _7286 <= _6540;
        57:
            _7286 <= _6527;
        58:
            _7286 <= _6514;
        59:
            _7286 <= _6501;
        60:
            _7286 <= _6488;
        61:
            _7286 <= _6475;
        62:
            _7286 <= _6462;
        63:
            _7286 <= _6449;
        64:
            _7286 <= _6436;
        65:
            _7286 <= _6423;
        66:
            _7286 <= _6410;
        67:
            _7286 <= _6397;
        68:
            _7286 <= _6384;
        69:
            _7286 <= _6371;
        70:
            _7286 <= _6358;
        71:
            _7286 <= _6345;
        72:
            _7286 <= _6332;
        73:
            _7286 <= _6319;
        74:
            _7286 <= _6306;
        75:
            _7286 <= _6293;
        76:
            _7286 <= _6280;
        77:
            _7286 <= _6267;
        78:
            _7286 <= _6254;
        79:
            _7286 <= _6241;
        80:
            _7286 <= _6228;
        81:
            _7286 <= _6215;
        82:
            _7286 <= _6202;
        83:
            _7286 <= _6189;
        84:
            _7286 <= _6176;
        85:
            _7286 <= _6163;
        86:
            _7286 <= _6150;
        87:
            _7286 <= _6137;
        88:
            _7286 <= _6124;
        89:
            _7286 <= _6111;
        90:
            _7286 <= _6098;
        91:
            _7286 <= _6085;
        92:
            _7286 <= _6072;
        93:
            _7286 <= _6059;
        94:
            _7286 <= _6046;
        95:
            _7286 <= _6033;
        96:
            _7286 <= _6020;
        97:
            _7286 <= _6007;
        98:
            _7286 <= _5994;
        99:
            _7286 <= _5981;
        100:
            _7286 <= _5968;
        101:
            _7286 <= _5955;
        102:
            _7286 <= _5942;
        103:
            _7286 <= _5929;
        104:
            _7286 <= _5916;
        105:
            _7286 <= _5903;
        106:
            _7286 <= _5890;
        107:
            _7286 <= _5877;
        108:
            _7286 <= _5864;
        109:
            _7286 <= _5851;
        110:
            _7286 <= _5838;
        111:
            _7286 <= _5825;
        112:
            _7286 <= _5812;
        113:
            _7286 <= _5799;
        114:
            _7286 <= _5786;
        115:
            _7286 <= _5773;
        116:
            _7286 <= _5760;
        117:
            _7286 <= _5747;
        118:
            _7286 <= _5734;
        119:
            _7286 <= _5721;
        120:
            _7286 <= _5708;
        121:
            _7286 <= _5695;
        122:
            _7286 <= _5682;
        123:
            _7286 <= _5669;
        124:
            _7286 <= _5656;
        125:
            _7286 <= _5643;
        126:
            _7286 <= _5630;
        127:
            _7286 <= _5617;
        128:
            _7286 <= _5604;
        129:
            _7286 <= _5591;
        130:
            _7286 <= _5578;
        131:
            _7286 <= _5565;
        132:
            _7286 <= _5552;
        133:
            _7286 <= _5539;
        134:
            _7286 <= _5526;
        135:
            _7286 <= _5513;
        136:
            _7286 <= _5500;
        137:
            _7286 <= _5487;
        138:
            _7286 <= _5474;
        139:
            _7286 <= _5461;
        140:
            _7286 <= _5448;
        141:
            _7286 <= _5435;
        142:
            _7286 <= _5422;
        143:
            _7286 <= _5409;
        144:
            _7286 <= _5396;
        145:
            _7286 <= _5383;
        146:
            _7286 <= _5370;
        147:
            _7286 <= _5357;
        148:
            _7286 <= _5344;
        149:
            _7286 <= _5331;
        150:
            _7286 <= _5318;
        151:
            _7286 <= _5305;
        152:
            _7286 <= _5292;
        153:
            _7286 <= _5279;
        154:
            _7286 <= _5266;
        155:
            _7286 <= _5253;
        156:
            _7286 <= _5240;
        157:
            _7286 <= _5227;
        158:
            _7286 <= _5214;
        159:
            _7286 <= _5201;
        160:
            _7286 <= _5188;
        161:
            _7286 <= _5175;
        162:
            _7286 <= _5162;
        163:
            _7286 <= _5149;
        164:
            _7286 <= _5136;
        165:
            _7286 <= _5123;
        166:
            _7286 <= _5110;
        167:
            _7286 <= _5097;
        168:
            _7286 <= _5084;
        169:
            _7286 <= _5071;
        170:
            _7286 <= _5058;
        171:
            _7286 <= _5045;
        172:
            _7286 <= _5032;
        173:
            _7286 <= _5019;
        174:
            _7286 <= _5006;
        175:
            _7286 <= _4993;
        176:
            _7286 <= _4980;
        177:
            _7286 <= _4967;
        178:
            _7286 <= _4954;
        179:
            _7286 <= _4941;
        180:
            _7286 <= _4928;
        181:
            _7286 <= _4915;
        182:
            _7286 <= _4902;
        183:
            _7286 <= _4889;
        184:
            _7286 <= _4876;
        185:
            _7286 <= _4863;
        186:
            _7286 <= _4850;
        187:
            _7286 <= _4837;
        188:
            _7286 <= _4824;
        189:
            _7286 <= _4811;
        190:
            _7286 <= _4798;
        191:
            _7286 <= _4785;
        192:
            _7286 <= _4772;
        193:
            _7286 <= _4759;
        194:
            _7286 <= _4746;
        195:
            _7286 <= _4733;
        196:
            _7286 <= _4720;
        197:
            _7286 <= _4707;
        198:
            _7286 <= _4694;
        199:
            _7286 <= _4681;
        200:
            _7286 <= _4668;
        201:
            _7286 <= _4655;
        202:
            _7286 <= _4642;
        203:
            _7286 <= _4629;
        204:
            _7286 <= _4616;
        205:
            _7286 <= _4603;
        206:
            _7286 <= _4590;
        207:
            _7286 <= _4577;
        208:
            _7286 <= _4564;
        209:
            _7286 <= _4551;
        210:
            _7286 <= _4538;
        211:
            _7286 <= _4525;
        212:
            _7286 <= _4512;
        213:
            _7286 <= _4499;
        214:
            _7286 <= _4486;
        215:
            _7286 <= _4473;
        216:
            _7286 <= _4460;
        217:
            _7286 <= _4447;
        218:
            _7286 <= _4434;
        219:
            _7286 <= _4421;
        220:
            _7286 <= _4408;
        221:
            _7286 <= _4395;
        222:
            _7286 <= _4382;
        223:
            _7286 <= _4369;
        224:
            _7286 <= _4356;
        225:
            _7286 <= _4343;
        226:
            _7286 <= _4330;
        227:
            _7286 <= _4317;
        228:
            _7286 <= _4304;
        229:
            _7286 <= _4291;
        230:
            _7286 <= _4278;
        231:
            _7286 <= _4265;
        232:
            _7286 <= _4252;
        233:
            _7286 <= _4239;
        234:
            _7286 <= _4226;
        235:
            _7286 <= _4213;
        236:
            _7286 <= _4200;
        237:
            _7286 <= _4187;
        238:
            _7286 <= _4174;
        239:
            _7286 <= _4161;
        240:
            _7286 <= _4148;
        241:
            _7286 <= _4135;
        242:
            _7286 <= _4122;
        243:
            _7286 <= _4109;
        244:
            _7286 <= _4096;
        245:
            _7286 <= _4083;
        246:
            _7286 <= _4070;
        247:
            _7286 <= _4057;
        248:
            _7286 <= _4044;
        249:
            _7286 <= _4031;
        250:
            _7286 <= _4018;
        251:
            _7286 <= _4005;
        252:
            _7286 <= _3992;
        253:
            _7286 <= _3979;
        254:
            _7286 <= _3966;
        default:
            _7286 <= _3953;
        endcase
    end
    assign _522 = id;
    assign _7304 = _7303 ? _522 : _7282;
    assign _7306 = _548 ? _567 : _7304;
    assign _523 = _7306;
    always @(posedge _539) begin
        if (_537)
            _7282 <= _567;
        else
            _7282 <= _523;
    end
    assign _7287 = _7282 < _7286;
    assign _7288 = ~ _7287;
    assign _7308 = _616 + _3919;
    assign _615 = _609 + _3919;
    assign _7310 = _565 ? _7309 : _609;
    assign _7312 = _548 ? _3935 : _7310;
    assign _524 = _7312;
    always @(posedge _539) begin
        if (_537)
            _609 <= _3935;
        else
            _609 <= _524;
    end
    assign _594 = _577 < _592;
    assign _595 = _594 ? _592 : _577;
    assign _526 = range_to;
    assign _592 = _526 + _7353;
    assign _593 = _580 ? _592 : _577;
    assign _589 = _569 & _573;
    assign _590 = _589 & _578;
    assign _596 = _590 ? _595 : _593;
    assign _587 = ~ _573;
    assign _588 = _569 & _587;
    assign _597 = _588 ? _592 : _596;
    assign _7313 = _565 ? _597 : _577;
    assign _7315 = _548 ? _567 : _7313;
    assign _527 = _7315;
    always @(posedge _539) begin
        if (_537)
            _577 <= _567;
        else
            _577 <= _527;
    end
    assign _529 = range_from;
    assign _578 = _529 < _577;
    assign _579 = ~ _578;
    assign _572 = 1'b0;
    assign _7316 = _569 ? vdd : _573;
    assign _7317 = _565 ? _7316 : _573;
    assign _7319 = _548 ? _572 : _7317;
    assign _530 = _7319;
    always @(posedge _539) begin
        if (_537)
            _573 <= _572;
        else
            _573 <= _530;
    end
    assign _574 = _569 & _573;
    assign _580 = _574 & _579;
    assign _616 = _580 ? _615 : _609;
    assign _7309 = _570 ? _7308 : _616;
    assign _7320 = _565 & _570;
    assign _7321 = _7320 ? _7309 : _7275;
    assign _7323 = _548 ? _3935 : _7321;
    assign _531 = _7323;
    always @(posedge _539) begin
        if (_537)
            _7275 <= _3935;
        else
            _7275 <= _531;
    end
    assign _7277 = _7275 == _3935;
    assign _7278 = ~ _7277;
    assign _7272 = _558 & _561;
    assign _7279 = _7272 & _7278;
    assign _7289 = _7279 & _7288;
    assign _7295 = _7289 & _7294;
    assign _7325 = ~ _7295;
    assign _552 = 2'b00;
    assign _557 = 2'b01;
    assign _555 = 2'b10;
    assign _533 = id_last;
    assign _535 = id_valid;
    assign _537 = clear;
    assign _539 = clock;
    assign vdd = 1'b1;
    assign _7328 = _7326 ? _572 : _561;
    assign _7329 = _7303 ? vdd : _7328;
    assign _7331 = _548 ? _572 : _7329;
    assign _540 = _7331;
    always @(posedge _539) begin
        if (_537)
            _561 <= _572;
        else
            _561 <= _540;
    end
    assign _562 = ~ _561;
    assign _563 = _558 & _562;
    assign _7303 = _563 & _535;
    assign _7335 = _7303 ? _533 : _7334;
    assign _7337 = _548 ? _572 : _7335;
    assign _541 = _7337;
    always @(posedge _539) begin
        if (_537)
            _7334 <= _572;
        else
            _7334 <= _541;
    end
    assign _7339 = _7326 & _7334;
    assign _7340 = _7339 ? _555 : _554;
    assign _543 = range_last;
    assign _545 = range_valid;
    assign _569 = _565 & _545;
    assign _570 = _569 & _543;
    assign _565 = _554 == _552;
    assign _7338 = _565 & _570;
    assign _7341 = _7338 ? _557 : _7340;
    assign _7342 = _548 ? _552 : _7341;
    assign _546 = _7342;
    always @(posedge _539) begin
        if (_537)
            _554 <= _552;
        else
            _554 <= _546;
    end
    assign _558 = _554 == _557;
    assign _7324 = _558 & _561;
    assign _7326 = _7324 & _7325;
    assign _7349 = _7326 & _7348;
    assign _7355 = _7349 ? _7354 : _7352;
    assign _548 = load;
    assign _7357 = _548 ? _567 : _7355;
    assign _549 = _7357;
    always @(posedge _539) begin
        if (_537)
            _7352 <= _567;
        else
            _7352 <= _549;
    end
    assign part1_result = _7352;
    assign part2_result = _568;
    assign range_ready = _565;
    assign id_ready = _563;
    assign done_ = _556;
    assign phase = _554;

endmodule
