module day3_opt_c (
    data,
    start,
    clear,
    clock,
    k,
    length,
    result,
    done_
);

    input [511:0] data;
    input start;
    input clear;
    input clock;
    input [3:0] k;
    input [7:0] length;
    output [63:0] result;
    output done_;

    wire _42;
    wire _45;
    wire _46;
    wire _1;
    reg _43;
    wire [3:0] _50;
    wire [3:0] _737;
    wire _738;
    wire _739;
    wire [3:0] _734;
    wire _735;
    wire _733;
    wire _736;
    wire _740;
    wire [3:0] _741;
    wire [3:0] _607;
    wire _608;
    wire _609;
    wire _605;
    wire _603;
    wire _606;
    wire _610;
    wire [3:0] _611;
    wire [3:0] _477;
    wire _478;
    wire _479;
    wire _475;
    wire _473;
    wire _476;
    wire _480;
    wire [3:0] _481;
    wire [3:0] _347;
    wire _348;
    wire _349;
    wire _345;
    wire _343;
    wire _346;
    wire _350;
    wire [3:0] _351;
    wire [3:0] _352;
    wire [3:0] _482;
    wire [3:0] _612;
    wire [3:0] _742;
    wire [7:0] _58;
    wire [7:0] _59;
    reg [3:0] _188;
    wire _53;
    wire [3:0] _189;
    wire [3:0] _190;
    wire [3:0] _743;
    wire [3:0] _3;
    reg [3:0] _51;
    wire [59:0] _985;
    wire [63:0] _986;
    wire [63:0] _982;
    wire [127:0] _983;
    wire [63:0] _984;
    wire [63:0] _987;
    wire [3:0] _727;
    wire _730;
    wire _731;
    wire [3:0] _613;
    wire _614;
    wire _725;
    wire _726;
    wire _732;
    wire [3:0] _752;
    wire [3:0] _597;
    wire _600;
    wire _601;
    wire _484;
    wire _595;
    wire _596;
    wire _602;
    wire [3:0] _728;
    wire [3:0] _467;
    wire _470;
    wire _471;
    wire _354;
    wire _465;
    wire _466;
    wire _472;
    wire [3:0] _598;
    wire [3:0] _336;
    wire _340;
    wire _341;
    wire _214;
    wire _334;
    wire _335;
    wire _342;
    wire [3:0] _468;
    wire [3:0] _469;
    wire [3:0] _599;
    wire [3:0] _729;
    wire [3:0] _753;
    wire [7:0] _747;
    wire [7:0] _748;
    reg [3:0] _749;
    wire _745;
    wire [3:0] _750;
    wire [3:0] _751;
    wire [3:0] _754;
    wire [3:0] _4;
    reg [3:0] _339;
    wire [63:0] _979;
    wire [127:0] _976;
    wire [63:0] _977;
    wire [63:0] _980;
    wire [3:0] _719;
    wire _722;
    wire _723;
    wire [3:0] _616;
    wire _617;
    wire _717;
    wire _718;
    wire _724;
    wire [3:0] _763;
    wire [3:0] _589;
    wire _592;
    wire _593;
    wire _487;
    wire _587;
    wire _588;
    wire _594;
    wire [3:0] _720;
    wire [3:0] _459;
    wire _462;
    wire _463;
    wire _357;
    wire _457;
    wire _458;
    wire _464;
    wire [3:0] _590;
    wire [3:0] _327;
    wire _331;
    wire _332;
    wire _217;
    wire _325;
    wire _326;
    wire _333;
    wire [3:0] _460;
    wire [3:0] _461;
    wire [3:0] _591;
    wire [3:0] _721;
    wire [3:0] _764;
    wire [7:0] _758;
    wire [7:0] _759;
    reg [3:0] _760;
    wire _756;
    wire [3:0] _761;
    wire [3:0] _762;
    wire [3:0] _765;
    wire [3:0] _5;
    reg [3:0] _330;
    wire [63:0] _972;
    wire [127:0] _969;
    wire [63:0] _970;
    wire [63:0] _973;
    wire [3:0] _711;
    wire _714;
    wire _715;
    wire [3:0] _619;
    wire _620;
    wire _709;
    wire _710;
    wire _716;
    wire [3:0] _774;
    wire [3:0] _581;
    wire _584;
    wire _585;
    wire _490;
    wire _579;
    wire _580;
    wire _586;
    wire [3:0] _712;
    wire [3:0] _451;
    wire _454;
    wire _455;
    wire _360;
    wire _449;
    wire _450;
    wire _456;
    wire [3:0] _582;
    wire [3:0] _318;
    wire _322;
    wire _323;
    wire _220;
    wire _316;
    wire _317;
    wire _324;
    wire [3:0] _452;
    wire [3:0] _453;
    wire [3:0] _583;
    wire [3:0] _713;
    wire [3:0] _775;
    wire [7:0] _769;
    wire [7:0] _770;
    reg [3:0] _771;
    wire _767;
    wire [3:0] _772;
    wire [3:0] _773;
    wire [3:0] _776;
    wire [3:0] _6;
    reg [3:0] _321;
    wire [63:0] _965;
    wire [127:0] _962;
    wire [63:0] _963;
    wire [63:0] _966;
    wire [3:0] _703;
    wire _706;
    wire _707;
    wire [3:0] _622;
    wire _623;
    wire _701;
    wire _702;
    wire _708;
    wire [3:0] _785;
    wire [3:0] _573;
    wire _576;
    wire _577;
    wire _493;
    wire _571;
    wire _572;
    wire _578;
    wire [3:0] _704;
    wire [3:0] _443;
    wire _446;
    wire _447;
    wire _363;
    wire _441;
    wire _442;
    wire _448;
    wire [3:0] _574;
    wire [3:0] _309;
    wire _313;
    wire _314;
    wire _223;
    wire _307;
    wire _308;
    wire _315;
    wire [3:0] _444;
    wire [3:0] _445;
    wire [3:0] _575;
    wire [3:0] _705;
    wire [3:0] _786;
    wire [7:0] _780;
    wire [7:0] _781;
    reg [3:0] _782;
    wire _778;
    wire [3:0] _783;
    wire [3:0] _784;
    wire [3:0] _787;
    wire [3:0] _7;
    reg [3:0] _312;
    wire [63:0] _958;
    wire [127:0] _955;
    wire [63:0] _956;
    wire [63:0] _959;
    wire [3:0] _695;
    wire _698;
    wire _699;
    wire [3:0] _625;
    wire _626;
    wire _693;
    wire _694;
    wire _700;
    wire [3:0] _796;
    wire [3:0] _565;
    wire _568;
    wire _569;
    wire _496;
    wire _563;
    wire _564;
    wire _570;
    wire [3:0] _696;
    wire [3:0] _435;
    wire _438;
    wire _439;
    wire _366;
    wire _433;
    wire _434;
    wire _440;
    wire [3:0] _566;
    wire [3:0] _300;
    wire _304;
    wire _305;
    wire _226;
    wire _298;
    wire _299;
    wire _306;
    wire [3:0] _436;
    wire [3:0] _437;
    wire [3:0] _567;
    wire [3:0] _697;
    wire [3:0] _797;
    wire [7:0] _791;
    wire [7:0] _792;
    reg [3:0] _793;
    wire _789;
    wire [3:0] _794;
    wire [3:0] _795;
    wire [3:0] _798;
    wire [3:0] _8;
    reg [3:0] _303;
    wire [63:0] _951;
    wire [127:0] _948;
    wire [63:0] _949;
    wire [63:0] _952;
    wire [3:0] _687;
    wire _690;
    wire _691;
    wire [3:0] _628;
    wire _629;
    wire _685;
    wire _686;
    wire _692;
    wire [3:0] _807;
    wire [3:0] _557;
    wire _560;
    wire _561;
    wire _499;
    wire _555;
    wire _556;
    wire _562;
    wire [3:0] _688;
    wire [3:0] _427;
    wire _430;
    wire _431;
    wire _369;
    wire _425;
    wire _426;
    wire _432;
    wire [3:0] _558;
    wire [3:0] _291;
    wire _295;
    wire _296;
    wire _229;
    wire _289;
    wire _290;
    wire _297;
    wire [3:0] _428;
    wire [3:0] _429;
    wire [3:0] _559;
    wire [3:0] _689;
    wire [3:0] _808;
    wire [7:0] _802;
    wire [7:0] _803;
    reg [3:0] _804;
    wire _800;
    wire [3:0] _805;
    wire [3:0] _806;
    wire [3:0] _809;
    wire [3:0] _9;
    reg [3:0] _294;
    wire [63:0] _944;
    wire [127:0] _941;
    wire [63:0] _942;
    wire [63:0] _945;
    wire [3:0] _679;
    wire _682;
    wire _683;
    wire [3:0] _631;
    wire _632;
    wire _677;
    wire _678;
    wire _684;
    wire [3:0] _818;
    wire [3:0] _549;
    wire _552;
    wire _553;
    wire _502;
    wire _547;
    wire _548;
    wire _554;
    wire [3:0] _680;
    wire [3:0] _419;
    wire _422;
    wire _423;
    wire _372;
    wire _417;
    wire _418;
    wire _424;
    wire [3:0] _550;
    wire [3:0] _282;
    wire _286;
    wire _287;
    wire _232;
    wire _280;
    wire _281;
    wire _288;
    wire [3:0] _420;
    wire [3:0] _421;
    wire [3:0] _551;
    wire [3:0] _681;
    wire [3:0] _819;
    wire [7:0] _813;
    wire [7:0] _814;
    reg [3:0] _815;
    wire _811;
    wire [3:0] _816;
    wire [3:0] _817;
    wire [3:0] _820;
    wire [3:0] _10;
    reg [3:0] _285;
    wire [63:0] _937;
    wire [127:0] _934;
    wire [63:0] _935;
    wire [63:0] _938;
    wire [3:0] _671;
    wire _674;
    wire _675;
    wire [3:0] _634;
    wire _635;
    wire _669;
    wire _670;
    wire _676;
    wire [3:0] _829;
    wire [3:0] _541;
    wire _544;
    wire _545;
    wire _505;
    wire _539;
    wire _540;
    wire _546;
    wire [3:0] _672;
    wire [3:0] _411;
    wire _414;
    wire _415;
    wire _375;
    wire _409;
    wire _410;
    wire _416;
    wire [3:0] _542;
    wire [3:0] _273;
    wire _277;
    wire _278;
    wire _235;
    wire _271;
    wire _272;
    wire _279;
    wire [3:0] _412;
    wire [3:0] _413;
    wire [3:0] _543;
    wire [3:0] _673;
    wire [3:0] _830;
    wire [7:0] _824;
    wire [7:0] _825;
    reg [3:0] _826;
    wire _822;
    wire [3:0] _827;
    wire [3:0] _828;
    wire [3:0] _831;
    wire [3:0] _11;
    reg [3:0] _276;
    wire [63:0] _930;
    wire [127:0] _927;
    wire [63:0] _928;
    wire [63:0] _931;
    wire [3:0] _663;
    wire _666;
    wire _667;
    wire [3:0] _637;
    wire _638;
    wire _661;
    wire _662;
    wire _668;
    wire [3:0] _840;
    wire [3:0] _533;
    wire _536;
    wire _537;
    wire _508;
    wire _531;
    wire _532;
    wire _538;
    wire [3:0] _664;
    wire [3:0] _403;
    wire _406;
    wire _407;
    wire _378;
    wire _401;
    wire _402;
    wire _408;
    wire [3:0] _534;
    wire [3:0] _264;
    wire _268;
    wire _269;
    wire _238;
    wire _262;
    wire _263;
    wire _270;
    wire [3:0] _404;
    wire [3:0] _405;
    wire [3:0] _535;
    wire [3:0] _665;
    wire [3:0] _841;
    wire [7:0] _835;
    wire [7:0] _836;
    reg [3:0] _837;
    wire _833;
    wire [3:0] _838;
    wire [3:0] _839;
    wire [3:0] _842;
    wire [3:0] _12;
    reg [3:0] _267;
    wire [63:0] _923;
    wire [127:0] _920;
    wire [63:0] _921;
    wire [63:0] _924;
    wire [3:0] _655;
    wire _658;
    wire _659;
    wire [3:0] _640;
    wire _641;
    wire _653;
    wire _654;
    wire _660;
    wire [3:0] _851;
    wire [3:0] _525;
    wire _528;
    wire _529;
    wire _511;
    wire _523;
    wire _524;
    wire _530;
    wire [3:0] _656;
    wire [3:0] _395;
    wire _398;
    wire _399;
    wire _381;
    wire _393;
    wire _394;
    wire _400;
    wire [3:0] _526;
    wire [3:0] _255;
    wire _259;
    wire _260;
    wire _241;
    wire _253;
    wire _254;
    wire _261;
    wire [3:0] _396;
    wire [3:0] _397;
    wire [3:0] _527;
    wire [3:0] _657;
    wire [3:0] _852;
    wire [7:0] _846;
    wire [7:0] _847;
    reg [3:0] _848;
    wire _844;
    wire [3:0] _849;
    wire [3:0] _850;
    wire [3:0] _853;
    wire [3:0] _13;
    reg [3:0] _258;
    wire [63:0] _916;
    wire [127:0] _913;
    wire [63:0] _914;
    wire [63:0] _917;
    wire [7:0] _646;
    reg [3:0] _647;
    wire _650;
    wire _651;
    wire _644;
    wire _652;
    wire [3:0] _860;
    wire [7:0] _516;
    reg [3:0] _517;
    wire _520;
    wire _521;
    wire _514;
    wire _522;
    wire [3:0] _648;
    wire [7:0] _386;
    reg [3:0] _387;
    wire _390;
    wire _391;
    wire _384;
    wire _392;
    wire [3:0] _518;
    reg [3:0] _246;
    wire _250;
    wire _251;
    wire _244;
    wire _252;
    wire [3:0] _388;
    wire [7:0] _206;
    wire _207;
    wire _208;
    wire _209;
    wire [3:0] _389;
    wire _203;
    wire _204;
    wire _205;
    wire [3:0] _519;
    wire _199;
    wire _200;
    wire _201;
    wire [3:0] _649;
    wire _195;
    wire _196;
    wire _197;
    wire [3:0] _861;
    wire [3:0] _187;
    wire [3:0] _186;
    wire [3:0] _185;
    wire [3:0] _184;
    wire [3:0] _183;
    wire [3:0] _182;
    wire [3:0] _181;
    wire [3:0] _180;
    wire [3:0] _179;
    wire [3:0] _178;
    wire [3:0] _177;
    wire [3:0] _176;
    wire [3:0] _175;
    wire [3:0] _174;
    wire [3:0] _173;
    wire [3:0] _172;
    wire [3:0] _171;
    wire [3:0] _170;
    wire [3:0] _169;
    wire [3:0] _168;
    wire [3:0] _167;
    wire [3:0] _166;
    wire [3:0] _165;
    wire [3:0] _164;
    wire [3:0] _163;
    wire [3:0] _162;
    wire [3:0] _161;
    wire [3:0] _160;
    wire [3:0] _159;
    wire [3:0] _158;
    wire [3:0] _157;
    wire [3:0] _156;
    wire [3:0] _155;
    wire [3:0] _154;
    wire [3:0] _153;
    wire [3:0] _152;
    wire [3:0] _151;
    wire [3:0] _150;
    wire [3:0] _149;
    wire [3:0] _148;
    wire [3:0] _147;
    wire [3:0] _146;
    wire [3:0] _145;
    wire [3:0] _144;
    wire [3:0] _143;
    wire [3:0] _142;
    wire [3:0] _141;
    wire [3:0] _140;
    wire [3:0] _139;
    wire [3:0] _138;
    wire [3:0] _137;
    wire [3:0] _136;
    wire [3:0] _135;
    wire [3:0] _134;
    wire [3:0] _133;
    wire [3:0] _132;
    wire [3:0] _131;
    wire [3:0] _130;
    wire [3:0] _129;
    wire [3:0] _128;
    wire [3:0] _127;
    wire [3:0] _126;
    wire [3:0] _125;
    wire [3:0] _124;
    wire [3:0] _123;
    wire [3:0] _122;
    wire [3:0] _121;
    wire [3:0] _120;
    wire [3:0] _119;
    wire [3:0] _118;
    wire [3:0] _117;
    wire [3:0] _116;
    wire [3:0] _115;
    wire [3:0] _114;
    wire [3:0] _113;
    wire [3:0] _112;
    wire [3:0] _111;
    wire [3:0] _110;
    wire [3:0] _109;
    wire [3:0] _108;
    wire [3:0] _107;
    wire [3:0] _106;
    wire [3:0] _105;
    wire [3:0] _104;
    wire [3:0] _103;
    wire [3:0] _102;
    wire [3:0] _101;
    wire [3:0] _100;
    wire [3:0] _99;
    wire [3:0] _98;
    wire [3:0] _97;
    wire [3:0] _96;
    wire [3:0] _95;
    wire [3:0] _94;
    wire [3:0] _93;
    wire [3:0] _92;
    wire [3:0] _91;
    wire [3:0] _90;
    wire [3:0] _89;
    wire [3:0] _88;
    wire [3:0] _87;
    wire [3:0] _86;
    wire [3:0] _85;
    wire [3:0] _84;
    wire [3:0] _83;
    wire [3:0] _82;
    wire [3:0] _81;
    wire [3:0] _80;
    wire [3:0] _79;
    wire [3:0] _78;
    wire [3:0] _77;
    wire [3:0] _76;
    wire [3:0] _75;
    wire [3:0] _74;
    wire [3:0] _73;
    wire [3:0] _72;
    wire [3:0] _71;
    wire [3:0] _70;
    wire [3:0] _69;
    wire [3:0] _68;
    wire [3:0] _67;
    wire [3:0] _66;
    wire [3:0] _65;
    wire [3:0] _64;
    wire [3:0] _63;
    wire [3:0] _62;
    wire [3:0] _61;
    wire [511:0] _15;
    wire [3:0] _60;
    reg [3:0] _857;
    wire _855;
    wire [3:0] _858;
    wire [3:0] _859;
    wire [3:0] _862;
    wire [3:0] _16;
    reg [3:0] _249;
    wire [63:0] _910;
    wire [63:0] _908;
    wire _907;
    wire [63:0] _911;
    wire _905;
    wire [63:0] _918;
    wire _903;
    wire [63:0] _925;
    wire _901;
    wire [63:0] _932;
    wire _899;
    wire [63:0] _939;
    wire _897;
    wire [63:0] _946;
    wire _895;
    wire [63:0] _953;
    wire _893;
    wire [63:0] _960;
    wire _891;
    wire [63:0] _967;
    wire _889;
    wire [63:0] _974;
    wire _887;
    wire [63:0] _981;
    wire _18;
    wire [1:0] _35;
    wire _36;
    wire [1:0] _37;
    wire [1:0] _879;
    wire vdd;
    wire _20;
    wire _22;
    wire [7:0] _869;
    wire [7:0] _871;
    wire [7:0] _864;
    wire [7:0] _865;
    wire [7:0] _872;
    wire [7:0] _23;
    reg [7:0] _193;
    wire _867;
    wire [1:0] _881;
    wire [3:0] _25;
    wire [7:0] _56;
    wire [7:0] _27;
    wire [7:0] _57;
    wire _874;
    wire [1:0] _877;
    wire [1:0] _878;
    wire _48;
    wire [1:0] _882;
    wire [1:0] _28;
    reg [1:0] _34;
    wire _38;
    wire _39;
    wire _40;
    wire [3:0] _883;
    wire [3:0] _29;
    reg [3:0] _213;
    wire _885;
    wire [63:0] _988;
    assign _42 = 1'b0;
    assign _45 = _40 ? _42 : _43;
    assign _46 = _36 ? vdd : _45;
    assign _1 = _46;
    always @(posedge _22) begin
        if (_20)
            _43 <= _42;
        else
            _43 <= _1;
    end
    assign _50 = 4'b0000;
    assign _737 = _732 ? _729 : _727;
    assign _738 = _737 < _612;
    assign _739 = ~ _738;
    assign _734 = 4'b1011;
    assign _735 = _734 < _213;
    assign _733 = _614 ? _732 : _42;
    assign _736 = _733 & _735;
    assign _740 = _736 & _739;
    assign _741 = _740 ? _737 : _612;
    assign _607 = _602 ? _599 : _597;
    assign _608 = _607 < _482;
    assign _609 = ~ _608;
    assign _605 = _734 < _213;
    assign _603 = _484 ? _602 : _42;
    assign _606 = _603 & _605;
    assign _610 = _606 & _609;
    assign _611 = _610 ? _607 : _482;
    assign _477 = _472 ? _469 : _467;
    assign _478 = _477 < _352;
    assign _479 = ~ _478;
    assign _475 = _734 < _213;
    assign _473 = _354 ? _472 : _42;
    assign _476 = _473 & _475;
    assign _480 = _476 & _479;
    assign _481 = _480 ? _477 : _352;
    assign _347 = _342 ? _339 : _336;
    assign _348 = _347 < _51;
    assign _349 = ~ _348;
    assign _345 = _734 < _213;
    assign _343 = _214 ? _342 : _42;
    assign _346 = _343 & _345;
    assign _350 = _346 & _349;
    assign _351 = _350 ? _347 : _51;
    assign _352 = _209 ? _351 : _51;
    assign _482 = _205 ? _481 : _352;
    assign _612 = _201 ? _611 : _482;
    assign _742 = _197 ? _741 : _612;
    assign _58 = 8'b00001011;
    assign _59 = _57 + _58;
    always @* begin
        case (_59)
        0:
            _188 <= _60;
        1:
            _188 <= _61;
        2:
            _188 <= _62;
        3:
            _188 <= _63;
        4:
            _188 <= _64;
        5:
            _188 <= _65;
        6:
            _188 <= _66;
        7:
            _188 <= _67;
        8:
            _188 <= _68;
        9:
            _188 <= _69;
        10:
            _188 <= _70;
        11:
            _188 <= _71;
        12:
            _188 <= _72;
        13:
            _188 <= _73;
        14:
            _188 <= _74;
        15:
            _188 <= _75;
        16:
            _188 <= _76;
        17:
            _188 <= _77;
        18:
            _188 <= _78;
        19:
            _188 <= _79;
        20:
            _188 <= _80;
        21:
            _188 <= _81;
        22:
            _188 <= _82;
        23:
            _188 <= _83;
        24:
            _188 <= _84;
        25:
            _188 <= _85;
        26:
            _188 <= _86;
        27:
            _188 <= _87;
        28:
            _188 <= _88;
        29:
            _188 <= _89;
        30:
            _188 <= _90;
        31:
            _188 <= _91;
        32:
            _188 <= _92;
        33:
            _188 <= _93;
        34:
            _188 <= _94;
        35:
            _188 <= _95;
        36:
            _188 <= _96;
        37:
            _188 <= _97;
        38:
            _188 <= _98;
        39:
            _188 <= _99;
        40:
            _188 <= _100;
        41:
            _188 <= _101;
        42:
            _188 <= _102;
        43:
            _188 <= _103;
        44:
            _188 <= _104;
        45:
            _188 <= _105;
        46:
            _188 <= _106;
        47:
            _188 <= _107;
        48:
            _188 <= _108;
        49:
            _188 <= _109;
        50:
            _188 <= _110;
        51:
            _188 <= _111;
        52:
            _188 <= _112;
        53:
            _188 <= _113;
        54:
            _188 <= _114;
        55:
            _188 <= _115;
        56:
            _188 <= _116;
        57:
            _188 <= _117;
        58:
            _188 <= _118;
        59:
            _188 <= _119;
        60:
            _188 <= _120;
        61:
            _188 <= _121;
        62:
            _188 <= _122;
        63:
            _188 <= _123;
        64:
            _188 <= _124;
        65:
            _188 <= _125;
        66:
            _188 <= _126;
        67:
            _188 <= _127;
        68:
            _188 <= _128;
        69:
            _188 <= _129;
        70:
            _188 <= _130;
        71:
            _188 <= _131;
        72:
            _188 <= _132;
        73:
            _188 <= _133;
        74:
            _188 <= _134;
        75:
            _188 <= _135;
        76:
            _188 <= _136;
        77:
            _188 <= _137;
        78:
            _188 <= _138;
        79:
            _188 <= _139;
        80:
            _188 <= _140;
        81:
            _188 <= _141;
        82:
            _188 <= _142;
        83:
            _188 <= _143;
        84:
            _188 <= _144;
        85:
            _188 <= _145;
        86:
            _188 <= _146;
        87:
            _188 <= _147;
        88:
            _188 <= _148;
        89:
            _188 <= _149;
        90:
            _188 <= _150;
        91:
            _188 <= _151;
        92:
            _188 <= _152;
        93:
            _188 <= _153;
        94:
            _188 <= _154;
        95:
            _188 <= _155;
        96:
            _188 <= _156;
        97:
            _188 <= _157;
        98:
            _188 <= _158;
        99:
            _188 <= _159;
        100:
            _188 <= _160;
        101:
            _188 <= _161;
        102:
            _188 <= _162;
        103:
            _188 <= _163;
        104:
            _188 <= _164;
        105:
            _188 <= _165;
        106:
            _188 <= _166;
        107:
            _188 <= _167;
        108:
            _188 <= _168;
        109:
            _188 <= _169;
        110:
            _188 <= _170;
        111:
            _188 <= _171;
        112:
            _188 <= _172;
        113:
            _188 <= _173;
        114:
            _188 <= _174;
        115:
            _188 <= _175;
        116:
            _188 <= _176;
        117:
            _188 <= _177;
        118:
            _188 <= _178;
        119:
            _188 <= _179;
        120:
            _188 <= _180;
        121:
            _188 <= _181;
        122:
            _188 <= _182;
        123:
            _188 <= _183;
        124:
            _188 <= _184;
        125:
            _188 <= _185;
        126:
            _188 <= _186;
        default:
            _188 <= _187;
        endcase
    end
    assign _53 = _734 < _25;
    assign _189 = _53 ? _188 : _50;
    assign _190 = _40 ? _189 : _51;
    assign _743 = _48 ? _742 : _190;
    assign _3 = _743;
    always @(posedge _22) begin
        if (_20)
            _51 <= _50;
        else
            _51 <= _3;
    end
    assign _985 = 60'b000000000000000000000000000000000000000000000000000000000000;
    assign _986 = { _985,
                    _51 };
    assign _982 = 64'b0000000000000000000000000000000000000000000000000000000000001010;
    assign _983 = _981 * _982;
    assign _984 = _983[63:0];
    assign _987 = _984 + _986;
    assign _727 = _724 ? _721 : _719;
    assign _730 = _727 < _729;
    assign _731 = ~ _730;
    assign _613 = 4'b1010;
    assign _614 = _613 < _213;
    assign _725 = _617 ? _724 : _42;
    assign _726 = _725 & _614;
    assign _732 = _726 & _731;
    assign _752 = _732 ? _727 : _729;
    assign _597 = _594 ? _591 : _589;
    assign _600 = _597 < _599;
    assign _601 = ~ _600;
    assign _484 = _613 < _213;
    assign _595 = _487 ? _594 : _42;
    assign _596 = _595 & _484;
    assign _602 = _596 & _601;
    assign _728 = _602 ? _597 : _599;
    assign _467 = _464 ? _461 : _459;
    assign _470 = _467 < _469;
    assign _471 = ~ _470;
    assign _354 = _613 < _213;
    assign _465 = _357 ? _464 : _42;
    assign _466 = _465 & _354;
    assign _472 = _466 & _471;
    assign _598 = _472 ? _467 : _469;
    assign _336 = _333 ? _330 : _327;
    assign _340 = _336 < _339;
    assign _341 = ~ _340;
    assign _214 = _613 < _213;
    assign _334 = _217 ? _333 : _42;
    assign _335 = _334 & _214;
    assign _342 = _335 & _341;
    assign _468 = _342 ? _336 : _339;
    assign _469 = _209 ? _468 : _339;
    assign _599 = _205 ? _598 : _469;
    assign _729 = _201 ? _728 : _599;
    assign _753 = _197 ? _752 : _729;
    assign _747 = 8'b00001010;
    assign _748 = _57 + _747;
    always @* begin
        case (_748)
        0:
            _749 <= _60;
        1:
            _749 <= _61;
        2:
            _749 <= _62;
        3:
            _749 <= _63;
        4:
            _749 <= _64;
        5:
            _749 <= _65;
        6:
            _749 <= _66;
        7:
            _749 <= _67;
        8:
            _749 <= _68;
        9:
            _749 <= _69;
        10:
            _749 <= _70;
        11:
            _749 <= _71;
        12:
            _749 <= _72;
        13:
            _749 <= _73;
        14:
            _749 <= _74;
        15:
            _749 <= _75;
        16:
            _749 <= _76;
        17:
            _749 <= _77;
        18:
            _749 <= _78;
        19:
            _749 <= _79;
        20:
            _749 <= _80;
        21:
            _749 <= _81;
        22:
            _749 <= _82;
        23:
            _749 <= _83;
        24:
            _749 <= _84;
        25:
            _749 <= _85;
        26:
            _749 <= _86;
        27:
            _749 <= _87;
        28:
            _749 <= _88;
        29:
            _749 <= _89;
        30:
            _749 <= _90;
        31:
            _749 <= _91;
        32:
            _749 <= _92;
        33:
            _749 <= _93;
        34:
            _749 <= _94;
        35:
            _749 <= _95;
        36:
            _749 <= _96;
        37:
            _749 <= _97;
        38:
            _749 <= _98;
        39:
            _749 <= _99;
        40:
            _749 <= _100;
        41:
            _749 <= _101;
        42:
            _749 <= _102;
        43:
            _749 <= _103;
        44:
            _749 <= _104;
        45:
            _749 <= _105;
        46:
            _749 <= _106;
        47:
            _749 <= _107;
        48:
            _749 <= _108;
        49:
            _749 <= _109;
        50:
            _749 <= _110;
        51:
            _749 <= _111;
        52:
            _749 <= _112;
        53:
            _749 <= _113;
        54:
            _749 <= _114;
        55:
            _749 <= _115;
        56:
            _749 <= _116;
        57:
            _749 <= _117;
        58:
            _749 <= _118;
        59:
            _749 <= _119;
        60:
            _749 <= _120;
        61:
            _749 <= _121;
        62:
            _749 <= _122;
        63:
            _749 <= _123;
        64:
            _749 <= _124;
        65:
            _749 <= _125;
        66:
            _749 <= _126;
        67:
            _749 <= _127;
        68:
            _749 <= _128;
        69:
            _749 <= _129;
        70:
            _749 <= _130;
        71:
            _749 <= _131;
        72:
            _749 <= _132;
        73:
            _749 <= _133;
        74:
            _749 <= _134;
        75:
            _749 <= _135;
        76:
            _749 <= _136;
        77:
            _749 <= _137;
        78:
            _749 <= _138;
        79:
            _749 <= _139;
        80:
            _749 <= _140;
        81:
            _749 <= _141;
        82:
            _749 <= _142;
        83:
            _749 <= _143;
        84:
            _749 <= _144;
        85:
            _749 <= _145;
        86:
            _749 <= _146;
        87:
            _749 <= _147;
        88:
            _749 <= _148;
        89:
            _749 <= _149;
        90:
            _749 <= _150;
        91:
            _749 <= _151;
        92:
            _749 <= _152;
        93:
            _749 <= _153;
        94:
            _749 <= _154;
        95:
            _749 <= _155;
        96:
            _749 <= _156;
        97:
            _749 <= _157;
        98:
            _749 <= _158;
        99:
            _749 <= _159;
        100:
            _749 <= _160;
        101:
            _749 <= _161;
        102:
            _749 <= _162;
        103:
            _749 <= _163;
        104:
            _749 <= _164;
        105:
            _749 <= _165;
        106:
            _749 <= _166;
        107:
            _749 <= _167;
        108:
            _749 <= _168;
        109:
            _749 <= _169;
        110:
            _749 <= _170;
        111:
            _749 <= _171;
        112:
            _749 <= _172;
        113:
            _749 <= _173;
        114:
            _749 <= _174;
        115:
            _749 <= _175;
        116:
            _749 <= _176;
        117:
            _749 <= _177;
        118:
            _749 <= _178;
        119:
            _749 <= _179;
        120:
            _749 <= _180;
        121:
            _749 <= _181;
        122:
            _749 <= _182;
        123:
            _749 <= _183;
        124:
            _749 <= _184;
        125:
            _749 <= _185;
        126:
            _749 <= _186;
        default:
            _749 <= _187;
        endcase
    end
    assign _745 = _613 < _25;
    assign _750 = _745 ? _749 : _50;
    assign _751 = _40 ? _750 : _339;
    assign _754 = _48 ? _753 : _751;
    assign _4 = _754;
    always @(posedge _22) begin
        if (_20)
            _339 <= _50;
        else
            _339 <= _4;
    end
    assign _979 = { _985,
                    _339 };
    assign _976 = _974 * _982;
    assign _977 = _976[63:0];
    assign _980 = _977 + _979;
    assign _719 = _716 ? _713 : _711;
    assign _722 = _719 < _721;
    assign _723 = ~ _722;
    assign _616 = 4'b1001;
    assign _617 = _616 < _213;
    assign _717 = _620 ? _716 : _42;
    assign _718 = _717 & _617;
    assign _724 = _718 & _723;
    assign _763 = _724 ? _719 : _721;
    assign _589 = _586 ? _583 : _581;
    assign _592 = _589 < _591;
    assign _593 = ~ _592;
    assign _487 = _616 < _213;
    assign _587 = _490 ? _586 : _42;
    assign _588 = _587 & _487;
    assign _594 = _588 & _593;
    assign _720 = _594 ? _589 : _591;
    assign _459 = _456 ? _453 : _451;
    assign _462 = _459 < _461;
    assign _463 = ~ _462;
    assign _357 = _616 < _213;
    assign _457 = _360 ? _456 : _42;
    assign _458 = _457 & _357;
    assign _464 = _458 & _463;
    assign _590 = _464 ? _459 : _461;
    assign _327 = _324 ? _321 : _318;
    assign _331 = _327 < _330;
    assign _332 = ~ _331;
    assign _217 = _616 < _213;
    assign _325 = _220 ? _324 : _42;
    assign _326 = _325 & _217;
    assign _333 = _326 & _332;
    assign _460 = _333 ? _327 : _330;
    assign _461 = _209 ? _460 : _330;
    assign _591 = _205 ? _590 : _461;
    assign _721 = _201 ? _720 : _591;
    assign _764 = _197 ? _763 : _721;
    assign _758 = 8'b00001001;
    assign _759 = _57 + _758;
    always @* begin
        case (_759)
        0:
            _760 <= _60;
        1:
            _760 <= _61;
        2:
            _760 <= _62;
        3:
            _760 <= _63;
        4:
            _760 <= _64;
        5:
            _760 <= _65;
        6:
            _760 <= _66;
        7:
            _760 <= _67;
        8:
            _760 <= _68;
        9:
            _760 <= _69;
        10:
            _760 <= _70;
        11:
            _760 <= _71;
        12:
            _760 <= _72;
        13:
            _760 <= _73;
        14:
            _760 <= _74;
        15:
            _760 <= _75;
        16:
            _760 <= _76;
        17:
            _760 <= _77;
        18:
            _760 <= _78;
        19:
            _760 <= _79;
        20:
            _760 <= _80;
        21:
            _760 <= _81;
        22:
            _760 <= _82;
        23:
            _760 <= _83;
        24:
            _760 <= _84;
        25:
            _760 <= _85;
        26:
            _760 <= _86;
        27:
            _760 <= _87;
        28:
            _760 <= _88;
        29:
            _760 <= _89;
        30:
            _760 <= _90;
        31:
            _760 <= _91;
        32:
            _760 <= _92;
        33:
            _760 <= _93;
        34:
            _760 <= _94;
        35:
            _760 <= _95;
        36:
            _760 <= _96;
        37:
            _760 <= _97;
        38:
            _760 <= _98;
        39:
            _760 <= _99;
        40:
            _760 <= _100;
        41:
            _760 <= _101;
        42:
            _760 <= _102;
        43:
            _760 <= _103;
        44:
            _760 <= _104;
        45:
            _760 <= _105;
        46:
            _760 <= _106;
        47:
            _760 <= _107;
        48:
            _760 <= _108;
        49:
            _760 <= _109;
        50:
            _760 <= _110;
        51:
            _760 <= _111;
        52:
            _760 <= _112;
        53:
            _760 <= _113;
        54:
            _760 <= _114;
        55:
            _760 <= _115;
        56:
            _760 <= _116;
        57:
            _760 <= _117;
        58:
            _760 <= _118;
        59:
            _760 <= _119;
        60:
            _760 <= _120;
        61:
            _760 <= _121;
        62:
            _760 <= _122;
        63:
            _760 <= _123;
        64:
            _760 <= _124;
        65:
            _760 <= _125;
        66:
            _760 <= _126;
        67:
            _760 <= _127;
        68:
            _760 <= _128;
        69:
            _760 <= _129;
        70:
            _760 <= _130;
        71:
            _760 <= _131;
        72:
            _760 <= _132;
        73:
            _760 <= _133;
        74:
            _760 <= _134;
        75:
            _760 <= _135;
        76:
            _760 <= _136;
        77:
            _760 <= _137;
        78:
            _760 <= _138;
        79:
            _760 <= _139;
        80:
            _760 <= _140;
        81:
            _760 <= _141;
        82:
            _760 <= _142;
        83:
            _760 <= _143;
        84:
            _760 <= _144;
        85:
            _760 <= _145;
        86:
            _760 <= _146;
        87:
            _760 <= _147;
        88:
            _760 <= _148;
        89:
            _760 <= _149;
        90:
            _760 <= _150;
        91:
            _760 <= _151;
        92:
            _760 <= _152;
        93:
            _760 <= _153;
        94:
            _760 <= _154;
        95:
            _760 <= _155;
        96:
            _760 <= _156;
        97:
            _760 <= _157;
        98:
            _760 <= _158;
        99:
            _760 <= _159;
        100:
            _760 <= _160;
        101:
            _760 <= _161;
        102:
            _760 <= _162;
        103:
            _760 <= _163;
        104:
            _760 <= _164;
        105:
            _760 <= _165;
        106:
            _760 <= _166;
        107:
            _760 <= _167;
        108:
            _760 <= _168;
        109:
            _760 <= _169;
        110:
            _760 <= _170;
        111:
            _760 <= _171;
        112:
            _760 <= _172;
        113:
            _760 <= _173;
        114:
            _760 <= _174;
        115:
            _760 <= _175;
        116:
            _760 <= _176;
        117:
            _760 <= _177;
        118:
            _760 <= _178;
        119:
            _760 <= _179;
        120:
            _760 <= _180;
        121:
            _760 <= _181;
        122:
            _760 <= _182;
        123:
            _760 <= _183;
        124:
            _760 <= _184;
        125:
            _760 <= _185;
        126:
            _760 <= _186;
        default:
            _760 <= _187;
        endcase
    end
    assign _756 = _616 < _25;
    assign _761 = _756 ? _760 : _50;
    assign _762 = _40 ? _761 : _330;
    assign _765 = _48 ? _764 : _762;
    assign _5 = _765;
    always @(posedge _22) begin
        if (_20)
            _330 <= _50;
        else
            _330 <= _5;
    end
    assign _972 = { _985,
                    _330 };
    assign _969 = _967 * _982;
    assign _970 = _969[63:0];
    assign _973 = _970 + _972;
    assign _711 = _708 ? _705 : _703;
    assign _714 = _711 < _713;
    assign _715 = ~ _714;
    assign _619 = 4'b1000;
    assign _620 = _619 < _213;
    assign _709 = _623 ? _708 : _42;
    assign _710 = _709 & _620;
    assign _716 = _710 & _715;
    assign _774 = _716 ? _711 : _713;
    assign _581 = _578 ? _575 : _573;
    assign _584 = _581 < _583;
    assign _585 = ~ _584;
    assign _490 = _619 < _213;
    assign _579 = _493 ? _578 : _42;
    assign _580 = _579 & _490;
    assign _586 = _580 & _585;
    assign _712 = _586 ? _581 : _583;
    assign _451 = _448 ? _445 : _443;
    assign _454 = _451 < _453;
    assign _455 = ~ _454;
    assign _360 = _619 < _213;
    assign _449 = _363 ? _448 : _42;
    assign _450 = _449 & _360;
    assign _456 = _450 & _455;
    assign _582 = _456 ? _451 : _453;
    assign _318 = _315 ? _312 : _309;
    assign _322 = _318 < _321;
    assign _323 = ~ _322;
    assign _220 = _619 < _213;
    assign _316 = _223 ? _315 : _42;
    assign _317 = _316 & _220;
    assign _324 = _317 & _323;
    assign _452 = _324 ? _318 : _321;
    assign _453 = _209 ? _452 : _321;
    assign _583 = _205 ? _582 : _453;
    assign _713 = _201 ? _712 : _583;
    assign _775 = _197 ? _774 : _713;
    assign _769 = 8'b00001000;
    assign _770 = _57 + _769;
    always @* begin
        case (_770)
        0:
            _771 <= _60;
        1:
            _771 <= _61;
        2:
            _771 <= _62;
        3:
            _771 <= _63;
        4:
            _771 <= _64;
        5:
            _771 <= _65;
        6:
            _771 <= _66;
        7:
            _771 <= _67;
        8:
            _771 <= _68;
        9:
            _771 <= _69;
        10:
            _771 <= _70;
        11:
            _771 <= _71;
        12:
            _771 <= _72;
        13:
            _771 <= _73;
        14:
            _771 <= _74;
        15:
            _771 <= _75;
        16:
            _771 <= _76;
        17:
            _771 <= _77;
        18:
            _771 <= _78;
        19:
            _771 <= _79;
        20:
            _771 <= _80;
        21:
            _771 <= _81;
        22:
            _771 <= _82;
        23:
            _771 <= _83;
        24:
            _771 <= _84;
        25:
            _771 <= _85;
        26:
            _771 <= _86;
        27:
            _771 <= _87;
        28:
            _771 <= _88;
        29:
            _771 <= _89;
        30:
            _771 <= _90;
        31:
            _771 <= _91;
        32:
            _771 <= _92;
        33:
            _771 <= _93;
        34:
            _771 <= _94;
        35:
            _771 <= _95;
        36:
            _771 <= _96;
        37:
            _771 <= _97;
        38:
            _771 <= _98;
        39:
            _771 <= _99;
        40:
            _771 <= _100;
        41:
            _771 <= _101;
        42:
            _771 <= _102;
        43:
            _771 <= _103;
        44:
            _771 <= _104;
        45:
            _771 <= _105;
        46:
            _771 <= _106;
        47:
            _771 <= _107;
        48:
            _771 <= _108;
        49:
            _771 <= _109;
        50:
            _771 <= _110;
        51:
            _771 <= _111;
        52:
            _771 <= _112;
        53:
            _771 <= _113;
        54:
            _771 <= _114;
        55:
            _771 <= _115;
        56:
            _771 <= _116;
        57:
            _771 <= _117;
        58:
            _771 <= _118;
        59:
            _771 <= _119;
        60:
            _771 <= _120;
        61:
            _771 <= _121;
        62:
            _771 <= _122;
        63:
            _771 <= _123;
        64:
            _771 <= _124;
        65:
            _771 <= _125;
        66:
            _771 <= _126;
        67:
            _771 <= _127;
        68:
            _771 <= _128;
        69:
            _771 <= _129;
        70:
            _771 <= _130;
        71:
            _771 <= _131;
        72:
            _771 <= _132;
        73:
            _771 <= _133;
        74:
            _771 <= _134;
        75:
            _771 <= _135;
        76:
            _771 <= _136;
        77:
            _771 <= _137;
        78:
            _771 <= _138;
        79:
            _771 <= _139;
        80:
            _771 <= _140;
        81:
            _771 <= _141;
        82:
            _771 <= _142;
        83:
            _771 <= _143;
        84:
            _771 <= _144;
        85:
            _771 <= _145;
        86:
            _771 <= _146;
        87:
            _771 <= _147;
        88:
            _771 <= _148;
        89:
            _771 <= _149;
        90:
            _771 <= _150;
        91:
            _771 <= _151;
        92:
            _771 <= _152;
        93:
            _771 <= _153;
        94:
            _771 <= _154;
        95:
            _771 <= _155;
        96:
            _771 <= _156;
        97:
            _771 <= _157;
        98:
            _771 <= _158;
        99:
            _771 <= _159;
        100:
            _771 <= _160;
        101:
            _771 <= _161;
        102:
            _771 <= _162;
        103:
            _771 <= _163;
        104:
            _771 <= _164;
        105:
            _771 <= _165;
        106:
            _771 <= _166;
        107:
            _771 <= _167;
        108:
            _771 <= _168;
        109:
            _771 <= _169;
        110:
            _771 <= _170;
        111:
            _771 <= _171;
        112:
            _771 <= _172;
        113:
            _771 <= _173;
        114:
            _771 <= _174;
        115:
            _771 <= _175;
        116:
            _771 <= _176;
        117:
            _771 <= _177;
        118:
            _771 <= _178;
        119:
            _771 <= _179;
        120:
            _771 <= _180;
        121:
            _771 <= _181;
        122:
            _771 <= _182;
        123:
            _771 <= _183;
        124:
            _771 <= _184;
        125:
            _771 <= _185;
        126:
            _771 <= _186;
        default:
            _771 <= _187;
        endcase
    end
    assign _767 = _619 < _25;
    assign _772 = _767 ? _771 : _50;
    assign _773 = _40 ? _772 : _321;
    assign _776 = _48 ? _775 : _773;
    assign _6 = _776;
    always @(posedge _22) begin
        if (_20)
            _321 <= _50;
        else
            _321 <= _6;
    end
    assign _965 = { _985,
                    _321 };
    assign _962 = _960 * _982;
    assign _963 = _962[63:0];
    assign _966 = _963 + _965;
    assign _703 = _700 ? _697 : _695;
    assign _706 = _703 < _705;
    assign _707 = ~ _706;
    assign _622 = 4'b0111;
    assign _623 = _622 < _213;
    assign _701 = _626 ? _700 : _42;
    assign _702 = _701 & _623;
    assign _708 = _702 & _707;
    assign _785 = _708 ? _703 : _705;
    assign _573 = _570 ? _567 : _565;
    assign _576 = _573 < _575;
    assign _577 = ~ _576;
    assign _493 = _622 < _213;
    assign _571 = _496 ? _570 : _42;
    assign _572 = _571 & _493;
    assign _578 = _572 & _577;
    assign _704 = _578 ? _573 : _575;
    assign _443 = _440 ? _437 : _435;
    assign _446 = _443 < _445;
    assign _447 = ~ _446;
    assign _363 = _622 < _213;
    assign _441 = _366 ? _440 : _42;
    assign _442 = _441 & _363;
    assign _448 = _442 & _447;
    assign _574 = _448 ? _443 : _445;
    assign _309 = _306 ? _303 : _300;
    assign _313 = _309 < _312;
    assign _314 = ~ _313;
    assign _223 = _622 < _213;
    assign _307 = _226 ? _306 : _42;
    assign _308 = _307 & _223;
    assign _315 = _308 & _314;
    assign _444 = _315 ? _309 : _312;
    assign _445 = _209 ? _444 : _312;
    assign _575 = _205 ? _574 : _445;
    assign _705 = _201 ? _704 : _575;
    assign _786 = _197 ? _785 : _705;
    assign _780 = 8'b00000111;
    assign _781 = _57 + _780;
    always @* begin
        case (_781)
        0:
            _782 <= _60;
        1:
            _782 <= _61;
        2:
            _782 <= _62;
        3:
            _782 <= _63;
        4:
            _782 <= _64;
        5:
            _782 <= _65;
        6:
            _782 <= _66;
        7:
            _782 <= _67;
        8:
            _782 <= _68;
        9:
            _782 <= _69;
        10:
            _782 <= _70;
        11:
            _782 <= _71;
        12:
            _782 <= _72;
        13:
            _782 <= _73;
        14:
            _782 <= _74;
        15:
            _782 <= _75;
        16:
            _782 <= _76;
        17:
            _782 <= _77;
        18:
            _782 <= _78;
        19:
            _782 <= _79;
        20:
            _782 <= _80;
        21:
            _782 <= _81;
        22:
            _782 <= _82;
        23:
            _782 <= _83;
        24:
            _782 <= _84;
        25:
            _782 <= _85;
        26:
            _782 <= _86;
        27:
            _782 <= _87;
        28:
            _782 <= _88;
        29:
            _782 <= _89;
        30:
            _782 <= _90;
        31:
            _782 <= _91;
        32:
            _782 <= _92;
        33:
            _782 <= _93;
        34:
            _782 <= _94;
        35:
            _782 <= _95;
        36:
            _782 <= _96;
        37:
            _782 <= _97;
        38:
            _782 <= _98;
        39:
            _782 <= _99;
        40:
            _782 <= _100;
        41:
            _782 <= _101;
        42:
            _782 <= _102;
        43:
            _782 <= _103;
        44:
            _782 <= _104;
        45:
            _782 <= _105;
        46:
            _782 <= _106;
        47:
            _782 <= _107;
        48:
            _782 <= _108;
        49:
            _782 <= _109;
        50:
            _782 <= _110;
        51:
            _782 <= _111;
        52:
            _782 <= _112;
        53:
            _782 <= _113;
        54:
            _782 <= _114;
        55:
            _782 <= _115;
        56:
            _782 <= _116;
        57:
            _782 <= _117;
        58:
            _782 <= _118;
        59:
            _782 <= _119;
        60:
            _782 <= _120;
        61:
            _782 <= _121;
        62:
            _782 <= _122;
        63:
            _782 <= _123;
        64:
            _782 <= _124;
        65:
            _782 <= _125;
        66:
            _782 <= _126;
        67:
            _782 <= _127;
        68:
            _782 <= _128;
        69:
            _782 <= _129;
        70:
            _782 <= _130;
        71:
            _782 <= _131;
        72:
            _782 <= _132;
        73:
            _782 <= _133;
        74:
            _782 <= _134;
        75:
            _782 <= _135;
        76:
            _782 <= _136;
        77:
            _782 <= _137;
        78:
            _782 <= _138;
        79:
            _782 <= _139;
        80:
            _782 <= _140;
        81:
            _782 <= _141;
        82:
            _782 <= _142;
        83:
            _782 <= _143;
        84:
            _782 <= _144;
        85:
            _782 <= _145;
        86:
            _782 <= _146;
        87:
            _782 <= _147;
        88:
            _782 <= _148;
        89:
            _782 <= _149;
        90:
            _782 <= _150;
        91:
            _782 <= _151;
        92:
            _782 <= _152;
        93:
            _782 <= _153;
        94:
            _782 <= _154;
        95:
            _782 <= _155;
        96:
            _782 <= _156;
        97:
            _782 <= _157;
        98:
            _782 <= _158;
        99:
            _782 <= _159;
        100:
            _782 <= _160;
        101:
            _782 <= _161;
        102:
            _782 <= _162;
        103:
            _782 <= _163;
        104:
            _782 <= _164;
        105:
            _782 <= _165;
        106:
            _782 <= _166;
        107:
            _782 <= _167;
        108:
            _782 <= _168;
        109:
            _782 <= _169;
        110:
            _782 <= _170;
        111:
            _782 <= _171;
        112:
            _782 <= _172;
        113:
            _782 <= _173;
        114:
            _782 <= _174;
        115:
            _782 <= _175;
        116:
            _782 <= _176;
        117:
            _782 <= _177;
        118:
            _782 <= _178;
        119:
            _782 <= _179;
        120:
            _782 <= _180;
        121:
            _782 <= _181;
        122:
            _782 <= _182;
        123:
            _782 <= _183;
        124:
            _782 <= _184;
        125:
            _782 <= _185;
        126:
            _782 <= _186;
        default:
            _782 <= _187;
        endcase
    end
    assign _778 = _622 < _25;
    assign _783 = _778 ? _782 : _50;
    assign _784 = _40 ? _783 : _312;
    assign _787 = _48 ? _786 : _784;
    assign _7 = _787;
    always @(posedge _22) begin
        if (_20)
            _312 <= _50;
        else
            _312 <= _7;
    end
    assign _958 = { _985,
                    _312 };
    assign _955 = _953 * _982;
    assign _956 = _955[63:0];
    assign _959 = _956 + _958;
    assign _695 = _692 ? _689 : _687;
    assign _698 = _695 < _697;
    assign _699 = ~ _698;
    assign _625 = 4'b0110;
    assign _626 = _625 < _213;
    assign _693 = _629 ? _692 : _42;
    assign _694 = _693 & _626;
    assign _700 = _694 & _699;
    assign _796 = _700 ? _695 : _697;
    assign _565 = _562 ? _559 : _557;
    assign _568 = _565 < _567;
    assign _569 = ~ _568;
    assign _496 = _625 < _213;
    assign _563 = _499 ? _562 : _42;
    assign _564 = _563 & _496;
    assign _570 = _564 & _569;
    assign _696 = _570 ? _565 : _567;
    assign _435 = _432 ? _429 : _427;
    assign _438 = _435 < _437;
    assign _439 = ~ _438;
    assign _366 = _625 < _213;
    assign _433 = _369 ? _432 : _42;
    assign _434 = _433 & _366;
    assign _440 = _434 & _439;
    assign _566 = _440 ? _435 : _437;
    assign _300 = _297 ? _294 : _291;
    assign _304 = _300 < _303;
    assign _305 = ~ _304;
    assign _226 = _625 < _213;
    assign _298 = _229 ? _297 : _42;
    assign _299 = _298 & _226;
    assign _306 = _299 & _305;
    assign _436 = _306 ? _300 : _303;
    assign _437 = _209 ? _436 : _303;
    assign _567 = _205 ? _566 : _437;
    assign _697 = _201 ? _696 : _567;
    assign _797 = _197 ? _796 : _697;
    assign _791 = 8'b00000110;
    assign _792 = _57 + _791;
    always @* begin
        case (_792)
        0:
            _793 <= _60;
        1:
            _793 <= _61;
        2:
            _793 <= _62;
        3:
            _793 <= _63;
        4:
            _793 <= _64;
        5:
            _793 <= _65;
        6:
            _793 <= _66;
        7:
            _793 <= _67;
        8:
            _793 <= _68;
        9:
            _793 <= _69;
        10:
            _793 <= _70;
        11:
            _793 <= _71;
        12:
            _793 <= _72;
        13:
            _793 <= _73;
        14:
            _793 <= _74;
        15:
            _793 <= _75;
        16:
            _793 <= _76;
        17:
            _793 <= _77;
        18:
            _793 <= _78;
        19:
            _793 <= _79;
        20:
            _793 <= _80;
        21:
            _793 <= _81;
        22:
            _793 <= _82;
        23:
            _793 <= _83;
        24:
            _793 <= _84;
        25:
            _793 <= _85;
        26:
            _793 <= _86;
        27:
            _793 <= _87;
        28:
            _793 <= _88;
        29:
            _793 <= _89;
        30:
            _793 <= _90;
        31:
            _793 <= _91;
        32:
            _793 <= _92;
        33:
            _793 <= _93;
        34:
            _793 <= _94;
        35:
            _793 <= _95;
        36:
            _793 <= _96;
        37:
            _793 <= _97;
        38:
            _793 <= _98;
        39:
            _793 <= _99;
        40:
            _793 <= _100;
        41:
            _793 <= _101;
        42:
            _793 <= _102;
        43:
            _793 <= _103;
        44:
            _793 <= _104;
        45:
            _793 <= _105;
        46:
            _793 <= _106;
        47:
            _793 <= _107;
        48:
            _793 <= _108;
        49:
            _793 <= _109;
        50:
            _793 <= _110;
        51:
            _793 <= _111;
        52:
            _793 <= _112;
        53:
            _793 <= _113;
        54:
            _793 <= _114;
        55:
            _793 <= _115;
        56:
            _793 <= _116;
        57:
            _793 <= _117;
        58:
            _793 <= _118;
        59:
            _793 <= _119;
        60:
            _793 <= _120;
        61:
            _793 <= _121;
        62:
            _793 <= _122;
        63:
            _793 <= _123;
        64:
            _793 <= _124;
        65:
            _793 <= _125;
        66:
            _793 <= _126;
        67:
            _793 <= _127;
        68:
            _793 <= _128;
        69:
            _793 <= _129;
        70:
            _793 <= _130;
        71:
            _793 <= _131;
        72:
            _793 <= _132;
        73:
            _793 <= _133;
        74:
            _793 <= _134;
        75:
            _793 <= _135;
        76:
            _793 <= _136;
        77:
            _793 <= _137;
        78:
            _793 <= _138;
        79:
            _793 <= _139;
        80:
            _793 <= _140;
        81:
            _793 <= _141;
        82:
            _793 <= _142;
        83:
            _793 <= _143;
        84:
            _793 <= _144;
        85:
            _793 <= _145;
        86:
            _793 <= _146;
        87:
            _793 <= _147;
        88:
            _793 <= _148;
        89:
            _793 <= _149;
        90:
            _793 <= _150;
        91:
            _793 <= _151;
        92:
            _793 <= _152;
        93:
            _793 <= _153;
        94:
            _793 <= _154;
        95:
            _793 <= _155;
        96:
            _793 <= _156;
        97:
            _793 <= _157;
        98:
            _793 <= _158;
        99:
            _793 <= _159;
        100:
            _793 <= _160;
        101:
            _793 <= _161;
        102:
            _793 <= _162;
        103:
            _793 <= _163;
        104:
            _793 <= _164;
        105:
            _793 <= _165;
        106:
            _793 <= _166;
        107:
            _793 <= _167;
        108:
            _793 <= _168;
        109:
            _793 <= _169;
        110:
            _793 <= _170;
        111:
            _793 <= _171;
        112:
            _793 <= _172;
        113:
            _793 <= _173;
        114:
            _793 <= _174;
        115:
            _793 <= _175;
        116:
            _793 <= _176;
        117:
            _793 <= _177;
        118:
            _793 <= _178;
        119:
            _793 <= _179;
        120:
            _793 <= _180;
        121:
            _793 <= _181;
        122:
            _793 <= _182;
        123:
            _793 <= _183;
        124:
            _793 <= _184;
        125:
            _793 <= _185;
        126:
            _793 <= _186;
        default:
            _793 <= _187;
        endcase
    end
    assign _789 = _625 < _25;
    assign _794 = _789 ? _793 : _50;
    assign _795 = _40 ? _794 : _303;
    assign _798 = _48 ? _797 : _795;
    assign _8 = _798;
    always @(posedge _22) begin
        if (_20)
            _303 <= _50;
        else
            _303 <= _8;
    end
    assign _951 = { _985,
                    _303 };
    assign _948 = _946 * _982;
    assign _949 = _948[63:0];
    assign _952 = _949 + _951;
    assign _687 = _684 ? _681 : _679;
    assign _690 = _687 < _689;
    assign _691 = ~ _690;
    assign _628 = 4'b0101;
    assign _629 = _628 < _213;
    assign _685 = _632 ? _684 : _42;
    assign _686 = _685 & _629;
    assign _692 = _686 & _691;
    assign _807 = _692 ? _687 : _689;
    assign _557 = _554 ? _551 : _549;
    assign _560 = _557 < _559;
    assign _561 = ~ _560;
    assign _499 = _628 < _213;
    assign _555 = _502 ? _554 : _42;
    assign _556 = _555 & _499;
    assign _562 = _556 & _561;
    assign _688 = _562 ? _557 : _559;
    assign _427 = _424 ? _421 : _419;
    assign _430 = _427 < _429;
    assign _431 = ~ _430;
    assign _369 = _628 < _213;
    assign _425 = _372 ? _424 : _42;
    assign _426 = _425 & _369;
    assign _432 = _426 & _431;
    assign _558 = _432 ? _427 : _429;
    assign _291 = _288 ? _285 : _282;
    assign _295 = _291 < _294;
    assign _296 = ~ _295;
    assign _229 = _628 < _213;
    assign _289 = _232 ? _288 : _42;
    assign _290 = _289 & _229;
    assign _297 = _290 & _296;
    assign _428 = _297 ? _291 : _294;
    assign _429 = _209 ? _428 : _294;
    assign _559 = _205 ? _558 : _429;
    assign _689 = _201 ? _688 : _559;
    assign _808 = _197 ? _807 : _689;
    assign _802 = 8'b00000101;
    assign _803 = _57 + _802;
    always @* begin
        case (_803)
        0:
            _804 <= _60;
        1:
            _804 <= _61;
        2:
            _804 <= _62;
        3:
            _804 <= _63;
        4:
            _804 <= _64;
        5:
            _804 <= _65;
        6:
            _804 <= _66;
        7:
            _804 <= _67;
        8:
            _804 <= _68;
        9:
            _804 <= _69;
        10:
            _804 <= _70;
        11:
            _804 <= _71;
        12:
            _804 <= _72;
        13:
            _804 <= _73;
        14:
            _804 <= _74;
        15:
            _804 <= _75;
        16:
            _804 <= _76;
        17:
            _804 <= _77;
        18:
            _804 <= _78;
        19:
            _804 <= _79;
        20:
            _804 <= _80;
        21:
            _804 <= _81;
        22:
            _804 <= _82;
        23:
            _804 <= _83;
        24:
            _804 <= _84;
        25:
            _804 <= _85;
        26:
            _804 <= _86;
        27:
            _804 <= _87;
        28:
            _804 <= _88;
        29:
            _804 <= _89;
        30:
            _804 <= _90;
        31:
            _804 <= _91;
        32:
            _804 <= _92;
        33:
            _804 <= _93;
        34:
            _804 <= _94;
        35:
            _804 <= _95;
        36:
            _804 <= _96;
        37:
            _804 <= _97;
        38:
            _804 <= _98;
        39:
            _804 <= _99;
        40:
            _804 <= _100;
        41:
            _804 <= _101;
        42:
            _804 <= _102;
        43:
            _804 <= _103;
        44:
            _804 <= _104;
        45:
            _804 <= _105;
        46:
            _804 <= _106;
        47:
            _804 <= _107;
        48:
            _804 <= _108;
        49:
            _804 <= _109;
        50:
            _804 <= _110;
        51:
            _804 <= _111;
        52:
            _804 <= _112;
        53:
            _804 <= _113;
        54:
            _804 <= _114;
        55:
            _804 <= _115;
        56:
            _804 <= _116;
        57:
            _804 <= _117;
        58:
            _804 <= _118;
        59:
            _804 <= _119;
        60:
            _804 <= _120;
        61:
            _804 <= _121;
        62:
            _804 <= _122;
        63:
            _804 <= _123;
        64:
            _804 <= _124;
        65:
            _804 <= _125;
        66:
            _804 <= _126;
        67:
            _804 <= _127;
        68:
            _804 <= _128;
        69:
            _804 <= _129;
        70:
            _804 <= _130;
        71:
            _804 <= _131;
        72:
            _804 <= _132;
        73:
            _804 <= _133;
        74:
            _804 <= _134;
        75:
            _804 <= _135;
        76:
            _804 <= _136;
        77:
            _804 <= _137;
        78:
            _804 <= _138;
        79:
            _804 <= _139;
        80:
            _804 <= _140;
        81:
            _804 <= _141;
        82:
            _804 <= _142;
        83:
            _804 <= _143;
        84:
            _804 <= _144;
        85:
            _804 <= _145;
        86:
            _804 <= _146;
        87:
            _804 <= _147;
        88:
            _804 <= _148;
        89:
            _804 <= _149;
        90:
            _804 <= _150;
        91:
            _804 <= _151;
        92:
            _804 <= _152;
        93:
            _804 <= _153;
        94:
            _804 <= _154;
        95:
            _804 <= _155;
        96:
            _804 <= _156;
        97:
            _804 <= _157;
        98:
            _804 <= _158;
        99:
            _804 <= _159;
        100:
            _804 <= _160;
        101:
            _804 <= _161;
        102:
            _804 <= _162;
        103:
            _804 <= _163;
        104:
            _804 <= _164;
        105:
            _804 <= _165;
        106:
            _804 <= _166;
        107:
            _804 <= _167;
        108:
            _804 <= _168;
        109:
            _804 <= _169;
        110:
            _804 <= _170;
        111:
            _804 <= _171;
        112:
            _804 <= _172;
        113:
            _804 <= _173;
        114:
            _804 <= _174;
        115:
            _804 <= _175;
        116:
            _804 <= _176;
        117:
            _804 <= _177;
        118:
            _804 <= _178;
        119:
            _804 <= _179;
        120:
            _804 <= _180;
        121:
            _804 <= _181;
        122:
            _804 <= _182;
        123:
            _804 <= _183;
        124:
            _804 <= _184;
        125:
            _804 <= _185;
        126:
            _804 <= _186;
        default:
            _804 <= _187;
        endcase
    end
    assign _800 = _628 < _25;
    assign _805 = _800 ? _804 : _50;
    assign _806 = _40 ? _805 : _294;
    assign _809 = _48 ? _808 : _806;
    assign _9 = _809;
    always @(posedge _22) begin
        if (_20)
            _294 <= _50;
        else
            _294 <= _9;
    end
    assign _944 = { _985,
                    _294 };
    assign _941 = _939 * _982;
    assign _942 = _941[63:0];
    assign _945 = _942 + _944;
    assign _679 = _676 ? _673 : _671;
    assign _682 = _679 < _681;
    assign _683 = ~ _682;
    assign _631 = 4'b0100;
    assign _632 = _631 < _213;
    assign _677 = _635 ? _676 : _42;
    assign _678 = _677 & _632;
    assign _684 = _678 & _683;
    assign _818 = _684 ? _679 : _681;
    assign _549 = _546 ? _543 : _541;
    assign _552 = _549 < _551;
    assign _553 = ~ _552;
    assign _502 = _631 < _213;
    assign _547 = _505 ? _546 : _42;
    assign _548 = _547 & _502;
    assign _554 = _548 & _553;
    assign _680 = _554 ? _549 : _551;
    assign _419 = _416 ? _413 : _411;
    assign _422 = _419 < _421;
    assign _423 = ~ _422;
    assign _372 = _631 < _213;
    assign _417 = _375 ? _416 : _42;
    assign _418 = _417 & _372;
    assign _424 = _418 & _423;
    assign _550 = _424 ? _419 : _421;
    assign _282 = _279 ? _276 : _273;
    assign _286 = _282 < _285;
    assign _287 = ~ _286;
    assign _232 = _631 < _213;
    assign _280 = _235 ? _279 : _42;
    assign _281 = _280 & _232;
    assign _288 = _281 & _287;
    assign _420 = _288 ? _282 : _285;
    assign _421 = _209 ? _420 : _285;
    assign _551 = _205 ? _550 : _421;
    assign _681 = _201 ? _680 : _551;
    assign _819 = _197 ? _818 : _681;
    assign _813 = 8'b00000100;
    assign _814 = _57 + _813;
    always @* begin
        case (_814)
        0:
            _815 <= _60;
        1:
            _815 <= _61;
        2:
            _815 <= _62;
        3:
            _815 <= _63;
        4:
            _815 <= _64;
        5:
            _815 <= _65;
        6:
            _815 <= _66;
        7:
            _815 <= _67;
        8:
            _815 <= _68;
        9:
            _815 <= _69;
        10:
            _815 <= _70;
        11:
            _815 <= _71;
        12:
            _815 <= _72;
        13:
            _815 <= _73;
        14:
            _815 <= _74;
        15:
            _815 <= _75;
        16:
            _815 <= _76;
        17:
            _815 <= _77;
        18:
            _815 <= _78;
        19:
            _815 <= _79;
        20:
            _815 <= _80;
        21:
            _815 <= _81;
        22:
            _815 <= _82;
        23:
            _815 <= _83;
        24:
            _815 <= _84;
        25:
            _815 <= _85;
        26:
            _815 <= _86;
        27:
            _815 <= _87;
        28:
            _815 <= _88;
        29:
            _815 <= _89;
        30:
            _815 <= _90;
        31:
            _815 <= _91;
        32:
            _815 <= _92;
        33:
            _815 <= _93;
        34:
            _815 <= _94;
        35:
            _815 <= _95;
        36:
            _815 <= _96;
        37:
            _815 <= _97;
        38:
            _815 <= _98;
        39:
            _815 <= _99;
        40:
            _815 <= _100;
        41:
            _815 <= _101;
        42:
            _815 <= _102;
        43:
            _815 <= _103;
        44:
            _815 <= _104;
        45:
            _815 <= _105;
        46:
            _815 <= _106;
        47:
            _815 <= _107;
        48:
            _815 <= _108;
        49:
            _815 <= _109;
        50:
            _815 <= _110;
        51:
            _815 <= _111;
        52:
            _815 <= _112;
        53:
            _815 <= _113;
        54:
            _815 <= _114;
        55:
            _815 <= _115;
        56:
            _815 <= _116;
        57:
            _815 <= _117;
        58:
            _815 <= _118;
        59:
            _815 <= _119;
        60:
            _815 <= _120;
        61:
            _815 <= _121;
        62:
            _815 <= _122;
        63:
            _815 <= _123;
        64:
            _815 <= _124;
        65:
            _815 <= _125;
        66:
            _815 <= _126;
        67:
            _815 <= _127;
        68:
            _815 <= _128;
        69:
            _815 <= _129;
        70:
            _815 <= _130;
        71:
            _815 <= _131;
        72:
            _815 <= _132;
        73:
            _815 <= _133;
        74:
            _815 <= _134;
        75:
            _815 <= _135;
        76:
            _815 <= _136;
        77:
            _815 <= _137;
        78:
            _815 <= _138;
        79:
            _815 <= _139;
        80:
            _815 <= _140;
        81:
            _815 <= _141;
        82:
            _815 <= _142;
        83:
            _815 <= _143;
        84:
            _815 <= _144;
        85:
            _815 <= _145;
        86:
            _815 <= _146;
        87:
            _815 <= _147;
        88:
            _815 <= _148;
        89:
            _815 <= _149;
        90:
            _815 <= _150;
        91:
            _815 <= _151;
        92:
            _815 <= _152;
        93:
            _815 <= _153;
        94:
            _815 <= _154;
        95:
            _815 <= _155;
        96:
            _815 <= _156;
        97:
            _815 <= _157;
        98:
            _815 <= _158;
        99:
            _815 <= _159;
        100:
            _815 <= _160;
        101:
            _815 <= _161;
        102:
            _815 <= _162;
        103:
            _815 <= _163;
        104:
            _815 <= _164;
        105:
            _815 <= _165;
        106:
            _815 <= _166;
        107:
            _815 <= _167;
        108:
            _815 <= _168;
        109:
            _815 <= _169;
        110:
            _815 <= _170;
        111:
            _815 <= _171;
        112:
            _815 <= _172;
        113:
            _815 <= _173;
        114:
            _815 <= _174;
        115:
            _815 <= _175;
        116:
            _815 <= _176;
        117:
            _815 <= _177;
        118:
            _815 <= _178;
        119:
            _815 <= _179;
        120:
            _815 <= _180;
        121:
            _815 <= _181;
        122:
            _815 <= _182;
        123:
            _815 <= _183;
        124:
            _815 <= _184;
        125:
            _815 <= _185;
        126:
            _815 <= _186;
        default:
            _815 <= _187;
        endcase
    end
    assign _811 = _631 < _25;
    assign _816 = _811 ? _815 : _50;
    assign _817 = _40 ? _816 : _285;
    assign _820 = _48 ? _819 : _817;
    assign _10 = _820;
    always @(posedge _22) begin
        if (_20)
            _285 <= _50;
        else
            _285 <= _10;
    end
    assign _937 = { _985,
                    _285 };
    assign _934 = _932 * _982;
    assign _935 = _934[63:0];
    assign _938 = _935 + _937;
    assign _671 = _668 ? _665 : _663;
    assign _674 = _671 < _673;
    assign _675 = ~ _674;
    assign _634 = 4'b0011;
    assign _635 = _634 < _213;
    assign _669 = _638 ? _668 : _42;
    assign _670 = _669 & _635;
    assign _676 = _670 & _675;
    assign _829 = _676 ? _671 : _673;
    assign _541 = _538 ? _535 : _533;
    assign _544 = _541 < _543;
    assign _545 = ~ _544;
    assign _505 = _634 < _213;
    assign _539 = _508 ? _538 : _42;
    assign _540 = _539 & _505;
    assign _546 = _540 & _545;
    assign _672 = _546 ? _541 : _543;
    assign _411 = _408 ? _405 : _403;
    assign _414 = _411 < _413;
    assign _415 = ~ _414;
    assign _375 = _634 < _213;
    assign _409 = _378 ? _408 : _42;
    assign _410 = _409 & _375;
    assign _416 = _410 & _415;
    assign _542 = _416 ? _411 : _413;
    assign _273 = _270 ? _267 : _264;
    assign _277 = _273 < _276;
    assign _278 = ~ _277;
    assign _235 = _634 < _213;
    assign _271 = _238 ? _270 : _42;
    assign _272 = _271 & _235;
    assign _279 = _272 & _278;
    assign _412 = _279 ? _273 : _276;
    assign _413 = _209 ? _412 : _276;
    assign _543 = _205 ? _542 : _413;
    assign _673 = _201 ? _672 : _543;
    assign _830 = _197 ? _829 : _673;
    assign _824 = 8'b00000011;
    assign _825 = _57 + _824;
    always @* begin
        case (_825)
        0:
            _826 <= _60;
        1:
            _826 <= _61;
        2:
            _826 <= _62;
        3:
            _826 <= _63;
        4:
            _826 <= _64;
        5:
            _826 <= _65;
        6:
            _826 <= _66;
        7:
            _826 <= _67;
        8:
            _826 <= _68;
        9:
            _826 <= _69;
        10:
            _826 <= _70;
        11:
            _826 <= _71;
        12:
            _826 <= _72;
        13:
            _826 <= _73;
        14:
            _826 <= _74;
        15:
            _826 <= _75;
        16:
            _826 <= _76;
        17:
            _826 <= _77;
        18:
            _826 <= _78;
        19:
            _826 <= _79;
        20:
            _826 <= _80;
        21:
            _826 <= _81;
        22:
            _826 <= _82;
        23:
            _826 <= _83;
        24:
            _826 <= _84;
        25:
            _826 <= _85;
        26:
            _826 <= _86;
        27:
            _826 <= _87;
        28:
            _826 <= _88;
        29:
            _826 <= _89;
        30:
            _826 <= _90;
        31:
            _826 <= _91;
        32:
            _826 <= _92;
        33:
            _826 <= _93;
        34:
            _826 <= _94;
        35:
            _826 <= _95;
        36:
            _826 <= _96;
        37:
            _826 <= _97;
        38:
            _826 <= _98;
        39:
            _826 <= _99;
        40:
            _826 <= _100;
        41:
            _826 <= _101;
        42:
            _826 <= _102;
        43:
            _826 <= _103;
        44:
            _826 <= _104;
        45:
            _826 <= _105;
        46:
            _826 <= _106;
        47:
            _826 <= _107;
        48:
            _826 <= _108;
        49:
            _826 <= _109;
        50:
            _826 <= _110;
        51:
            _826 <= _111;
        52:
            _826 <= _112;
        53:
            _826 <= _113;
        54:
            _826 <= _114;
        55:
            _826 <= _115;
        56:
            _826 <= _116;
        57:
            _826 <= _117;
        58:
            _826 <= _118;
        59:
            _826 <= _119;
        60:
            _826 <= _120;
        61:
            _826 <= _121;
        62:
            _826 <= _122;
        63:
            _826 <= _123;
        64:
            _826 <= _124;
        65:
            _826 <= _125;
        66:
            _826 <= _126;
        67:
            _826 <= _127;
        68:
            _826 <= _128;
        69:
            _826 <= _129;
        70:
            _826 <= _130;
        71:
            _826 <= _131;
        72:
            _826 <= _132;
        73:
            _826 <= _133;
        74:
            _826 <= _134;
        75:
            _826 <= _135;
        76:
            _826 <= _136;
        77:
            _826 <= _137;
        78:
            _826 <= _138;
        79:
            _826 <= _139;
        80:
            _826 <= _140;
        81:
            _826 <= _141;
        82:
            _826 <= _142;
        83:
            _826 <= _143;
        84:
            _826 <= _144;
        85:
            _826 <= _145;
        86:
            _826 <= _146;
        87:
            _826 <= _147;
        88:
            _826 <= _148;
        89:
            _826 <= _149;
        90:
            _826 <= _150;
        91:
            _826 <= _151;
        92:
            _826 <= _152;
        93:
            _826 <= _153;
        94:
            _826 <= _154;
        95:
            _826 <= _155;
        96:
            _826 <= _156;
        97:
            _826 <= _157;
        98:
            _826 <= _158;
        99:
            _826 <= _159;
        100:
            _826 <= _160;
        101:
            _826 <= _161;
        102:
            _826 <= _162;
        103:
            _826 <= _163;
        104:
            _826 <= _164;
        105:
            _826 <= _165;
        106:
            _826 <= _166;
        107:
            _826 <= _167;
        108:
            _826 <= _168;
        109:
            _826 <= _169;
        110:
            _826 <= _170;
        111:
            _826 <= _171;
        112:
            _826 <= _172;
        113:
            _826 <= _173;
        114:
            _826 <= _174;
        115:
            _826 <= _175;
        116:
            _826 <= _176;
        117:
            _826 <= _177;
        118:
            _826 <= _178;
        119:
            _826 <= _179;
        120:
            _826 <= _180;
        121:
            _826 <= _181;
        122:
            _826 <= _182;
        123:
            _826 <= _183;
        124:
            _826 <= _184;
        125:
            _826 <= _185;
        126:
            _826 <= _186;
        default:
            _826 <= _187;
        endcase
    end
    assign _822 = _634 < _25;
    assign _827 = _822 ? _826 : _50;
    assign _828 = _40 ? _827 : _276;
    assign _831 = _48 ? _830 : _828;
    assign _11 = _831;
    always @(posedge _22) begin
        if (_20)
            _276 <= _50;
        else
            _276 <= _11;
    end
    assign _930 = { _985,
                    _276 };
    assign _927 = _925 * _982;
    assign _928 = _927[63:0];
    assign _931 = _928 + _930;
    assign _663 = _660 ? _657 : _655;
    assign _666 = _663 < _665;
    assign _667 = ~ _666;
    assign _637 = 4'b0010;
    assign _638 = _637 < _213;
    assign _661 = _641 ? _660 : _42;
    assign _662 = _661 & _638;
    assign _668 = _662 & _667;
    assign _840 = _668 ? _663 : _665;
    assign _533 = _530 ? _527 : _525;
    assign _536 = _533 < _535;
    assign _537 = ~ _536;
    assign _508 = _637 < _213;
    assign _531 = _511 ? _530 : _42;
    assign _532 = _531 & _508;
    assign _538 = _532 & _537;
    assign _664 = _538 ? _533 : _535;
    assign _403 = _400 ? _397 : _395;
    assign _406 = _403 < _405;
    assign _407 = ~ _406;
    assign _378 = _637 < _213;
    assign _401 = _381 ? _400 : _42;
    assign _402 = _401 & _378;
    assign _408 = _402 & _407;
    assign _534 = _408 ? _403 : _405;
    assign _264 = _261 ? _258 : _255;
    assign _268 = _264 < _267;
    assign _269 = ~ _268;
    assign _238 = _637 < _213;
    assign _262 = _241 ? _261 : _42;
    assign _263 = _262 & _238;
    assign _270 = _263 & _269;
    assign _404 = _270 ? _264 : _267;
    assign _405 = _209 ? _404 : _267;
    assign _535 = _205 ? _534 : _405;
    assign _665 = _201 ? _664 : _535;
    assign _841 = _197 ? _840 : _665;
    assign _835 = 8'b00000010;
    assign _836 = _57 + _835;
    always @* begin
        case (_836)
        0:
            _837 <= _60;
        1:
            _837 <= _61;
        2:
            _837 <= _62;
        3:
            _837 <= _63;
        4:
            _837 <= _64;
        5:
            _837 <= _65;
        6:
            _837 <= _66;
        7:
            _837 <= _67;
        8:
            _837 <= _68;
        9:
            _837 <= _69;
        10:
            _837 <= _70;
        11:
            _837 <= _71;
        12:
            _837 <= _72;
        13:
            _837 <= _73;
        14:
            _837 <= _74;
        15:
            _837 <= _75;
        16:
            _837 <= _76;
        17:
            _837 <= _77;
        18:
            _837 <= _78;
        19:
            _837 <= _79;
        20:
            _837 <= _80;
        21:
            _837 <= _81;
        22:
            _837 <= _82;
        23:
            _837 <= _83;
        24:
            _837 <= _84;
        25:
            _837 <= _85;
        26:
            _837 <= _86;
        27:
            _837 <= _87;
        28:
            _837 <= _88;
        29:
            _837 <= _89;
        30:
            _837 <= _90;
        31:
            _837 <= _91;
        32:
            _837 <= _92;
        33:
            _837 <= _93;
        34:
            _837 <= _94;
        35:
            _837 <= _95;
        36:
            _837 <= _96;
        37:
            _837 <= _97;
        38:
            _837 <= _98;
        39:
            _837 <= _99;
        40:
            _837 <= _100;
        41:
            _837 <= _101;
        42:
            _837 <= _102;
        43:
            _837 <= _103;
        44:
            _837 <= _104;
        45:
            _837 <= _105;
        46:
            _837 <= _106;
        47:
            _837 <= _107;
        48:
            _837 <= _108;
        49:
            _837 <= _109;
        50:
            _837 <= _110;
        51:
            _837 <= _111;
        52:
            _837 <= _112;
        53:
            _837 <= _113;
        54:
            _837 <= _114;
        55:
            _837 <= _115;
        56:
            _837 <= _116;
        57:
            _837 <= _117;
        58:
            _837 <= _118;
        59:
            _837 <= _119;
        60:
            _837 <= _120;
        61:
            _837 <= _121;
        62:
            _837 <= _122;
        63:
            _837 <= _123;
        64:
            _837 <= _124;
        65:
            _837 <= _125;
        66:
            _837 <= _126;
        67:
            _837 <= _127;
        68:
            _837 <= _128;
        69:
            _837 <= _129;
        70:
            _837 <= _130;
        71:
            _837 <= _131;
        72:
            _837 <= _132;
        73:
            _837 <= _133;
        74:
            _837 <= _134;
        75:
            _837 <= _135;
        76:
            _837 <= _136;
        77:
            _837 <= _137;
        78:
            _837 <= _138;
        79:
            _837 <= _139;
        80:
            _837 <= _140;
        81:
            _837 <= _141;
        82:
            _837 <= _142;
        83:
            _837 <= _143;
        84:
            _837 <= _144;
        85:
            _837 <= _145;
        86:
            _837 <= _146;
        87:
            _837 <= _147;
        88:
            _837 <= _148;
        89:
            _837 <= _149;
        90:
            _837 <= _150;
        91:
            _837 <= _151;
        92:
            _837 <= _152;
        93:
            _837 <= _153;
        94:
            _837 <= _154;
        95:
            _837 <= _155;
        96:
            _837 <= _156;
        97:
            _837 <= _157;
        98:
            _837 <= _158;
        99:
            _837 <= _159;
        100:
            _837 <= _160;
        101:
            _837 <= _161;
        102:
            _837 <= _162;
        103:
            _837 <= _163;
        104:
            _837 <= _164;
        105:
            _837 <= _165;
        106:
            _837 <= _166;
        107:
            _837 <= _167;
        108:
            _837 <= _168;
        109:
            _837 <= _169;
        110:
            _837 <= _170;
        111:
            _837 <= _171;
        112:
            _837 <= _172;
        113:
            _837 <= _173;
        114:
            _837 <= _174;
        115:
            _837 <= _175;
        116:
            _837 <= _176;
        117:
            _837 <= _177;
        118:
            _837 <= _178;
        119:
            _837 <= _179;
        120:
            _837 <= _180;
        121:
            _837 <= _181;
        122:
            _837 <= _182;
        123:
            _837 <= _183;
        124:
            _837 <= _184;
        125:
            _837 <= _185;
        126:
            _837 <= _186;
        default:
            _837 <= _187;
        endcase
    end
    assign _833 = _637 < _25;
    assign _838 = _833 ? _837 : _50;
    assign _839 = _40 ? _838 : _267;
    assign _842 = _48 ? _841 : _839;
    assign _12 = _842;
    always @(posedge _22) begin
        if (_20)
            _267 <= _50;
        else
            _267 <= _12;
    end
    assign _923 = { _985,
                    _267 };
    assign _920 = _918 * _982;
    assign _921 = _920[63:0];
    assign _924 = _921 + _923;
    assign _655 = _652 ? _649 : _647;
    assign _658 = _655 < _657;
    assign _659 = ~ _658;
    assign _640 = 4'b0001;
    assign _641 = _640 < _213;
    assign _653 = _644 ? _652 : _42;
    assign _654 = _653 & _641;
    assign _660 = _654 & _659;
    assign _851 = _660 ? _655 : _657;
    assign _525 = _522 ? _519 : _517;
    assign _528 = _525 < _527;
    assign _529 = ~ _528;
    assign _511 = _640 < _213;
    assign _523 = _514 ? _522 : _42;
    assign _524 = _523 & _511;
    assign _530 = _524 & _529;
    assign _656 = _530 ? _525 : _527;
    assign _395 = _392 ? _389 : _387;
    assign _398 = _395 < _397;
    assign _399 = ~ _398;
    assign _381 = _640 < _213;
    assign _393 = _384 ? _392 : _42;
    assign _394 = _393 & _381;
    assign _400 = _394 & _399;
    assign _526 = _400 ? _395 : _397;
    assign _255 = _252 ? _249 : _246;
    assign _259 = _255 < _258;
    assign _260 = ~ _259;
    assign _241 = _640 < _213;
    assign _253 = _244 ? _252 : _42;
    assign _254 = _253 & _241;
    assign _261 = _254 & _260;
    assign _396 = _261 ? _255 : _258;
    assign _397 = _209 ? _396 : _258;
    assign _527 = _205 ? _526 : _397;
    assign _657 = _201 ? _656 : _527;
    assign _852 = _197 ? _851 : _657;
    assign _846 = 8'b00000001;
    assign _847 = _57 + _846;
    always @* begin
        case (_847)
        0:
            _848 <= _60;
        1:
            _848 <= _61;
        2:
            _848 <= _62;
        3:
            _848 <= _63;
        4:
            _848 <= _64;
        5:
            _848 <= _65;
        6:
            _848 <= _66;
        7:
            _848 <= _67;
        8:
            _848 <= _68;
        9:
            _848 <= _69;
        10:
            _848 <= _70;
        11:
            _848 <= _71;
        12:
            _848 <= _72;
        13:
            _848 <= _73;
        14:
            _848 <= _74;
        15:
            _848 <= _75;
        16:
            _848 <= _76;
        17:
            _848 <= _77;
        18:
            _848 <= _78;
        19:
            _848 <= _79;
        20:
            _848 <= _80;
        21:
            _848 <= _81;
        22:
            _848 <= _82;
        23:
            _848 <= _83;
        24:
            _848 <= _84;
        25:
            _848 <= _85;
        26:
            _848 <= _86;
        27:
            _848 <= _87;
        28:
            _848 <= _88;
        29:
            _848 <= _89;
        30:
            _848 <= _90;
        31:
            _848 <= _91;
        32:
            _848 <= _92;
        33:
            _848 <= _93;
        34:
            _848 <= _94;
        35:
            _848 <= _95;
        36:
            _848 <= _96;
        37:
            _848 <= _97;
        38:
            _848 <= _98;
        39:
            _848 <= _99;
        40:
            _848 <= _100;
        41:
            _848 <= _101;
        42:
            _848 <= _102;
        43:
            _848 <= _103;
        44:
            _848 <= _104;
        45:
            _848 <= _105;
        46:
            _848 <= _106;
        47:
            _848 <= _107;
        48:
            _848 <= _108;
        49:
            _848 <= _109;
        50:
            _848 <= _110;
        51:
            _848 <= _111;
        52:
            _848 <= _112;
        53:
            _848 <= _113;
        54:
            _848 <= _114;
        55:
            _848 <= _115;
        56:
            _848 <= _116;
        57:
            _848 <= _117;
        58:
            _848 <= _118;
        59:
            _848 <= _119;
        60:
            _848 <= _120;
        61:
            _848 <= _121;
        62:
            _848 <= _122;
        63:
            _848 <= _123;
        64:
            _848 <= _124;
        65:
            _848 <= _125;
        66:
            _848 <= _126;
        67:
            _848 <= _127;
        68:
            _848 <= _128;
        69:
            _848 <= _129;
        70:
            _848 <= _130;
        71:
            _848 <= _131;
        72:
            _848 <= _132;
        73:
            _848 <= _133;
        74:
            _848 <= _134;
        75:
            _848 <= _135;
        76:
            _848 <= _136;
        77:
            _848 <= _137;
        78:
            _848 <= _138;
        79:
            _848 <= _139;
        80:
            _848 <= _140;
        81:
            _848 <= _141;
        82:
            _848 <= _142;
        83:
            _848 <= _143;
        84:
            _848 <= _144;
        85:
            _848 <= _145;
        86:
            _848 <= _146;
        87:
            _848 <= _147;
        88:
            _848 <= _148;
        89:
            _848 <= _149;
        90:
            _848 <= _150;
        91:
            _848 <= _151;
        92:
            _848 <= _152;
        93:
            _848 <= _153;
        94:
            _848 <= _154;
        95:
            _848 <= _155;
        96:
            _848 <= _156;
        97:
            _848 <= _157;
        98:
            _848 <= _158;
        99:
            _848 <= _159;
        100:
            _848 <= _160;
        101:
            _848 <= _161;
        102:
            _848 <= _162;
        103:
            _848 <= _163;
        104:
            _848 <= _164;
        105:
            _848 <= _165;
        106:
            _848 <= _166;
        107:
            _848 <= _167;
        108:
            _848 <= _168;
        109:
            _848 <= _169;
        110:
            _848 <= _170;
        111:
            _848 <= _171;
        112:
            _848 <= _172;
        113:
            _848 <= _173;
        114:
            _848 <= _174;
        115:
            _848 <= _175;
        116:
            _848 <= _176;
        117:
            _848 <= _177;
        118:
            _848 <= _178;
        119:
            _848 <= _179;
        120:
            _848 <= _180;
        121:
            _848 <= _181;
        122:
            _848 <= _182;
        123:
            _848 <= _183;
        124:
            _848 <= _184;
        125:
            _848 <= _185;
        126:
            _848 <= _186;
        default:
            _848 <= _187;
        endcase
    end
    assign _844 = _640 < _25;
    assign _849 = _844 ? _848 : _50;
    assign _850 = _40 ? _849 : _258;
    assign _853 = _48 ? _852 : _850;
    assign _13 = _853;
    always @(posedge _22) begin
        if (_20)
            _258 <= _50;
        else
            _258 <= _13;
    end
    assign _916 = { _985,
                    _258 };
    assign _913 = _911 * _982;
    assign _914 = _913[63:0];
    assign _917 = _914 + _916;
    assign _646 = _193 - _824;
    always @* begin
        case (_646)
        0:
            _647 <= _60;
        1:
            _647 <= _61;
        2:
            _647 <= _62;
        3:
            _647 <= _63;
        4:
            _647 <= _64;
        5:
            _647 <= _65;
        6:
            _647 <= _66;
        7:
            _647 <= _67;
        8:
            _647 <= _68;
        9:
            _647 <= _69;
        10:
            _647 <= _70;
        11:
            _647 <= _71;
        12:
            _647 <= _72;
        13:
            _647 <= _73;
        14:
            _647 <= _74;
        15:
            _647 <= _75;
        16:
            _647 <= _76;
        17:
            _647 <= _77;
        18:
            _647 <= _78;
        19:
            _647 <= _79;
        20:
            _647 <= _80;
        21:
            _647 <= _81;
        22:
            _647 <= _82;
        23:
            _647 <= _83;
        24:
            _647 <= _84;
        25:
            _647 <= _85;
        26:
            _647 <= _86;
        27:
            _647 <= _87;
        28:
            _647 <= _88;
        29:
            _647 <= _89;
        30:
            _647 <= _90;
        31:
            _647 <= _91;
        32:
            _647 <= _92;
        33:
            _647 <= _93;
        34:
            _647 <= _94;
        35:
            _647 <= _95;
        36:
            _647 <= _96;
        37:
            _647 <= _97;
        38:
            _647 <= _98;
        39:
            _647 <= _99;
        40:
            _647 <= _100;
        41:
            _647 <= _101;
        42:
            _647 <= _102;
        43:
            _647 <= _103;
        44:
            _647 <= _104;
        45:
            _647 <= _105;
        46:
            _647 <= _106;
        47:
            _647 <= _107;
        48:
            _647 <= _108;
        49:
            _647 <= _109;
        50:
            _647 <= _110;
        51:
            _647 <= _111;
        52:
            _647 <= _112;
        53:
            _647 <= _113;
        54:
            _647 <= _114;
        55:
            _647 <= _115;
        56:
            _647 <= _116;
        57:
            _647 <= _117;
        58:
            _647 <= _118;
        59:
            _647 <= _119;
        60:
            _647 <= _120;
        61:
            _647 <= _121;
        62:
            _647 <= _122;
        63:
            _647 <= _123;
        64:
            _647 <= _124;
        65:
            _647 <= _125;
        66:
            _647 <= _126;
        67:
            _647 <= _127;
        68:
            _647 <= _128;
        69:
            _647 <= _129;
        70:
            _647 <= _130;
        71:
            _647 <= _131;
        72:
            _647 <= _132;
        73:
            _647 <= _133;
        74:
            _647 <= _134;
        75:
            _647 <= _135;
        76:
            _647 <= _136;
        77:
            _647 <= _137;
        78:
            _647 <= _138;
        79:
            _647 <= _139;
        80:
            _647 <= _140;
        81:
            _647 <= _141;
        82:
            _647 <= _142;
        83:
            _647 <= _143;
        84:
            _647 <= _144;
        85:
            _647 <= _145;
        86:
            _647 <= _146;
        87:
            _647 <= _147;
        88:
            _647 <= _148;
        89:
            _647 <= _149;
        90:
            _647 <= _150;
        91:
            _647 <= _151;
        92:
            _647 <= _152;
        93:
            _647 <= _153;
        94:
            _647 <= _154;
        95:
            _647 <= _155;
        96:
            _647 <= _156;
        97:
            _647 <= _157;
        98:
            _647 <= _158;
        99:
            _647 <= _159;
        100:
            _647 <= _160;
        101:
            _647 <= _161;
        102:
            _647 <= _162;
        103:
            _647 <= _163;
        104:
            _647 <= _164;
        105:
            _647 <= _165;
        106:
            _647 <= _166;
        107:
            _647 <= _167;
        108:
            _647 <= _168;
        109:
            _647 <= _169;
        110:
            _647 <= _170;
        111:
            _647 <= _171;
        112:
            _647 <= _172;
        113:
            _647 <= _173;
        114:
            _647 <= _174;
        115:
            _647 <= _175;
        116:
            _647 <= _176;
        117:
            _647 <= _177;
        118:
            _647 <= _178;
        119:
            _647 <= _179;
        120:
            _647 <= _180;
        121:
            _647 <= _181;
        122:
            _647 <= _182;
        123:
            _647 <= _183;
        124:
            _647 <= _184;
        125:
            _647 <= _185;
        126:
            _647 <= _186;
        default:
            _647 <= _187;
        endcase
    end
    assign _650 = _647 < _649;
    assign _651 = ~ _650;
    assign _644 = _50 < _213;
    assign _652 = _644 & _651;
    assign _860 = _652 ? _647 : _649;
    assign _516 = _193 - _835;
    always @* begin
        case (_516)
        0:
            _517 <= _60;
        1:
            _517 <= _61;
        2:
            _517 <= _62;
        3:
            _517 <= _63;
        4:
            _517 <= _64;
        5:
            _517 <= _65;
        6:
            _517 <= _66;
        7:
            _517 <= _67;
        8:
            _517 <= _68;
        9:
            _517 <= _69;
        10:
            _517 <= _70;
        11:
            _517 <= _71;
        12:
            _517 <= _72;
        13:
            _517 <= _73;
        14:
            _517 <= _74;
        15:
            _517 <= _75;
        16:
            _517 <= _76;
        17:
            _517 <= _77;
        18:
            _517 <= _78;
        19:
            _517 <= _79;
        20:
            _517 <= _80;
        21:
            _517 <= _81;
        22:
            _517 <= _82;
        23:
            _517 <= _83;
        24:
            _517 <= _84;
        25:
            _517 <= _85;
        26:
            _517 <= _86;
        27:
            _517 <= _87;
        28:
            _517 <= _88;
        29:
            _517 <= _89;
        30:
            _517 <= _90;
        31:
            _517 <= _91;
        32:
            _517 <= _92;
        33:
            _517 <= _93;
        34:
            _517 <= _94;
        35:
            _517 <= _95;
        36:
            _517 <= _96;
        37:
            _517 <= _97;
        38:
            _517 <= _98;
        39:
            _517 <= _99;
        40:
            _517 <= _100;
        41:
            _517 <= _101;
        42:
            _517 <= _102;
        43:
            _517 <= _103;
        44:
            _517 <= _104;
        45:
            _517 <= _105;
        46:
            _517 <= _106;
        47:
            _517 <= _107;
        48:
            _517 <= _108;
        49:
            _517 <= _109;
        50:
            _517 <= _110;
        51:
            _517 <= _111;
        52:
            _517 <= _112;
        53:
            _517 <= _113;
        54:
            _517 <= _114;
        55:
            _517 <= _115;
        56:
            _517 <= _116;
        57:
            _517 <= _117;
        58:
            _517 <= _118;
        59:
            _517 <= _119;
        60:
            _517 <= _120;
        61:
            _517 <= _121;
        62:
            _517 <= _122;
        63:
            _517 <= _123;
        64:
            _517 <= _124;
        65:
            _517 <= _125;
        66:
            _517 <= _126;
        67:
            _517 <= _127;
        68:
            _517 <= _128;
        69:
            _517 <= _129;
        70:
            _517 <= _130;
        71:
            _517 <= _131;
        72:
            _517 <= _132;
        73:
            _517 <= _133;
        74:
            _517 <= _134;
        75:
            _517 <= _135;
        76:
            _517 <= _136;
        77:
            _517 <= _137;
        78:
            _517 <= _138;
        79:
            _517 <= _139;
        80:
            _517 <= _140;
        81:
            _517 <= _141;
        82:
            _517 <= _142;
        83:
            _517 <= _143;
        84:
            _517 <= _144;
        85:
            _517 <= _145;
        86:
            _517 <= _146;
        87:
            _517 <= _147;
        88:
            _517 <= _148;
        89:
            _517 <= _149;
        90:
            _517 <= _150;
        91:
            _517 <= _151;
        92:
            _517 <= _152;
        93:
            _517 <= _153;
        94:
            _517 <= _154;
        95:
            _517 <= _155;
        96:
            _517 <= _156;
        97:
            _517 <= _157;
        98:
            _517 <= _158;
        99:
            _517 <= _159;
        100:
            _517 <= _160;
        101:
            _517 <= _161;
        102:
            _517 <= _162;
        103:
            _517 <= _163;
        104:
            _517 <= _164;
        105:
            _517 <= _165;
        106:
            _517 <= _166;
        107:
            _517 <= _167;
        108:
            _517 <= _168;
        109:
            _517 <= _169;
        110:
            _517 <= _170;
        111:
            _517 <= _171;
        112:
            _517 <= _172;
        113:
            _517 <= _173;
        114:
            _517 <= _174;
        115:
            _517 <= _175;
        116:
            _517 <= _176;
        117:
            _517 <= _177;
        118:
            _517 <= _178;
        119:
            _517 <= _179;
        120:
            _517 <= _180;
        121:
            _517 <= _181;
        122:
            _517 <= _182;
        123:
            _517 <= _183;
        124:
            _517 <= _184;
        125:
            _517 <= _185;
        126:
            _517 <= _186;
        default:
            _517 <= _187;
        endcase
    end
    assign _520 = _517 < _519;
    assign _521 = ~ _520;
    assign _514 = _50 < _213;
    assign _522 = _514 & _521;
    assign _648 = _522 ? _517 : _519;
    assign _386 = _193 - _846;
    always @* begin
        case (_386)
        0:
            _387 <= _60;
        1:
            _387 <= _61;
        2:
            _387 <= _62;
        3:
            _387 <= _63;
        4:
            _387 <= _64;
        5:
            _387 <= _65;
        6:
            _387 <= _66;
        7:
            _387 <= _67;
        8:
            _387 <= _68;
        9:
            _387 <= _69;
        10:
            _387 <= _70;
        11:
            _387 <= _71;
        12:
            _387 <= _72;
        13:
            _387 <= _73;
        14:
            _387 <= _74;
        15:
            _387 <= _75;
        16:
            _387 <= _76;
        17:
            _387 <= _77;
        18:
            _387 <= _78;
        19:
            _387 <= _79;
        20:
            _387 <= _80;
        21:
            _387 <= _81;
        22:
            _387 <= _82;
        23:
            _387 <= _83;
        24:
            _387 <= _84;
        25:
            _387 <= _85;
        26:
            _387 <= _86;
        27:
            _387 <= _87;
        28:
            _387 <= _88;
        29:
            _387 <= _89;
        30:
            _387 <= _90;
        31:
            _387 <= _91;
        32:
            _387 <= _92;
        33:
            _387 <= _93;
        34:
            _387 <= _94;
        35:
            _387 <= _95;
        36:
            _387 <= _96;
        37:
            _387 <= _97;
        38:
            _387 <= _98;
        39:
            _387 <= _99;
        40:
            _387 <= _100;
        41:
            _387 <= _101;
        42:
            _387 <= _102;
        43:
            _387 <= _103;
        44:
            _387 <= _104;
        45:
            _387 <= _105;
        46:
            _387 <= _106;
        47:
            _387 <= _107;
        48:
            _387 <= _108;
        49:
            _387 <= _109;
        50:
            _387 <= _110;
        51:
            _387 <= _111;
        52:
            _387 <= _112;
        53:
            _387 <= _113;
        54:
            _387 <= _114;
        55:
            _387 <= _115;
        56:
            _387 <= _116;
        57:
            _387 <= _117;
        58:
            _387 <= _118;
        59:
            _387 <= _119;
        60:
            _387 <= _120;
        61:
            _387 <= _121;
        62:
            _387 <= _122;
        63:
            _387 <= _123;
        64:
            _387 <= _124;
        65:
            _387 <= _125;
        66:
            _387 <= _126;
        67:
            _387 <= _127;
        68:
            _387 <= _128;
        69:
            _387 <= _129;
        70:
            _387 <= _130;
        71:
            _387 <= _131;
        72:
            _387 <= _132;
        73:
            _387 <= _133;
        74:
            _387 <= _134;
        75:
            _387 <= _135;
        76:
            _387 <= _136;
        77:
            _387 <= _137;
        78:
            _387 <= _138;
        79:
            _387 <= _139;
        80:
            _387 <= _140;
        81:
            _387 <= _141;
        82:
            _387 <= _142;
        83:
            _387 <= _143;
        84:
            _387 <= _144;
        85:
            _387 <= _145;
        86:
            _387 <= _146;
        87:
            _387 <= _147;
        88:
            _387 <= _148;
        89:
            _387 <= _149;
        90:
            _387 <= _150;
        91:
            _387 <= _151;
        92:
            _387 <= _152;
        93:
            _387 <= _153;
        94:
            _387 <= _154;
        95:
            _387 <= _155;
        96:
            _387 <= _156;
        97:
            _387 <= _157;
        98:
            _387 <= _158;
        99:
            _387 <= _159;
        100:
            _387 <= _160;
        101:
            _387 <= _161;
        102:
            _387 <= _162;
        103:
            _387 <= _163;
        104:
            _387 <= _164;
        105:
            _387 <= _165;
        106:
            _387 <= _166;
        107:
            _387 <= _167;
        108:
            _387 <= _168;
        109:
            _387 <= _169;
        110:
            _387 <= _170;
        111:
            _387 <= _171;
        112:
            _387 <= _172;
        113:
            _387 <= _173;
        114:
            _387 <= _174;
        115:
            _387 <= _175;
        116:
            _387 <= _176;
        117:
            _387 <= _177;
        118:
            _387 <= _178;
        119:
            _387 <= _179;
        120:
            _387 <= _180;
        121:
            _387 <= _181;
        122:
            _387 <= _182;
        123:
            _387 <= _183;
        124:
            _387 <= _184;
        125:
            _387 <= _185;
        126:
            _387 <= _186;
        default:
            _387 <= _187;
        endcase
    end
    assign _390 = _387 < _389;
    assign _391 = ~ _390;
    assign _384 = _50 < _213;
    assign _392 = _384 & _391;
    assign _518 = _392 ? _387 : _389;
    always @* begin
        case (_193)
        0:
            _246 <= _60;
        1:
            _246 <= _61;
        2:
            _246 <= _62;
        3:
            _246 <= _63;
        4:
            _246 <= _64;
        5:
            _246 <= _65;
        6:
            _246 <= _66;
        7:
            _246 <= _67;
        8:
            _246 <= _68;
        9:
            _246 <= _69;
        10:
            _246 <= _70;
        11:
            _246 <= _71;
        12:
            _246 <= _72;
        13:
            _246 <= _73;
        14:
            _246 <= _74;
        15:
            _246 <= _75;
        16:
            _246 <= _76;
        17:
            _246 <= _77;
        18:
            _246 <= _78;
        19:
            _246 <= _79;
        20:
            _246 <= _80;
        21:
            _246 <= _81;
        22:
            _246 <= _82;
        23:
            _246 <= _83;
        24:
            _246 <= _84;
        25:
            _246 <= _85;
        26:
            _246 <= _86;
        27:
            _246 <= _87;
        28:
            _246 <= _88;
        29:
            _246 <= _89;
        30:
            _246 <= _90;
        31:
            _246 <= _91;
        32:
            _246 <= _92;
        33:
            _246 <= _93;
        34:
            _246 <= _94;
        35:
            _246 <= _95;
        36:
            _246 <= _96;
        37:
            _246 <= _97;
        38:
            _246 <= _98;
        39:
            _246 <= _99;
        40:
            _246 <= _100;
        41:
            _246 <= _101;
        42:
            _246 <= _102;
        43:
            _246 <= _103;
        44:
            _246 <= _104;
        45:
            _246 <= _105;
        46:
            _246 <= _106;
        47:
            _246 <= _107;
        48:
            _246 <= _108;
        49:
            _246 <= _109;
        50:
            _246 <= _110;
        51:
            _246 <= _111;
        52:
            _246 <= _112;
        53:
            _246 <= _113;
        54:
            _246 <= _114;
        55:
            _246 <= _115;
        56:
            _246 <= _116;
        57:
            _246 <= _117;
        58:
            _246 <= _118;
        59:
            _246 <= _119;
        60:
            _246 <= _120;
        61:
            _246 <= _121;
        62:
            _246 <= _122;
        63:
            _246 <= _123;
        64:
            _246 <= _124;
        65:
            _246 <= _125;
        66:
            _246 <= _126;
        67:
            _246 <= _127;
        68:
            _246 <= _128;
        69:
            _246 <= _129;
        70:
            _246 <= _130;
        71:
            _246 <= _131;
        72:
            _246 <= _132;
        73:
            _246 <= _133;
        74:
            _246 <= _134;
        75:
            _246 <= _135;
        76:
            _246 <= _136;
        77:
            _246 <= _137;
        78:
            _246 <= _138;
        79:
            _246 <= _139;
        80:
            _246 <= _140;
        81:
            _246 <= _141;
        82:
            _246 <= _142;
        83:
            _246 <= _143;
        84:
            _246 <= _144;
        85:
            _246 <= _145;
        86:
            _246 <= _146;
        87:
            _246 <= _147;
        88:
            _246 <= _148;
        89:
            _246 <= _149;
        90:
            _246 <= _150;
        91:
            _246 <= _151;
        92:
            _246 <= _152;
        93:
            _246 <= _153;
        94:
            _246 <= _154;
        95:
            _246 <= _155;
        96:
            _246 <= _156;
        97:
            _246 <= _157;
        98:
            _246 <= _158;
        99:
            _246 <= _159;
        100:
            _246 <= _160;
        101:
            _246 <= _161;
        102:
            _246 <= _162;
        103:
            _246 <= _163;
        104:
            _246 <= _164;
        105:
            _246 <= _165;
        106:
            _246 <= _166;
        107:
            _246 <= _167;
        108:
            _246 <= _168;
        109:
            _246 <= _169;
        110:
            _246 <= _170;
        111:
            _246 <= _171;
        112:
            _246 <= _172;
        113:
            _246 <= _173;
        114:
            _246 <= _174;
        115:
            _246 <= _175;
        116:
            _246 <= _176;
        117:
            _246 <= _177;
        118:
            _246 <= _178;
        119:
            _246 <= _179;
        120:
            _246 <= _180;
        121:
            _246 <= _181;
        122:
            _246 <= _182;
        123:
            _246 <= _183;
        124:
            _246 <= _184;
        125:
            _246 <= _185;
        126:
            _246 <= _186;
        default:
            _246 <= _187;
        endcase
    end
    assign _250 = _246 < _249;
    assign _251 = ~ _250;
    assign _244 = _50 < _213;
    assign _252 = _244 & _251;
    assign _388 = _252 ? _246 : _249;
    assign _206 = 8'b00000000;
    assign _207 = _193 < _206;
    assign _208 = ~ _207;
    assign _209 = _48 & _208;
    assign _389 = _209 ? _388 : _249;
    assign _203 = _193 < _846;
    assign _204 = ~ _203;
    assign _205 = _48 & _204;
    assign _519 = _205 ? _518 : _389;
    assign _199 = _193 < _835;
    assign _200 = ~ _199;
    assign _201 = _48 & _200;
    assign _649 = _201 ? _648 : _519;
    assign _195 = _193 < _824;
    assign _196 = ~ _195;
    assign _197 = _48 & _196;
    assign _861 = _197 ? _860 : _649;
    assign _187 = _15[511:508];
    assign _186 = _15[507:504];
    assign _185 = _15[503:500];
    assign _184 = _15[499:496];
    assign _183 = _15[495:492];
    assign _182 = _15[491:488];
    assign _181 = _15[487:484];
    assign _180 = _15[483:480];
    assign _179 = _15[479:476];
    assign _178 = _15[475:472];
    assign _177 = _15[471:468];
    assign _176 = _15[467:464];
    assign _175 = _15[463:460];
    assign _174 = _15[459:456];
    assign _173 = _15[455:452];
    assign _172 = _15[451:448];
    assign _171 = _15[447:444];
    assign _170 = _15[443:440];
    assign _169 = _15[439:436];
    assign _168 = _15[435:432];
    assign _167 = _15[431:428];
    assign _166 = _15[427:424];
    assign _165 = _15[423:420];
    assign _164 = _15[419:416];
    assign _163 = _15[415:412];
    assign _162 = _15[411:408];
    assign _161 = _15[407:404];
    assign _160 = _15[403:400];
    assign _159 = _15[399:396];
    assign _158 = _15[395:392];
    assign _157 = _15[391:388];
    assign _156 = _15[387:384];
    assign _155 = _15[383:380];
    assign _154 = _15[379:376];
    assign _153 = _15[375:372];
    assign _152 = _15[371:368];
    assign _151 = _15[367:364];
    assign _150 = _15[363:360];
    assign _149 = _15[359:356];
    assign _148 = _15[355:352];
    assign _147 = _15[351:348];
    assign _146 = _15[347:344];
    assign _145 = _15[343:340];
    assign _144 = _15[339:336];
    assign _143 = _15[335:332];
    assign _142 = _15[331:328];
    assign _141 = _15[327:324];
    assign _140 = _15[323:320];
    assign _139 = _15[319:316];
    assign _138 = _15[315:312];
    assign _137 = _15[311:308];
    assign _136 = _15[307:304];
    assign _135 = _15[303:300];
    assign _134 = _15[299:296];
    assign _133 = _15[295:292];
    assign _132 = _15[291:288];
    assign _131 = _15[287:284];
    assign _130 = _15[283:280];
    assign _129 = _15[279:276];
    assign _128 = _15[275:272];
    assign _127 = _15[271:268];
    assign _126 = _15[267:264];
    assign _125 = _15[263:260];
    assign _124 = _15[259:256];
    assign _123 = _15[255:252];
    assign _122 = _15[251:248];
    assign _121 = _15[247:244];
    assign _120 = _15[243:240];
    assign _119 = _15[239:236];
    assign _118 = _15[235:232];
    assign _117 = _15[231:228];
    assign _116 = _15[227:224];
    assign _115 = _15[223:220];
    assign _114 = _15[219:216];
    assign _113 = _15[215:212];
    assign _112 = _15[211:208];
    assign _111 = _15[207:204];
    assign _110 = _15[203:200];
    assign _109 = _15[199:196];
    assign _108 = _15[195:192];
    assign _107 = _15[191:188];
    assign _106 = _15[187:184];
    assign _105 = _15[183:180];
    assign _104 = _15[179:176];
    assign _103 = _15[175:172];
    assign _102 = _15[171:168];
    assign _101 = _15[167:164];
    assign _100 = _15[163:160];
    assign _99 = _15[159:156];
    assign _98 = _15[155:152];
    assign _97 = _15[151:148];
    assign _96 = _15[147:144];
    assign _95 = _15[143:140];
    assign _94 = _15[139:136];
    assign _93 = _15[135:132];
    assign _92 = _15[131:128];
    assign _91 = _15[127:124];
    assign _90 = _15[123:120];
    assign _89 = _15[119:116];
    assign _88 = _15[115:112];
    assign _87 = _15[111:108];
    assign _86 = _15[107:104];
    assign _85 = _15[103:100];
    assign _84 = _15[99:96];
    assign _83 = _15[95:92];
    assign _82 = _15[91:88];
    assign _81 = _15[87:84];
    assign _80 = _15[83:80];
    assign _79 = _15[79:76];
    assign _78 = _15[75:72];
    assign _77 = _15[71:68];
    assign _76 = _15[67:64];
    assign _75 = _15[63:60];
    assign _74 = _15[59:56];
    assign _73 = _15[55:52];
    assign _72 = _15[51:48];
    assign _71 = _15[47:44];
    assign _70 = _15[43:40];
    assign _69 = _15[39:36];
    assign _68 = _15[35:32];
    assign _67 = _15[31:28];
    assign _66 = _15[27:24];
    assign _65 = _15[23:20];
    assign _64 = _15[19:16];
    assign _63 = _15[15:12];
    assign _62 = _15[11:8];
    assign _61 = _15[7:4];
    assign _15 = data;
    assign _60 = _15[3:0];
    always @* begin
        case (_57)
        0:
            _857 <= _60;
        1:
            _857 <= _61;
        2:
            _857 <= _62;
        3:
            _857 <= _63;
        4:
            _857 <= _64;
        5:
            _857 <= _65;
        6:
            _857 <= _66;
        7:
            _857 <= _67;
        8:
            _857 <= _68;
        9:
            _857 <= _69;
        10:
            _857 <= _70;
        11:
            _857 <= _71;
        12:
            _857 <= _72;
        13:
            _857 <= _73;
        14:
            _857 <= _74;
        15:
            _857 <= _75;
        16:
            _857 <= _76;
        17:
            _857 <= _77;
        18:
            _857 <= _78;
        19:
            _857 <= _79;
        20:
            _857 <= _80;
        21:
            _857 <= _81;
        22:
            _857 <= _82;
        23:
            _857 <= _83;
        24:
            _857 <= _84;
        25:
            _857 <= _85;
        26:
            _857 <= _86;
        27:
            _857 <= _87;
        28:
            _857 <= _88;
        29:
            _857 <= _89;
        30:
            _857 <= _90;
        31:
            _857 <= _91;
        32:
            _857 <= _92;
        33:
            _857 <= _93;
        34:
            _857 <= _94;
        35:
            _857 <= _95;
        36:
            _857 <= _96;
        37:
            _857 <= _97;
        38:
            _857 <= _98;
        39:
            _857 <= _99;
        40:
            _857 <= _100;
        41:
            _857 <= _101;
        42:
            _857 <= _102;
        43:
            _857 <= _103;
        44:
            _857 <= _104;
        45:
            _857 <= _105;
        46:
            _857 <= _106;
        47:
            _857 <= _107;
        48:
            _857 <= _108;
        49:
            _857 <= _109;
        50:
            _857 <= _110;
        51:
            _857 <= _111;
        52:
            _857 <= _112;
        53:
            _857 <= _113;
        54:
            _857 <= _114;
        55:
            _857 <= _115;
        56:
            _857 <= _116;
        57:
            _857 <= _117;
        58:
            _857 <= _118;
        59:
            _857 <= _119;
        60:
            _857 <= _120;
        61:
            _857 <= _121;
        62:
            _857 <= _122;
        63:
            _857 <= _123;
        64:
            _857 <= _124;
        65:
            _857 <= _125;
        66:
            _857 <= _126;
        67:
            _857 <= _127;
        68:
            _857 <= _128;
        69:
            _857 <= _129;
        70:
            _857 <= _130;
        71:
            _857 <= _131;
        72:
            _857 <= _132;
        73:
            _857 <= _133;
        74:
            _857 <= _134;
        75:
            _857 <= _135;
        76:
            _857 <= _136;
        77:
            _857 <= _137;
        78:
            _857 <= _138;
        79:
            _857 <= _139;
        80:
            _857 <= _140;
        81:
            _857 <= _141;
        82:
            _857 <= _142;
        83:
            _857 <= _143;
        84:
            _857 <= _144;
        85:
            _857 <= _145;
        86:
            _857 <= _146;
        87:
            _857 <= _147;
        88:
            _857 <= _148;
        89:
            _857 <= _149;
        90:
            _857 <= _150;
        91:
            _857 <= _151;
        92:
            _857 <= _152;
        93:
            _857 <= _153;
        94:
            _857 <= _154;
        95:
            _857 <= _155;
        96:
            _857 <= _156;
        97:
            _857 <= _157;
        98:
            _857 <= _158;
        99:
            _857 <= _159;
        100:
            _857 <= _160;
        101:
            _857 <= _161;
        102:
            _857 <= _162;
        103:
            _857 <= _163;
        104:
            _857 <= _164;
        105:
            _857 <= _165;
        106:
            _857 <= _166;
        107:
            _857 <= _167;
        108:
            _857 <= _168;
        109:
            _857 <= _169;
        110:
            _857 <= _170;
        111:
            _857 <= _171;
        112:
            _857 <= _172;
        113:
            _857 <= _173;
        114:
            _857 <= _174;
        115:
            _857 <= _175;
        116:
            _857 <= _176;
        117:
            _857 <= _177;
        118:
            _857 <= _178;
        119:
            _857 <= _179;
        120:
            _857 <= _180;
        121:
            _857 <= _181;
        122:
            _857 <= _182;
        123:
            _857 <= _183;
        124:
            _857 <= _184;
        125:
            _857 <= _185;
        126:
            _857 <= _186;
        default:
            _857 <= _187;
        endcase
    end
    assign _855 = _50 < _25;
    assign _858 = _855 ? _857 : _50;
    assign _859 = _40 ? _858 : _249;
    assign _862 = _48 ? _861 : _859;
    assign _16 = _862;
    always @(posedge _22) begin
        if (_20)
            _249 <= _50;
        else
            _249 <= _16;
    end
    assign _910 = { _985,
                    _249 };
    assign _908 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign _907 = _50 < _213;
    assign _911 = _907 ? _910 : _908;
    assign _905 = _640 < _213;
    assign _918 = _905 ? _917 : _911;
    assign _903 = _637 < _213;
    assign _925 = _903 ? _924 : _918;
    assign _901 = _634 < _213;
    assign _932 = _901 ? _931 : _925;
    assign _899 = _631 < _213;
    assign _939 = _899 ? _938 : _932;
    assign _897 = _628 < _213;
    assign _946 = _897 ? _945 : _939;
    assign _895 = _625 < _213;
    assign _953 = _895 ? _952 : _946;
    assign _893 = _622 < _213;
    assign _960 = _893 ? _959 : _953;
    assign _891 = _619 < _213;
    assign _967 = _891 ? _966 : _960;
    assign _889 = _616 < _213;
    assign _974 = _889 ? _973 : _967;
    assign _887 = _613 < _213;
    assign _981 = _887 ? _980 : _974;
    assign _18 = start;
    assign _35 = 2'b10;
    assign _36 = _34 == _35;
    assign _37 = 2'b00;
    assign _879 = 2'b01;
    assign vdd = 1'b1;
    assign _20 = clear;
    assign _22 = clock;
    assign _869 = _193 - _813;
    assign _871 = _867 ? _206 : _869;
    assign _864 = _57 - _846;
    assign _865 = _40 ? _864 : _193;
    assign _872 = _48 ? _871 : _865;
    assign _23 = _872;
    always @(posedge _22) begin
        if (_20)
            _193 <= _206;
        else
            _193 <= _23;
    end
    assign _867 = _193 < _813;
    assign _881 = _867 ? _35 : _879;
    assign _25 = k;
    assign _56 = { _50,
                   _25 };
    assign _27 = length;
    assign _57 = _27 - _56;
    assign _874 = _57 == _206;
    assign _877 = _874 ? _35 : _879;
    assign _878 = _40 ? _877 : _34;
    assign _48 = _34 == _879;
    assign _882 = _48 ? _881 : _878;
    assign _28 = _882;
    always @(posedge _22) begin
        if (_20)
            _34 <= _37;
        else
            _34 <= _28;
    end
    assign _38 = _34 == _37;
    assign _39 = _38 | _36;
    assign _40 = _39 & _18;
    assign _883 = _40 ? _25 : _213;
    assign _29 = _883;
    always @(posedge _22) begin
        if (_20)
            _213 <= _50;
        else
            _213 <= _29;
    end
    assign _885 = _734 < _213;
    assign _988 = _885 ? _987 : _981;
    assign result = _988;
    assign done_ = _43;

endmodule
