module day2 (
    from_,
    to_,
    last,
    clear,
    clock,
    pair_valid,
    load,
    sum_p1,
    sum_p2,
    ready,
    done_,
    family_index
);

    input [63:0] from_;
    input [63:0] to_;
    input last;
    input clear;
    input clock;
    input pair_valid;
    input load;
    output [63:0] sum_p1;
    output [63:0] sum_p2;
    output ready;
    output done_;
    output [3:0] family_index;

    wire [63:0] _45;
    wire _766;
    wire _747;
    wire _749;
    wire _751;
    wire _753;
    wire _755;
    wire _757;
    wire _759;
    wire _761;
    wire _763;
    wire _765;
    wire _767;
    wire _768;
    wire _769;
    wire _770;
    wire [63:0] _1933;
    wire [63:0] _1934;
    wire _42;
    wire _43;
    wire [63:0] _1935;
    wire [63:0] _1937;
    wire [63:0] _4;
    reg [63:0] _46;
    wire _1945;
    wire _1947;
    wire _1949;
    wire _1951;
    wire _1953;
    wire _1954;
    wire _1955;
    wire _1956;
    wire _1957;
    wire _1958;
    wire _1959;
    wire _1961;
    wire _1963;
    wire _1964;
    wire [63:0] _1966;
    wire [63:0] _1967;
    wire _1938;
    wire _1939;
    wire [63:0] _1968;
    wire [63:0] _1970;
    wire [63:0] _5;
    reg [63:0] _1942;
    wire [63:0] _1974;
    wire [63:0] _1975;
    wire _1925;
    wire [63:0] _1922;
    wire [63:0] _1923;
    wire [62:0] _1924;
    wire [63:0] _1926;
    wire _1927;
    wire _1928;
    wire _1916;
    wire [63:0] _1913;
    wire [63:0] _1914;
    wire [62:0] _1915;
    wire [63:0] _1917;
    wire _1918;
    wire _1919;
    wire _1907;
    wire [63:0] _1904;
    wire [63:0] _1905;
    wire [62:0] _1906;
    wire [63:0] _1908;
    wire _1909;
    wire _1910;
    wire _1898;
    wire [63:0] _1895;
    wire [63:0] _1896;
    wire [62:0] _1897;
    wire [63:0] _1899;
    wire _1900;
    wire _1901;
    wire _1889;
    wire [63:0] _1886;
    wire [63:0] _1887;
    wire [62:0] _1888;
    wire [63:0] _1890;
    wire _1891;
    wire _1892;
    wire _1880;
    wire [63:0] _1877;
    wire [63:0] _1878;
    wire [62:0] _1879;
    wire [63:0] _1881;
    wire _1882;
    wire _1883;
    wire _1871;
    wire [63:0] _1868;
    wire [63:0] _1869;
    wire [62:0] _1870;
    wire [63:0] _1872;
    wire _1873;
    wire _1874;
    wire _1862;
    wire [63:0] _1859;
    wire [63:0] _1860;
    wire [62:0] _1861;
    wire [63:0] _1863;
    wire _1864;
    wire _1865;
    wire _1853;
    wire [63:0] _1850;
    wire [63:0] _1851;
    wire [62:0] _1852;
    wire [63:0] _1854;
    wire _1855;
    wire _1856;
    wire _1844;
    wire [63:0] _1841;
    wire [63:0] _1842;
    wire [62:0] _1843;
    wire [63:0] _1845;
    wire _1846;
    wire _1847;
    wire _1835;
    wire [63:0] _1832;
    wire [63:0] _1833;
    wire [62:0] _1834;
    wire [63:0] _1836;
    wire _1837;
    wire _1838;
    wire _1826;
    wire [63:0] _1823;
    wire [63:0] _1824;
    wire [62:0] _1825;
    wire [63:0] _1827;
    wire _1828;
    wire _1829;
    wire _1817;
    wire [63:0] _1814;
    wire [63:0] _1815;
    wire [62:0] _1816;
    wire [63:0] _1818;
    wire _1819;
    wire _1820;
    wire _1808;
    wire [63:0] _1805;
    wire [63:0] _1806;
    wire [62:0] _1807;
    wire [63:0] _1809;
    wire _1810;
    wire _1811;
    wire _1799;
    wire [63:0] _1796;
    wire [63:0] _1797;
    wire [62:0] _1798;
    wire [63:0] _1800;
    wire _1801;
    wire _1802;
    wire _1790;
    wire [63:0] _1787;
    wire [63:0] _1788;
    wire [62:0] _1789;
    wire [63:0] _1791;
    wire _1792;
    wire _1793;
    wire _1781;
    wire [63:0] _1778;
    wire [63:0] _1779;
    wire [62:0] _1780;
    wire [63:0] _1782;
    wire _1783;
    wire _1784;
    wire _1772;
    wire [63:0] _1769;
    wire [63:0] _1770;
    wire [62:0] _1771;
    wire [63:0] _1773;
    wire _1774;
    wire _1775;
    wire _1763;
    wire [63:0] _1760;
    wire [63:0] _1761;
    wire [62:0] _1762;
    wire [63:0] _1764;
    wire _1765;
    wire _1766;
    wire _1754;
    wire [63:0] _1751;
    wire [63:0] _1752;
    wire [62:0] _1753;
    wire [63:0] _1755;
    wire _1756;
    wire _1757;
    wire _1745;
    wire [63:0] _1742;
    wire [63:0] _1743;
    wire [62:0] _1744;
    wire [63:0] _1746;
    wire _1747;
    wire _1748;
    wire _1736;
    wire [63:0] _1733;
    wire [63:0] _1734;
    wire [62:0] _1735;
    wire [63:0] _1737;
    wire _1738;
    wire _1739;
    wire _1727;
    wire [63:0] _1724;
    wire [63:0] _1725;
    wire [62:0] _1726;
    wire [63:0] _1728;
    wire _1729;
    wire _1730;
    wire _1718;
    wire [63:0] _1715;
    wire [63:0] _1716;
    wire [62:0] _1717;
    wire [63:0] _1719;
    wire _1720;
    wire _1721;
    wire _1709;
    wire [63:0] _1706;
    wire [63:0] _1707;
    wire [62:0] _1708;
    wire [63:0] _1710;
    wire _1711;
    wire _1712;
    wire _1700;
    wire [63:0] _1697;
    wire [63:0] _1698;
    wire [62:0] _1699;
    wire [63:0] _1701;
    wire _1702;
    wire _1703;
    wire _1691;
    wire [63:0] _1688;
    wire [63:0] _1689;
    wire [62:0] _1690;
    wire [63:0] _1692;
    wire _1693;
    wire _1694;
    wire _1682;
    wire [63:0] _1679;
    wire [63:0] _1680;
    wire [62:0] _1681;
    wire [63:0] _1683;
    wire _1684;
    wire _1685;
    wire _1673;
    wire [63:0] _1670;
    wire [63:0] _1671;
    wire [62:0] _1672;
    wire [63:0] _1674;
    wire _1675;
    wire _1676;
    wire _1664;
    wire [63:0] _1661;
    wire [63:0] _1662;
    wire [62:0] _1663;
    wire [63:0] _1665;
    wire _1666;
    wire _1667;
    wire _1655;
    wire [63:0] _1652;
    wire [63:0] _1653;
    wire [62:0] _1654;
    wire [63:0] _1656;
    wire _1657;
    wire _1658;
    wire _1646;
    wire [63:0] _1643;
    wire [63:0] _1644;
    wire [62:0] _1645;
    wire [63:0] _1647;
    wire _1648;
    wire _1649;
    wire _1637;
    wire [63:0] _1634;
    wire [63:0] _1635;
    wire [62:0] _1636;
    wire [63:0] _1638;
    wire _1639;
    wire _1640;
    wire _1628;
    wire [63:0] _1625;
    wire [63:0] _1626;
    wire [62:0] _1627;
    wire [63:0] _1629;
    wire _1630;
    wire _1631;
    wire _1619;
    wire [63:0] _1616;
    wire [63:0] _1617;
    wire [62:0] _1618;
    wire [63:0] _1620;
    wire _1621;
    wire _1622;
    wire _1610;
    wire [63:0] _1607;
    wire [63:0] _1608;
    wire [62:0] _1609;
    wire [63:0] _1611;
    wire _1612;
    wire _1613;
    wire _1601;
    wire [63:0] _1598;
    wire [63:0] _1599;
    wire [62:0] _1600;
    wire [63:0] _1602;
    wire _1603;
    wire _1604;
    wire _1592;
    wire [63:0] _1589;
    wire [63:0] _1590;
    wire [62:0] _1591;
    wire [63:0] _1593;
    wire _1594;
    wire _1595;
    wire _1583;
    wire [63:0] _1580;
    wire [63:0] _1581;
    wire [62:0] _1582;
    wire [63:0] _1584;
    wire _1585;
    wire _1586;
    wire _1574;
    wire [63:0] _1571;
    wire [63:0] _1572;
    wire [62:0] _1573;
    wire [63:0] _1575;
    wire _1576;
    wire _1577;
    wire _1565;
    wire [63:0] _1562;
    wire [63:0] _1563;
    wire [62:0] _1564;
    wire [63:0] _1566;
    wire _1567;
    wire _1568;
    wire _1556;
    wire [63:0] _1553;
    wire [63:0] _1554;
    wire [62:0] _1555;
    wire [63:0] _1557;
    wire _1558;
    wire _1559;
    wire _1547;
    wire [63:0] _1544;
    wire [63:0] _1545;
    wire [62:0] _1546;
    wire [63:0] _1548;
    wire _1549;
    wire _1550;
    wire _1538;
    wire [63:0] _1535;
    wire [63:0] _1536;
    wire [62:0] _1537;
    wire [63:0] _1539;
    wire _1540;
    wire _1541;
    wire _1529;
    wire [63:0] _1526;
    wire [63:0] _1527;
    wire [62:0] _1528;
    wire [63:0] _1530;
    wire _1531;
    wire _1532;
    wire _1520;
    wire [63:0] _1517;
    wire [63:0] _1518;
    wire [62:0] _1519;
    wire [63:0] _1521;
    wire _1522;
    wire _1523;
    wire _1511;
    wire [63:0] _1508;
    wire [63:0] _1509;
    wire [62:0] _1510;
    wire [63:0] _1512;
    wire _1513;
    wire _1514;
    wire _1502;
    wire [63:0] _1499;
    wire [63:0] _1500;
    wire [62:0] _1501;
    wire [63:0] _1503;
    wire _1504;
    wire _1505;
    wire _1493;
    wire [63:0] _1490;
    wire [63:0] _1491;
    wire [62:0] _1492;
    wire [63:0] _1494;
    wire _1495;
    wire _1496;
    wire _1484;
    wire [63:0] _1481;
    wire [63:0] _1482;
    wire [62:0] _1483;
    wire [63:0] _1485;
    wire _1486;
    wire _1487;
    wire _1475;
    wire [63:0] _1472;
    wire [63:0] _1473;
    wire [62:0] _1474;
    wire [63:0] _1476;
    wire _1477;
    wire _1478;
    wire _1466;
    wire [63:0] _1463;
    wire [63:0] _1464;
    wire [62:0] _1465;
    wire [63:0] _1467;
    wire _1468;
    wire _1469;
    wire _1457;
    wire [63:0] _1454;
    wire [63:0] _1455;
    wire [62:0] _1456;
    wire [63:0] _1458;
    wire _1459;
    wire _1460;
    wire _1448;
    wire [63:0] _1445;
    wire [63:0] _1446;
    wire [62:0] _1447;
    wire [63:0] _1449;
    wire _1450;
    wire _1451;
    wire _1439;
    wire [63:0] _1436;
    wire [63:0] _1437;
    wire [62:0] _1438;
    wire [63:0] _1440;
    wire _1441;
    wire _1442;
    wire _1430;
    wire [63:0] _1427;
    wire [63:0] _1428;
    wire [62:0] _1429;
    wire [63:0] _1431;
    wire _1432;
    wire _1433;
    wire _1421;
    wire [63:0] _1418;
    wire [63:0] _1419;
    wire [62:0] _1420;
    wire [63:0] _1422;
    wire _1423;
    wire _1424;
    wire _1412;
    wire [63:0] _1409;
    wire [63:0] _1410;
    wire [62:0] _1411;
    wire [63:0] _1413;
    wire _1414;
    wire _1415;
    wire _1403;
    wire [63:0] _1400;
    wire [63:0] _1401;
    wire [62:0] _1402;
    wire [63:0] _1404;
    wire _1405;
    wire _1406;
    wire _1394;
    wire [63:0] _1391;
    wire [63:0] _1392;
    wire [62:0] _1393;
    wire [63:0] _1395;
    wire _1396;
    wire _1397;
    wire _1385;
    wire [63:0] _1382;
    wire [63:0] _1383;
    wire [62:0] _1384;
    wire [63:0] _1386;
    wire _1387;
    wire _1388;
    wire _1376;
    wire [63:0] _1373;
    wire [63:0] _1374;
    wire [62:0] _1375;
    wire [63:0] _1377;
    wire _1378;
    wire _1379;
    wire _1367;
    wire [63:0] _1364;
    wire [63:0] _1365;
    wire [62:0] _1366;
    wire [63:0] _1368;
    wire _1369;
    wire _1370;
    wire [63:0] _1359;
    wire [63:0] _1353;
    wire [63:0] _1354;
    wire [127:0] _1355;
    wire [63:0] _1356;
    wire _1357;
    wire [62:0] _1352;
    wire [63:0] _1358;
    wire _1360;
    wire _1361;
    wire [63:0] _1362;
    wire [62:0] _1363;
    wire [63:0] _1371;
    wire [62:0] _1372;
    wire [63:0] _1380;
    wire [62:0] _1381;
    wire [63:0] _1389;
    wire [62:0] _1390;
    wire [63:0] _1398;
    wire [62:0] _1399;
    wire [63:0] _1407;
    wire [62:0] _1408;
    wire [63:0] _1416;
    wire [62:0] _1417;
    wire [63:0] _1425;
    wire [62:0] _1426;
    wire [63:0] _1434;
    wire [62:0] _1435;
    wire [63:0] _1443;
    wire [62:0] _1444;
    wire [63:0] _1452;
    wire [62:0] _1453;
    wire [63:0] _1461;
    wire [62:0] _1462;
    wire [63:0] _1470;
    wire [62:0] _1471;
    wire [63:0] _1479;
    wire [62:0] _1480;
    wire [63:0] _1488;
    wire [62:0] _1489;
    wire [63:0] _1497;
    wire [62:0] _1498;
    wire [63:0] _1506;
    wire [62:0] _1507;
    wire [63:0] _1515;
    wire [62:0] _1516;
    wire [63:0] _1524;
    wire [62:0] _1525;
    wire [63:0] _1533;
    wire [62:0] _1534;
    wire [63:0] _1542;
    wire [62:0] _1543;
    wire [63:0] _1551;
    wire [62:0] _1552;
    wire [63:0] _1560;
    wire [62:0] _1561;
    wire [63:0] _1569;
    wire [62:0] _1570;
    wire [63:0] _1578;
    wire [62:0] _1579;
    wire [63:0] _1587;
    wire [62:0] _1588;
    wire [63:0] _1596;
    wire [62:0] _1597;
    wire [63:0] _1605;
    wire [62:0] _1606;
    wire [63:0] _1614;
    wire [62:0] _1615;
    wire [63:0] _1623;
    wire [62:0] _1624;
    wire [63:0] _1632;
    wire [62:0] _1633;
    wire [63:0] _1641;
    wire [62:0] _1642;
    wire [63:0] _1650;
    wire [62:0] _1651;
    wire [63:0] _1659;
    wire [62:0] _1660;
    wire [63:0] _1668;
    wire [62:0] _1669;
    wire [63:0] _1677;
    wire [62:0] _1678;
    wire [63:0] _1686;
    wire [62:0] _1687;
    wire [63:0] _1695;
    wire [62:0] _1696;
    wire [63:0] _1704;
    wire [62:0] _1705;
    wire [63:0] _1713;
    wire [62:0] _1714;
    wire [63:0] _1722;
    wire [62:0] _1723;
    wire [63:0] _1731;
    wire [62:0] _1732;
    wire [63:0] _1740;
    wire [62:0] _1741;
    wire [63:0] _1749;
    wire [62:0] _1750;
    wire [63:0] _1758;
    wire [62:0] _1759;
    wire [63:0] _1767;
    wire [62:0] _1768;
    wire [63:0] _1776;
    wire [62:0] _1777;
    wire [63:0] _1785;
    wire [62:0] _1786;
    wire [63:0] _1794;
    wire [62:0] _1795;
    wire [63:0] _1803;
    wire [62:0] _1804;
    wire [63:0] _1812;
    wire [62:0] _1813;
    wire [63:0] _1821;
    wire [62:0] _1822;
    wire [63:0] _1830;
    wire [62:0] _1831;
    wire [63:0] _1839;
    wire [62:0] _1840;
    wire [63:0] _1848;
    wire [62:0] _1849;
    wire [63:0] _1857;
    wire [62:0] _1858;
    wire [63:0] _1866;
    wire [62:0] _1867;
    wire [63:0] _1875;
    wire [62:0] _1876;
    wire [63:0] _1884;
    wire [62:0] _1885;
    wire [63:0] _1893;
    wire [62:0] _1894;
    wire [63:0] _1902;
    wire [62:0] _1903;
    wire [63:0] _1911;
    wire [62:0] _1912;
    wire [63:0] _1920;
    wire [62:0] _1921;
    wire [63:0] _1929;
    wire [127:0] _1930;
    wire [63:0] _1931;
    wire _1342;
    wire [63:0] _1339;
    wire [63:0] _1340;
    wire [62:0] _1341;
    wire [63:0] _1343;
    wire _1344;
    wire _1345;
    wire _1333;
    wire [63:0] _1330;
    wire [63:0] _1331;
    wire [62:0] _1332;
    wire [63:0] _1334;
    wire _1335;
    wire _1336;
    wire _1324;
    wire [63:0] _1321;
    wire [63:0] _1322;
    wire [62:0] _1323;
    wire [63:0] _1325;
    wire _1326;
    wire _1327;
    wire _1315;
    wire [63:0] _1312;
    wire [63:0] _1313;
    wire [62:0] _1314;
    wire [63:0] _1316;
    wire _1317;
    wire _1318;
    wire _1306;
    wire [63:0] _1303;
    wire [63:0] _1304;
    wire [62:0] _1305;
    wire [63:0] _1307;
    wire _1308;
    wire _1309;
    wire _1297;
    wire [63:0] _1294;
    wire [63:0] _1295;
    wire [62:0] _1296;
    wire [63:0] _1298;
    wire _1299;
    wire _1300;
    wire _1288;
    wire [63:0] _1285;
    wire [63:0] _1286;
    wire [62:0] _1287;
    wire [63:0] _1289;
    wire _1290;
    wire _1291;
    wire _1279;
    wire [63:0] _1276;
    wire [63:0] _1277;
    wire [62:0] _1278;
    wire [63:0] _1280;
    wire _1281;
    wire _1282;
    wire _1270;
    wire [63:0] _1267;
    wire [63:0] _1268;
    wire [62:0] _1269;
    wire [63:0] _1271;
    wire _1272;
    wire _1273;
    wire _1261;
    wire [63:0] _1258;
    wire [63:0] _1259;
    wire [62:0] _1260;
    wire [63:0] _1262;
    wire _1263;
    wire _1264;
    wire _1252;
    wire [63:0] _1249;
    wire [63:0] _1250;
    wire [62:0] _1251;
    wire [63:0] _1253;
    wire _1254;
    wire _1255;
    wire _1243;
    wire [63:0] _1240;
    wire [63:0] _1241;
    wire [62:0] _1242;
    wire [63:0] _1244;
    wire _1245;
    wire _1246;
    wire _1234;
    wire [63:0] _1231;
    wire [63:0] _1232;
    wire [62:0] _1233;
    wire [63:0] _1235;
    wire _1236;
    wire _1237;
    wire _1225;
    wire [63:0] _1222;
    wire [63:0] _1223;
    wire [62:0] _1224;
    wire [63:0] _1226;
    wire _1227;
    wire _1228;
    wire _1216;
    wire [63:0] _1213;
    wire [63:0] _1214;
    wire [62:0] _1215;
    wire [63:0] _1217;
    wire _1218;
    wire _1219;
    wire _1207;
    wire [63:0] _1204;
    wire [63:0] _1205;
    wire [62:0] _1206;
    wire [63:0] _1208;
    wire _1209;
    wire _1210;
    wire _1198;
    wire [63:0] _1195;
    wire [63:0] _1196;
    wire [62:0] _1197;
    wire [63:0] _1199;
    wire _1200;
    wire _1201;
    wire _1189;
    wire [63:0] _1186;
    wire [63:0] _1187;
    wire [62:0] _1188;
    wire [63:0] _1190;
    wire _1191;
    wire _1192;
    wire _1180;
    wire [63:0] _1177;
    wire [63:0] _1178;
    wire [62:0] _1179;
    wire [63:0] _1181;
    wire _1182;
    wire _1183;
    wire _1171;
    wire [63:0] _1168;
    wire [63:0] _1169;
    wire [62:0] _1170;
    wire [63:0] _1172;
    wire _1173;
    wire _1174;
    wire _1162;
    wire [63:0] _1159;
    wire [63:0] _1160;
    wire [62:0] _1161;
    wire [63:0] _1163;
    wire _1164;
    wire _1165;
    wire _1153;
    wire [63:0] _1150;
    wire [63:0] _1151;
    wire [62:0] _1152;
    wire [63:0] _1154;
    wire _1155;
    wire _1156;
    wire _1144;
    wire [63:0] _1141;
    wire [63:0] _1142;
    wire [62:0] _1143;
    wire [63:0] _1145;
    wire _1146;
    wire _1147;
    wire _1135;
    wire [63:0] _1132;
    wire [63:0] _1133;
    wire [62:0] _1134;
    wire [63:0] _1136;
    wire _1137;
    wire _1138;
    wire _1126;
    wire [63:0] _1123;
    wire [63:0] _1124;
    wire [62:0] _1125;
    wire [63:0] _1127;
    wire _1128;
    wire _1129;
    wire _1117;
    wire [63:0] _1114;
    wire [63:0] _1115;
    wire [62:0] _1116;
    wire [63:0] _1118;
    wire _1119;
    wire _1120;
    wire _1108;
    wire [63:0] _1105;
    wire [63:0] _1106;
    wire [62:0] _1107;
    wire [63:0] _1109;
    wire _1110;
    wire _1111;
    wire _1099;
    wire [63:0] _1096;
    wire [63:0] _1097;
    wire [62:0] _1098;
    wire [63:0] _1100;
    wire _1101;
    wire _1102;
    wire _1090;
    wire [63:0] _1087;
    wire [63:0] _1088;
    wire [62:0] _1089;
    wire [63:0] _1091;
    wire _1092;
    wire _1093;
    wire _1081;
    wire [63:0] _1078;
    wire [63:0] _1079;
    wire [62:0] _1080;
    wire [63:0] _1082;
    wire _1083;
    wire _1084;
    wire _1072;
    wire [63:0] _1069;
    wire [63:0] _1070;
    wire [62:0] _1071;
    wire [63:0] _1073;
    wire _1074;
    wire _1075;
    wire _1063;
    wire [63:0] _1060;
    wire [63:0] _1061;
    wire [62:0] _1062;
    wire [63:0] _1064;
    wire _1065;
    wire _1066;
    wire _1054;
    wire [63:0] _1051;
    wire [63:0] _1052;
    wire [62:0] _1053;
    wire [63:0] _1055;
    wire _1056;
    wire _1057;
    wire _1045;
    wire [63:0] _1042;
    wire [63:0] _1043;
    wire [62:0] _1044;
    wire [63:0] _1046;
    wire _1047;
    wire _1048;
    wire _1036;
    wire [63:0] _1033;
    wire [63:0] _1034;
    wire [62:0] _1035;
    wire [63:0] _1037;
    wire _1038;
    wire _1039;
    wire _1027;
    wire [63:0] _1024;
    wire [63:0] _1025;
    wire [62:0] _1026;
    wire [63:0] _1028;
    wire _1029;
    wire _1030;
    wire _1018;
    wire [63:0] _1015;
    wire [63:0] _1016;
    wire [62:0] _1017;
    wire [63:0] _1019;
    wire _1020;
    wire _1021;
    wire _1009;
    wire [63:0] _1006;
    wire [63:0] _1007;
    wire [62:0] _1008;
    wire [63:0] _1010;
    wire _1011;
    wire _1012;
    wire _1000;
    wire [63:0] _997;
    wire [63:0] _998;
    wire [62:0] _999;
    wire [63:0] _1001;
    wire _1002;
    wire _1003;
    wire _991;
    wire [63:0] _988;
    wire [63:0] _989;
    wire [62:0] _990;
    wire [63:0] _992;
    wire _993;
    wire _994;
    wire _982;
    wire [63:0] _979;
    wire [63:0] _980;
    wire [62:0] _981;
    wire [63:0] _983;
    wire _984;
    wire _985;
    wire _973;
    wire [63:0] _970;
    wire [63:0] _971;
    wire [62:0] _972;
    wire [63:0] _974;
    wire _975;
    wire _976;
    wire _964;
    wire [63:0] _961;
    wire [63:0] _962;
    wire [62:0] _963;
    wire [63:0] _965;
    wire _966;
    wire _967;
    wire _955;
    wire [63:0] _952;
    wire [63:0] _953;
    wire [62:0] _954;
    wire [63:0] _956;
    wire _957;
    wire _958;
    wire _946;
    wire [63:0] _943;
    wire [63:0] _944;
    wire [62:0] _945;
    wire [63:0] _947;
    wire _948;
    wire _949;
    wire _937;
    wire [63:0] _934;
    wire [63:0] _935;
    wire [62:0] _936;
    wire [63:0] _938;
    wire _939;
    wire _940;
    wire _928;
    wire [63:0] _925;
    wire [63:0] _926;
    wire [62:0] _927;
    wire [63:0] _929;
    wire _930;
    wire _931;
    wire _919;
    wire [63:0] _916;
    wire [63:0] _917;
    wire [62:0] _918;
    wire [63:0] _920;
    wire _921;
    wire _922;
    wire _910;
    wire [63:0] _907;
    wire [63:0] _908;
    wire [62:0] _909;
    wire [63:0] _911;
    wire _912;
    wire _913;
    wire _901;
    wire [63:0] _898;
    wire [63:0] _899;
    wire [62:0] _900;
    wire [63:0] _902;
    wire _903;
    wire _904;
    wire _892;
    wire [63:0] _889;
    wire [63:0] _890;
    wire [62:0] _891;
    wire [63:0] _893;
    wire _894;
    wire _895;
    wire _883;
    wire [63:0] _880;
    wire [63:0] _881;
    wire [62:0] _882;
    wire [63:0] _884;
    wire _885;
    wire _886;
    wire _874;
    wire [63:0] _871;
    wire [63:0] _872;
    wire [62:0] _873;
    wire [63:0] _875;
    wire _876;
    wire _877;
    wire _865;
    wire [63:0] _862;
    wire [63:0] _863;
    wire [62:0] _864;
    wire [63:0] _866;
    wire _867;
    wire _868;
    wire _856;
    wire [63:0] _853;
    wire [63:0] _854;
    wire [62:0] _855;
    wire [63:0] _857;
    wire _858;
    wire _859;
    wire _847;
    wire [63:0] _844;
    wire [63:0] _845;
    wire [62:0] _846;
    wire [63:0] _848;
    wire _849;
    wire _850;
    wire _838;
    wire [63:0] _835;
    wire [63:0] _836;
    wire [62:0] _837;
    wire [63:0] _839;
    wire _840;
    wire _841;
    wire _829;
    wire [63:0] _826;
    wire [63:0] _827;
    wire [62:0] _828;
    wire [63:0] _830;
    wire _831;
    wire _832;
    wire _820;
    wire [63:0] _817;
    wire [63:0] _818;
    wire [62:0] _819;
    wire [63:0] _821;
    wire _822;
    wire _823;
    wire _811;
    wire [63:0] _808;
    wire [63:0] _809;
    wire [62:0] _810;
    wire [63:0] _812;
    wire _813;
    wire _814;
    wire _802;
    wire [63:0] _799;
    wire [63:0] _800;
    wire [62:0] _801;
    wire [63:0] _803;
    wire _804;
    wire _805;
    wire _793;
    wire [63:0] _790;
    wire [63:0] _791;
    wire [62:0] _792;
    wire [63:0] _794;
    wire _795;
    wire _796;
    wire _784;
    wire [63:0] _781;
    wire [63:0] _782;
    wire [62:0] _783;
    wire [63:0] _785;
    wire _786;
    wire _787;
    wire [63:0] _774;
    wire _775;
    wire [63:0] _776;
    wire _777;
    wire _778;
    wire [63:0] _779;
    wire [62:0] _780;
    wire [63:0] _788;
    wire [62:0] _789;
    wire [63:0] _797;
    wire [62:0] _798;
    wire [63:0] _806;
    wire [62:0] _807;
    wire [63:0] _815;
    wire [62:0] _816;
    wire [63:0] _824;
    wire [62:0] _825;
    wire [63:0] _833;
    wire [62:0] _834;
    wire [63:0] _842;
    wire [62:0] _843;
    wire [63:0] _851;
    wire [62:0] _852;
    wire [63:0] _860;
    wire [62:0] _861;
    wire [63:0] _869;
    wire [62:0] _870;
    wire [63:0] _878;
    wire [62:0] _879;
    wire [63:0] _887;
    wire [62:0] _888;
    wire [63:0] _896;
    wire [62:0] _897;
    wire [63:0] _905;
    wire [62:0] _906;
    wire [63:0] _914;
    wire [62:0] _915;
    wire [63:0] _923;
    wire [62:0] _924;
    wire [63:0] _932;
    wire [62:0] _933;
    wire [63:0] _941;
    wire [62:0] _942;
    wire [63:0] _950;
    wire [62:0] _951;
    wire [63:0] _959;
    wire [62:0] _960;
    wire [63:0] _968;
    wire [62:0] _969;
    wire [63:0] _977;
    wire [62:0] _978;
    wire [63:0] _986;
    wire [62:0] _987;
    wire [63:0] _995;
    wire [62:0] _996;
    wire [63:0] _1004;
    wire [62:0] _1005;
    wire [63:0] _1013;
    wire [62:0] _1014;
    wire [63:0] _1022;
    wire [62:0] _1023;
    wire [63:0] _1031;
    wire [62:0] _1032;
    wire [63:0] _1040;
    wire [62:0] _1041;
    wire [63:0] _1049;
    wire [62:0] _1050;
    wire [63:0] _1058;
    wire [62:0] _1059;
    wire [63:0] _1067;
    wire [62:0] _1068;
    wire [63:0] _1076;
    wire [62:0] _1077;
    wire [63:0] _1085;
    wire [62:0] _1086;
    wire [63:0] _1094;
    wire [62:0] _1095;
    wire [63:0] _1103;
    wire [62:0] _1104;
    wire [63:0] _1112;
    wire [62:0] _1113;
    wire [63:0] _1121;
    wire [62:0] _1122;
    wire [63:0] _1130;
    wire [62:0] _1131;
    wire [63:0] _1139;
    wire [62:0] _1140;
    wire [63:0] _1148;
    wire [62:0] _1149;
    wire [63:0] _1157;
    wire [62:0] _1158;
    wire [63:0] _1166;
    wire [62:0] _1167;
    wire [63:0] _1175;
    wire [62:0] _1176;
    wire [63:0] _1184;
    wire [62:0] _1185;
    wire [63:0] _1193;
    wire [62:0] _1194;
    wire [63:0] _1202;
    wire [62:0] _1203;
    wire [63:0] _1211;
    wire [62:0] _1212;
    wire [63:0] _1220;
    wire [62:0] _1221;
    wire [63:0] _1229;
    wire [62:0] _1230;
    wire [63:0] _1238;
    wire [62:0] _1239;
    wire [63:0] _1247;
    wire [62:0] _1248;
    wire [63:0] _1256;
    wire [62:0] _1257;
    wire [63:0] _1265;
    wire [62:0] _1266;
    wire [63:0] _1274;
    wire [62:0] _1275;
    wire [63:0] _1283;
    wire [62:0] _1284;
    wire [63:0] _1292;
    wire [62:0] _1293;
    wire [63:0] _1301;
    wire [62:0] _1302;
    wire [63:0] _1310;
    wire [62:0] _1311;
    wire [63:0] _1319;
    wire [62:0] _1320;
    wire [63:0] _1328;
    wire [62:0] _1329;
    wire [63:0] _1337;
    wire [62:0] _1338;
    wire [63:0] _1346;
    wire [63:0] _1348;
    wire [127:0] _1349;
    wire [63:0] _1350;
    wire [63:0] _1932;
    wire _2010;
    wire _2011;
    wire _2012;
    wire _2013;
    wire _2014;
    wire _2016;
    wire _2018;
    wire _2020;
    wire _2022;
    wire _2024;
    wire _2026;
    wire _2028;
    wire _2030;
    wire _734;
    wire [63:0] _731;
    wire [63:0] _732;
    wire [62:0] _733;
    wire [63:0] _735;
    wire _736;
    wire _737;
    wire _725;
    wire [63:0] _722;
    wire [63:0] _723;
    wire [62:0] _724;
    wire [63:0] _726;
    wire _727;
    wire _728;
    wire _716;
    wire [63:0] _713;
    wire [63:0] _714;
    wire [62:0] _715;
    wire [63:0] _717;
    wire _718;
    wire _719;
    wire _707;
    wire [63:0] _704;
    wire [63:0] _705;
    wire [62:0] _706;
    wire [63:0] _708;
    wire _709;
    wire _710;
    wire _698;
    wire [63:0] _695;
    wire [63:0] _696;
    wire [62:0] _697;
    wire [63:0] _699;
    wire _700;
    wire _701;
    wire _689;
    wire [63:0] _686;
    wire [63:0] _687;
    wire [62:0] _688;
    wire [63:0] _690;
    wire _691;
    wire _692;
    wire _680;
    wire [63:0] _677;
    wire [63:0] _678;
    wire [62:0] _679;
    wire [63:0] _681;
    wire _682;
    wire _683;
    wire _671;
    wire [63:0] _668;
    wire [63:0] _669;
    wire [62:0] _670;
    wire [63:0] _672;
    wire _673;
    wire _674;
    wire _662;
    wire [63:0] _659;
    wire [63:0] _660;
    wire [62:0] _661;
    wire [63:0] _663;
    wire _664;
    wire _665;
    wire _653;
    wire [63:0] _650;
    wire [63:0] _651;
    wire [62:0] _652;
    wire [63:0] _654;
    wire _655;
    wire _656;
    wire _644;
    wire [63:0] _641;
    wire [63:0] _642;
    wire [62:0] _643;
    wire [63:0] _645;
    wire _646;
    wire _647;
    wire _635;
    wire [63:0] _632;
    wire [63:0] _633;
    wire [62:0] _634;
    wire [63:0] _636;
    wire _637;
    wire _638;
    wire _626;
    wire [63:0] _623;
    wire [63:0] _624;
    wire [62:0] _625;
    wire [63:0] _627;
    wire _628;
    wire _629;
    wire _617;
    wire [63:0] _614;
    wire [63:0] _615;
    wire [62:0] _616;
    wire [63:0] _618;
    wire _619;
    wire _620;
    wire _608;
    wire [63:0] _605;
    wire [63:0] _606;
    wire [62:0] _607;
    wire [63:0] _609;
    wire _610;
    wire _611;
    wire _599;
    wire [63:0] _596;
    wire [63:0] _597;
    wire [62:0] _598;
    wire [63:0] _600;
    wire _601;
    wire _602;
    wire _590;
    wire [63:0] _587;
    wire [63:0] _588;
    wire [62:0] _589;
    wire [63:0] _591;
    wire _592;
    wire _593;
    wire _581;
    wire [63:0] _578;
    wire [63:0] _579;
    wire [62:0] _580;
    wire [63:0] _582;
    wire _583;
    wire _584;
    wire _572;
    wire [63:0] _569;
    wire [63:0] _570;
    wire [62:0] _571;
    wire [63:0] _573;
    wire _574;
    wire _575;
    wire _563;
    wire [63:0] _560;
    wire [63:0] _561;
    wire [62:0] _562;
    wire [63:0] _564;
    wire _565;
    wire _566;
    wire _554;
    wire [63:0] _551;
    wire [63:0] _552;
    wire [62:0] _553;
    wire [63:0] _555;
    wire _556;
    wire _557;
    wire _545;
    wire [63:0] _542;
    wire [63:0] _543;
    wire [62:0] _544;
    wire [63:0] _546;
    wire _547;
    wire _548;
    wire _536;
    wire [63:0] _533;
    wire [63:0] _534;
    wire [62:0] _535;
    wire [63:0] _537;
    wire _538;
    wire _539;
    wire _527;
    wire [63:0] _524;
    wire [63:0] _525;
    wire [62:0] _526;
    wire [63:0] _528;
    wire _529;
    wire _530;
    wire _518;
    wire [63:0] _515;
    wire [63:0] _516;
    wire [62:0] _517;
    wire [63:0] _519;
    wire _520;
    wire _521;
    wire _509;
    wire [63:0] _506;
    wire [63:0] _507;
    wire [62:0] _508;
    wire [63:0] _510;
    wire _511;
    wire _512;
    wire _500;
    wire [63:0] _497;
    wire [63:0] _498;
    wire [62:0] _499;
    wire [63:0] _501;
    wire _502;
    wire _503;
    wire _491;
    wire [63:0] _488;
    wire [63:0] _489;
    wire [62:0] _490;
    wire [63:0] _492;
    wire _493;
    wire _494;
    wire _482;
    wire [63:0] _479;
    wire [63:0] _480;
    wire [62:0] _481;
    wire [63:0] _483;
    wire _484;
    wire _485;
    wire _473;
    wire [63:0] _470;
    wire [63:0] _471;
    wire [62:0] _472;
    wire [63:0] _474;
    wire _475;
    wire _476;
    wire _464;
    wire [63:0] _461;
    wire [63:0] _462;
    wire [62:0] _463;
    wire [63:0] _465;
    wire _466;
    wire _467;
    wire _455;
    wire [63:0] _452;
    wire [63:0] _453;
    wire [62:0] _454;
    wire [63:0] _456;
    wire _457;
    wire _458;
    wire _446;
    wire [63:0] _443;
    wire [63:0] _444;
    wire [62:0] _445;
    wire [63:0] _447;
    wire _448;
    wire _449;
    wire _437;
    wire [63:0] _434;
    wire [63:0] _435;
    wire [62:0] _436;
    wire [63:0] _438;
    wire _439;
    wire _440;
    wire _428;
    wire [63:0] _425;
    wire [63:0] _426;
    wire [62:0] _427;
    wire [63:0] _429;
    wire _430;
    wire _431;
    wire _419;
    wire [63:0] _416;
    wire [63:0] _417;
    wire [62:0] _418;
    wire [63:0] _420;
    wire _421;
    wire _422;
    wire _410;
    wire [63:0] _407;
    wire [63:0] _408;
    wire [62:0] _409;
    wire [63:0] _411;
    wire _412;
    wire _413;
    wire _401;
    wire [63:0] _398;
    wire [63:0] _399;
    wire [62:0] _400;
    wire [63:0] _402;
    wire _403;
    wire _404;
    wire _392;
    wire [63:0] _389;
    wire [63:0] _390;
    wire [62:0] _391;
    wire [63:0] _393;
    wire _394;
    wire _395;
    wire _383;
    wire [63:0] _380;
    wire [63:0] _381;
    wire [62:0] _382;
    wire [63:0] _384;
    wire _385;
    wire _386;
    wire _374;
    wire [63:0] _371;
    wire [63:0] _372;
    wire [62:0] _373;
    wire [63:0] _375;
    wire _376;
    wire _377;
    wire _365;
    wire [63:0] _362;
    wire [63:0] _363;
    wire [62:0] _364;
    wire [63:0] _366;
    wire _367;
    wire _368;
    wire _356;
    wire [63:0] _353;
    wire [63:0] _354;
    wire [62:0] _355;
    wire [63:0] _357;
    wire _358;
    wire _359;
    wire _347;
    wire [63:0] _344;
    wire [63:0] _345;
    wire [62:0] _346;
    wire [63:0] _348;
    wire _349;
    wire _350;
    wire _338;
    wire [63:0] _335;
    wire [63:0] _336;
    wire [62:0] _337;
    wire [63:0] _339;
    wire _340;
    wire _341;
    wire _329;
    wire [63:0] _326;
    wire [63:0] _327;
    wire [62:0] _328;
    wire [63:0] _330;
    wire _331;
    wire _332;
    wire _320;
    wire [63:0] _317;
    wire [63:0] _318;
    wire [62:0] _319;
    wire [63:0] _321;
    wire _322;
    wire _323;
    wire _311;
    wire [63:0] _308;
    wire [63:0] _309;
    wire [62:0] _310;
    wire [63:0] _312;
    wire _313;
    wire _314;
    wire _302;
    wire [63:0] _299;
    wire [63:0] _300;
    wire [62:0] _301;
    wire [63:0] _303;
    wire _304;
    wire _305;
    wire _293;
    wire [63:0] _290;
    wire [63:0] _291;
    wire [62:0] _292;
    wire [63:0] _294;
    wire _295;
    wire _296;
    wire _284;
    wire [63:0] _281;
    wire [63:0] _282;
    wire [62:0] _283;
    wire [63:0] _285;
    wire _286;
    wire _287;
    wire _275;
    wire [63:0] _272;
    wire [63:0] _273;
    wire [62:0] _274;
    wire [63:0] _276;
    wire _277;
    wire _278;
    wire _266;
    wire [63:0] _263;
    wire [63:0] _264;
    wire [62:0] _265;
    wire [63:0] _267;
    wire _268;
    wire _269;
    wire _257;
    wire [63:0] _254;
    wire [63:0] _255;
    wire [62:0] _256;
    wire [63:0] _258;
    wire _259;
    wire _260;
    wire _248;
    wire [63:0] _245;
    wire [63:0] _246;
    wire [62:0] _247;
    wire [63:0] _249;
    wire _250;
    wire _251;
    wire _239;
    wire [63:0] _236;
    wire [63:0] _237;
    wire [62:0] _238;
    wire [63:0] _240;
    wire _241;
    wire _242;
    wire _230;
    wire [63:0] _227;
    wire [63:0] _228;
    wire [62:0] _229;
    wire [63:0] _231;
    wire _232;
    wire _233;
    wire _221;
    wire [63:0] _218;
    wire [63:0] _219;
    wire [62:0] _220;
    wire [63:0] _222;
    wire _223;
    wire _224;
    wire _212;
    wire [63:0] _209;
    wire [63:0] _210;
    wire [62:0] _211;
    wire [63:0] _213;
    wire _214;
    wire _215;
    wire _203;
    wire [63:0] _200;
    wire [63:0] _201;
    wire [62:0] _202;
    wire [63:0] _204;
    wire _205;
    wire _206;
    wire _194;
    wire [63:0] _191;
    wire [63:0] _192;
    wire [62:0] _193;
    wire [63:0] _195;
    wire _196;
    wire _197;
    wire _185;
    wire [63:0] _182;
    wire [63:0] _183;
    wire [62:0] _184;
    wire [63:0] _186;
    wire _187;
    wire _188;
    wire _176;
    wire [63:0] _173;
    wire [63:0] _174;
    wire [62:0] _175;
    wire [63:0] _177;
    wire _178;
    wire _179;
    wire [63:0] _162;
    wire [63:0] _160;
    wire [63:0] _158;
    wire [63:0] _156;
    wire [63:0] _154;
    wire [63:0] _152;
    wire [63:0] _150;
    wire [63:0] _148;
    wire [63:0] _146;
    wire [63:0] _144;
    wire [63:0] _142;
    wire [63:0] _140;
    wire [63:0] _138;
    wire [63:0] _139;
    wire [63:0] _141;
    wire [63:0] _143;
    wire [63:0] _145;
    wire [63:0] _147;
    wire [63:0] _149;
    wire [63:0] _151;
    wire [63:0] _153;
    wire [63:0] _155;
    wire [63:0] _157;
    wire [63:0] _159;
    wire [63:0] _161;
    wire [63:0] _163;
    wire [63:0] _165;
    wire [63:0] _8;
    wire [63:0] _1977;
    wire [63:0] _1979;
    wire [63:0] _9;
    reg [63:0] _136;
    wire [63:0] _166;
    wire _167;
    wire [63:0] _168;
    wire _169;
    wire _170;
    wire [63:0] _171;
    wire [62:0] _172;
    wire [63:0] _180;
    wire [62:0] _181;
    wire [63:0] _189;
    wire [62:0] _190;
    wire [63:0] _198;
    wire [62:0] _199;
    wire [63:0] _207;
    wire [62:0] _208;
    wire [63:0] _216;
    wire [62:0] _217;
    wire [63:0] _225;
    wire [62:0] _226;
    wire [63:0] _234;
    wire [62:0] _235;
    wire [63:0] _243;
    wire [62:0] _244;
    wire [63:0] _252;
    wire [62:0] _253;
    wire [63:0] _261;
    wire [62:0] _262;
    wire [63:0] _270;
    wire [62:0] _271;
    wire [63:0] _279;
    wire [62:0] _280;
    wire [63:0] _288;
    wire [62:0] _289;
    wire [63:0] _297;
    wire [62:0] _298;
    wire [63:0] _306;
    wire [62:0] _307;
    wire [63:0] _315;
    wire [62:0] _316;
    wire [63:0] _324;
    wire [62:0] _325;
    wire [63:0] _333;
    wire [62:0] _334;
    wire [63:0] _342;
    wire [62:0] _343;
    wire [63:0] _351;
    wire [62:0] _352;
    wire [63:0] _360;
    wire [62:0] _361;
    wire [63:0] _369;
    wire [62:0] _370;
    wire [63:0] _378;
    wire [62:0] _379;
    wire [63:0] _387;
    wire [62:0] _388;
    wire [63:0] _396;
    wire [62:0] _397;
    wire [63:0] _405;
    wire [62:0] _406;
    wire [63:0] _414;
    wire [62:0] _415;
    wire [63:0] _423;
    wire [62:0] _424;
    wire [63:0] _432;
    wire [62:0] _433;
    wire [63:0] _441;
    wire [62:0] _442;
    wire [63:0] _450;
    wire [62:0] _451;
    wire [63:0] _459;
    wire [62:0] _460;
    wire [63:0] _468;
    wire [62:0] _469;
    wire [63:0] _477;
    wire [62:0] _478;
    wire [63:0] _486;
    wire [62:0] _487;
    wire [63:0] _495;
    wire [62:0] _496;
    wire [63:0] _504;
    wire [62:0] _505;
    wire [63:0] _513;
    wire [62:0] _514;
    wire [63:0] _522;
    wire [62:0] _523;
    wire [63:0] _531;
    wire [62:0] _532;
    wire [63:0] _540;
    wire [62:0] _541;
    wire [63:0] _549;
    wire [62:0] _550;
    wire [63:0] _558;
    wire [62:0] _559;
    wire [63:0] _567;
    wire [62:0] _568;
    wire [63:0] _576;
    wire [62:0] _577;
    wire [63:0] _585;
    wire [62:0] _586;
    wire [63:0] _594;
    wire [62:0] _595;
    wire [63:0] _603;
    wire [62:0] _604;
    wire [63:0] _612;
    wire [62:0] _613;
    wire [63:0] _621;
    wire [62:0] _622;
    wire [63:0] _630;
    wire [62:0] _631;
    wire [63:0] _639;
    wire [62:0] _640;
    wire [63:0] _648;
    wire [62:0] _649;
    wire [63:0] _657;
    wire [62:0] _658;
    wire [63:0] _666;
    wire [62:0] _667;
    wire [63:0] _675;
    wire [62:0] _676;
    wire [63:0] _684;
    wire [62:0] _685;
    wire [63:0] _693;
    wire [62:0] _694;
    wire [63:0] _702;
    wire [62:0] _703;
    wire [63:0] _711;
    wire [62:0] _712;
    wire [63:0] _720;
    wire [62:0] _721;
    wire [63:0] _729;
    wire [62:0] _730;
    wire [63:0] _738;
    wire [127:0] _739;
    wire [63:0] _740;
    wire [63:0] _126;
    wire [63:0] _124;
    wire [63:0] _120;
    wire [63:0] _114;
    wire [63:0] _112;
    wire [63:0] _110;
    wire [63:0] _108;
    wire [63:0] _107;
    wire [63:0] _109;
    wire [63:0] _111;
    wire [63:0] _113;
    wire [63:0] _115;
    wire [63:0] _117;
    wire [63:0] _119;
    wire [63:0] _121;
    wire [63:0] _123;
    wire [63:0] _125;
    wire [63:0] _127;
    wire [63:0] _129;
    wire [63:0] _131;
    wire _741;
    wire [63:0] _742;
    wire [63:0] _101;
    wire [63:0] _99;
    wire [63:0] _95;
    wire [63:0] _93;
    wire [63:0] _89;
    wire [63:0] _87;
    wire [63:0] _83;
    wire [63:0] _79;
    wire [63:0] _77;
    wire [3:0] _74;
    wire _75;
    wire [63:0] _78;
    wire [3:0] _72;
    wire _73;
    wire [63:0] _80;
    wire [3:0] _70;
    wire _71;
    wire [63:0] _82;
    wire [3:0] _68;
    wire _69;
    wire [63:0] _84;
    wire [3:0] _66;
    wire _67;
    wire [63:0] _86;
    wire [3:0] _64;
    wire _65;
    wire [63:0] _88;
    wire [3:0] _62;
    wire _63;
    wire [63:0] _90;
    wire [3:0] _60;
    wire _61;
    wire [63:0] _92;
    wire [3:0] _58;
    wire _59;
    wire [63:0] _94;
    wire [3:0] _56;
    wire _57;
    wire [63:0] _96;
    wire [3:0] _54;
    wire _55;
    wire [63:0] _98;
    wire [3:0] _52;
    wire _53;
    wire [63:0] _100;
    wire [3:0] _50;
    wire _51;
    wire [63:0] _102;
    wire [63:0] _11;
    wire [63:0] _1980;
    wire [63:0] _1982;
    wire [63:0] _12;
    reg [63:0] _49;
    wire _103;
    wire [63:0] _104;
    wire _743;
    wire _744;
    wire _2031;
    wire [63:0] _2033;
    wire [63:0] _2034;
    wire _2008;
    wire _2004;
    wire _14;
    wire _1986;
    wire _1988;
    wire _15;
    reg _1985;
    wire vdd;
    wire _17;
    wire _19;
    wire [3:0] _1990;
    wire [3:0] _1991;
    wire [3:0] _1993;
    wire [3:0] _1995;
    wire [3:0] _20;
    reg [3:0] _32;
    wire _1997;
    wire _1998;
    wire _1999;
    wire _2000;
    wire _2002;
    wire _21;
    reg _35;
    wire _40;
    wire _39;
    wire _41;
    wire _23;
    wire _1976;
    wire _2005;
    wire _2007;
    wire _24;
    reg _38;
    wire _2009;
    wire [63:0] _2035;
    wire _26;
    wire [63:0] _2037;
    wire [63:0] _27;
    reg [63:0] _1973;
    assign _45 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign _766 = 1'b0;
    assign _747 = _75 ? _766 : _766;
    assign _749 = _73 ? _766 : _747;
    assign _751 = _71 ? _766 : _749;
    assign _753 = _69 ? _766 : _751;
    assign _755 = _67 ? _766 : _753;
    assign _757 = _65 ? _766 : _755;
    assign _759 = _63 ? _766 : _757;
    assign _761 = _61 ? _766 : _759;
    assign _763 = _59 ? _766 : _761;
    assign _765 = _57 ? _766 : _763;
    assign _767 = _55 ? _766 : _765;
    assign _768 = _53 ? vdd : _767;
    assign _769 = _51 ? vdd : _768;
    assign _770 = _744 & _769;
    assign _1933 = _770 ? _1932 : _45;
    assign _1934 = _46 + _1933;
    assign _42 = ~ _35;
    assign _43 = _38 & _42;
    assign _1935 = _43 ? _1934 : _46;
    assign _1937 = _26 ? _45 : _1935;
    assign _4 = _1937;
    always @(posedge _19) begin
        if (_17)
            _46 <= _45;
        else
            _46 <= _4;
    end
    assign _1945 = _75 ? _766 : _766;
    assign _1947 = _73 ? _766 : _1945;
    assign _1949 = _71 ? _766 : _1947;
    assign _1951 = _69 ? _766 : _1949;
    assign _1953 = _67 ? _766 : _1951;
    assign _1954 = _65 ? vdd : _1953;
    assign _1955 = _63 ? vdd : _1954;
    assign _1956 = _61 ? vdd : _1955;
    assign _1957 = _59 ? vdd : _1956;
    assign _1958 = _57 ? vdd : _1957;
    assign _1959 = _55 ? vdd : _1958;
    assign _1961 = _53 ? _766 : _1959;
    assign _1963 = _51 ? _766 : _1961;
    assign _1964 = _744 & _1963;
    assign _1966 = _1964 ? _1932 : _45;
    assign _1967 = _1942 + _1966;
    assign _1938 = ~ _35;
    assign _1939 = _38 & _1938;
    assign _1968 = _1939 ? _1967 : _1942;
    assign _1970 = _26 ? _45 : _1968;
    assign _5 = _1970;
    always @(posedge _19) begin
        if (_17)
            _1942 <= _45;
        else
            _1942 <= _5;
    end
    assign _1974 = _1973 + _1942;
    assign _1975 = _1974 - _46;
    assign _1925 = _1356[0:0];
    assign _1922 = _1917 - _1359;
    assign _1923 = _1919 ? _1922 : _1917;
    assign _1924 = _1923[62:0];
    assign _1926 = { _1924,
                     _1925 };
    assign _1927 = _1926 < _1359;
    assign _1928 = ~ _1927;
    assign _1916 = _1356[1:1];
    assign _1913 = _1908 - _1359;
    assign _1914 = _1910 ? _1913 : _1908;
    assign _1915 = _1914[62:0];
    assign _1917 = { _1915,
                     _1916 };
    assign _1918 = _1917 < _1359;
    assign _1919 = ~ _1918;
    assign _1907 = _1356[2:2];
    assign _1904 = _1899 - _1359;
    assign _1905 = _1901 ? _1904 : _1899;
    assign _1906 = _1905[62:0];
    assign _1908 = { _1906,
                     _1907 };
    assign _1909 = _1908 < _1359;
    assign _1910 = ~ _1909;
    assign _1898 = _1356[3:3];
    assign _1895 = _1890 - _1359;
    assign _1896 = _1892 ? _1895 : _1890;
    assign _1897 = _1896[62:0];
    assign _1899 = { _1897,
                     _1898 };
    assign _1900 = _1899 < _1359;
    assign _1901 = ~ _1900;
    assign _1889 = _1356[4:4];
    assign _1886 = _1881 - _1359;
    assign _1887 = _1883 ? _1886 : _1881;
    assign _1888 = _1887[62:0];
    assign _1890 = { _1888,
                     _1889 };
    assign _1891 = _1890 < _1359;
    assign _1892 = ~ _1891;
    assign _1880 = _1356[5:5];
    assign _1877 = _1872 - _1359;
    assign _1878 = _1874 ? _1877 : _1872;
    assign _1879 = _1878[62:0];
    assign _1881 = { _1879,
                     _1880 };
    assign _1882 = _1881 < _1359;
    assign _1883 = ~ _1882;
    assign _1871 = _1356[6:6];
    assign _1868 = _1863 - _1359;
    assign _1869 = _1865 ? _1868 : _1863;
    assign _1870 = _1869[62:0];
    assign _1872 = { _1870,
                     _1871 };
    assign _1873 = _1872 < _1359;
    assign _1874 = ~ _1873;
    assign _1862 = _1356[7:7];
    assign _1859 = _1854 - _1359;
    assign _1860 = _1856 ? _1859 : _1854;
    assign _1861 = _1860[62:0];
    assign _1863 = { _1861,
                     _1862 };
    assign _1864 = _1863 < _1359;
    assign _1865 = ~ _1864;
    assign _1853 = _1356[8:8];
    assign _1850 = _1845 - _1359;
    assign _1851 = _1847 ? _1850 : _1845;
    assign _1852 = _1851[62:0];
    assign _1854 = { _1852,
                     _1853 };
    assign _1855 = _1854 < _1359;
    assign _1856 = ~ _1855;
    assign _1844 = _1356[9:9];
    assign _1841 = _1836 - _1359;
    assign _1842 = _1838 ? _1841 : _1836;
    assign _1843 = _1842[62:0];
    assign _1845 = { _1843,
                     _1844 };
    assign _1846 = _1845 < _1359;
    assign _1847 = ~ _1846;
    assign _1835 = _1356[10:10];
    assign _1832 = _1827 - _1359;
    assign _1833 = _1829 ? _1832 : _1827;
    assign _1834 = _1833[62:0];
    assign _1836 = { _1834,
                     _1835 };
    assign _1837 = _1836 < _1359;
    assign _1838 = ~ _1837;
    assign _1826 = _1356[11:11];
    assign _1823 = _1818 - _1359;
    assign _1824 = _1820 ? _1823 : _1818;
    assign _1825 = _1824[62:0];
    assign _1827 = { _1825,
                     _1826 };
    assign _1828 = _1827 < _1359;
    assign _1829 = ~ _1828;
    assign _1817 = _1356[12:12];
    assign _1814 = _1809 - _1359;
    assign _1815 = _1811 ? _1814 : _1809;
    assign _1816 = _1815[62:0];
    assign _1818 = { _1816,
                     _1817 };
    assign _1819 = _1818 < _1359;
    assign _1820 = ~ _1819;
    assign _1808 = _1356[13:13];
    assign _1805 = _1800 - _1359;
    assign _1806 = _1802 ? _1805 : _1800;
    assign _1807 = _1806[62:0];
    assign _1809 = { _1807,
                     _1808 };
    assign _1810 = _1809 < _1359;
    assign _1811 = ~ _1810;
    assign _1799 = _1356[14:14];
    assign _1796 = _1791 - _1359;
    assign _1797 = _1793 ? _1796 : _1791;
    assign _1798 = _1797[62:0];
    assign _1800 = { _1798,
                     _1799 };
    assign _1801 = _1800 < _1359;
    assign _1802 = ~ _1801;
    assign _1790 = _1356[15:15];
    assign _1787 = _1782 - _1359;
    assign _1788 = _1784 ? _1787 : _1782;
    assign _1789 = _1788[62:0];
    assign _1791 = { _1789,
                     _1790 };
    assign _1792 = _1791 < _1359;
    assign _1793 = ~ _1792;
    assign _1781 = _1356[16:16];
    assign _1778 = _1773 - _1359;
    assign _1779 = _1775 ? _1778 : _1773;
    assign _1780 = _1779[62:0];
    assign _1782 = { _1780,
                     _1781 };
    assign _1783 = _1782 < _1359;
    assign _1784 = ~ _1783;
    assign _1772 = _1356[17:17];
    assign _1769 = _1764 - _1359;
    assign _1770 = _1766 ? _1769 : _1764;
    assign _1771 = _1770[62:0];
    assign _1773 = { _1771,
                     _1772 };
    assign _1774 = _1773 < _1359;
    assign _1775 = ~ _1774;
    assign _1763 = _1356[18:18];
    assign _1760 = _1755 - _1359;
    assign _1761 = _1757 ? _1760 : _1755;
    assign _1762 = _1761[62:0];
    assign _1764 = { _1762,
                     _1763 };
    assign _1765 = _1764 < _1359;
    assign _1766 = ~ _1765;
    assign _1754 = _1356[19:19];
    assign _1751 = _1746 - _1359;
    assign _1752 = _1748 ? _1751 : _1746;
    assign _1753 = _1752[62:0];
    assign _1755 = { _1753,
                     _1754 };
    assign _1756 = _1755 < _1359;
    assign _1757 = ~ _1756;
    assign _1745 = _1356[20:20];
    assign _1742 = _1737 - _1359;
    assign _1743 = _1739 ? _1742 : _1737;
    assign _1744 = _1743[62:0];
    assign _1746 = { _1744,
                     _1745 };
    assign _1747 = _1746 < _1359;
    assign _1748 = ~ _1747;
    assign _1736 = _1356[21:21];
    assign _1733 = _1728 - _1359;
    assign _1734 = _1730 ? _1733 : _1728;
    assign _1735 = _1734[62:0];
    assign _1737 = { _1735,
                     _1736 };
    assign _1738 = _1737 < _1359;
    assign _1739 = ~ _1738;
    assign _1727 = _1356[22:22];
    assign _1724 = _1719 - _1359;
    assign _1725 = _1721 ? _1724 : _1719;
    assign _1726 = _1725[62:0];
    assign _1728 = { _1726,
                     _1727 };
    assign _1729 = _1728 < _1359;
    assign _1730 = ~ _1729;
    assign _1718 = _1356[23:23];
    assign _1715 = _1710 - _1359;
    assign _1716 = _1712 ? _1715 : _1710;
    assign _1717 = _1716[62:0];
    assign _1719 = { _1717,
                     _1718 };
    assign _1720 = _1719 < _1359;
    assign _1721 = ~ _1720;
    assign _1709 = _1356[24:24];
    assign _1706 = _1701 - _1359;
    assign _1707 = _1703 ? _1706 : _1701;
    assign _1708 = _1707[62:0];
    assign _1710 = { _1708,
                     _1709 };
    assign _1711 = _1710 < _1359;
    assign _1712 = ~ _1711;
    assign _1700 = _1356[25:25];
    assign _1697 = _1692 - _1359;
    assign _1698 = _1694 ? _1697 : _1692;
    assign _1699 = _1698[62:0];
    assign _1701 = { _1699,
                     _1700 };
    assign _1702 = _1701 < _1359;
    assign _1703 = ~ _1702;
    assign _1691 = _1356[26:26];
    assign _1688 = _1683 - _1359;
    assign _1689 = _1685 ? _1688 : _1683;
    assign _1690 = _1689[62:0];
    assign _1692 = { _1690,
                     _1691 };
    assign _1693 = _1692 < _1359;
    assign _1694 = ~ _1693;
    assign _1682 = _1356[27:27];
    assign _1679 = _1674 - _1359;
    assign _1680 = _1676 ? _1679 : _1674;
    assign _1681 = _1680[62:0];
    assign _1683 = { _1681,
                     _1682 };
    assign _1684 = _1683 < _1359;
    assign _1685 = ~ _1684;
    assign _1673 = _1356[28:28];
    assign _1670 = _1665 - _1359;
    assign _1671 = _1667 ? _1670 : _1665;
    assign _1672 = _1671[62:0];
    assign _1674 = { _1672,
                     _1673 };
    assign _1675 = _1674 < _1359;
    assign _1676 = ~ _1675;
    assign _1664 = _1356[29:29];
    assign _1661 = _1656 - _1359;
    assign _1662 = _1658 ? _1661 : _1656;
    assign _1663 = _1662[62:0];
    assign _1665 = { _1663,
                     _1664 };
    assign _1666 = _1665 < _1359;
    assign _1667 = ~ _1666;
    assign _1655 = _1356[30:30];
    assign _1652 = _1647 - _1359;
    assign _1653 = _1649 ? _1652 : _1647;
    assign _1654 = _1653[62:0];
    assign _1656 = { _1654,
                     _1655 };
    assign _1657 = _1656 < _1359;
    assign _1658 = ~ _1657;
    assign _1646 = _1356[31:31];
    assign _1643 = _1638 - _1359;
    assign _1644 = _1640 ? _1643 : _1638;
    assign _1645 = _1644[62:0];
    assign _1647 = { _1645,
                     _1646 };
    assign _1648 = _1647 < _1359;
    assign _1649 = ~ _1648;
    assign _1637 = _1356[32:32];
    assign _1634 = _1629 - _1359;
    assign _1635 = _1631 ? _1634 : _1629;
    assign _1636 = _1635[62:0];
    assign _1638 = { _1636,
                     _1637 };
    assign _1639 = _1638 < _1359;
    assign _1640 = ~ _1639;
    assign _1628 = _1356[33:33];
    assign _1625 = _1620 - _1359;
    assign _1626 = _1622 ? _1625 : _1620;
    assign _1627 = _1626[62:0];
    assign _1629 = { _1627,
                     _1628 };
    assign _1630 = _1629 < _1359;
    assign _1631 = ~ _1630;
    assign _1619 = _1356[34:34];
    assign _1616 = _1611 - _1359;
    assign _1617 = _1613 ? _1616 : _1611;
    assign _1618 = _1617[62:0];
    assign _1620 = { _1618,
                     _1619 };
    assign _1621 = _1620 < _1359;
    assign _1622 = ~ _1621;
    assign _1610 = _1356[35:35];
    assign _1607 = _1602 - _1359;
    assign _1608 = _1604 ? _1607 : _1602;
    assign _1609 = _1608[62:0];
    assign _1611 = { _1609,
                     _1610 };
    assign _1612 = _1611 < _1359;
    assign _1613 = ~ _1612;
    assign _1601 = _1356[36:36];
    assign _1598 = _1593 - _1359;
    assign _1599 = _1595 ? _1598 : _1593;
    assign _1600 = _1599[62:0];
    assign _1602 = { _1600,
                     _1601 };
    assign _1603 = _1602 < _1359;
    assign _1604 = ~ _1603;
    assign _1592 = _1356[37:37];
    assign _1589 = _1584 - _1359;
    assign _1590 = _1586 ? _1589 : _1584;
    assign _1591 = _1590[62:0];
    assign _1593 = { _1591,
                     _1592 };
    assign _1594 = _1593 < _1359;
    assign _1595 = ~ _1594;
    assign _1583 = _1356[38:38];
    assign _1580 = _1575 - _1359;
    assign _1581 = _1577 ? _1580 : _1575;
    assign _1582 = _1581[62:0];
    assign _1584 = { _1582,
                     _1583 };
    assign _1585 = _1584 < _1359;
    assign _1586 = ~ _1585;
    assign _1574 = _1356[39:39];
    assign _1571 = _1566 - _1359;
    assign _1572 = _1568 ? _1571 : _1566;
    assign _1573 = _1572[62:0];
    assign _1575 = { _1573,
                     _1574 };
    assign _1576 = _1575 < _1359;
    assign _1577 = ~ _1576;
    assign _1565 = _1356[40:40];
    assign _1562 = _1557 - _1359;
    assign _1563 = _1559 ? _1562 : _1557;
    assign _1564 = _1563[62:0];
    assign _1566 = { _1564,
                     _1565 };
    assign _1567 = _1566 < _1359;
    assign _1568 = ~ _1567;
    assign _1556 = _1356[41:41];
    assign _1553 = _1548 - _1359;
    assign _1554 = _1550 ? _1553 : _1548;
    assign _1555 = _1554[62:0];
    assign _1557 = { _1555,
                     _1556 };
    assign _1558 = _1557 < _1359;
    assign _1559 = ~ _1558;
    assign _1547 = _1356[42:42];
    assign _1544 = _1539 - _1359;
    assign _1545 = _1541 ? _1544 : _1539;
    assign _1546 = _1545[62:0];
    assign _1548 = { _1546,
                     _1547 };
    assign _1549 = _1548 < _1359;
    assign _1550 = ~ _1549;
    assign _1538 = _1356[43:43];
    assign _1535 = _1530 - _1359;
    assign _1536 = _1532 ? _1535 : _1530;
    assign _1537 = _1536[62:0];
    assign _1539 = { _1537,
                     _1538 };
    assign _1540 = _1539 < _1359;
    assign _1541 = ~ _1540;
    assign _1529 = _1356[44:44];
    assign _1526 = _1521 - _1359;
    assign _1527 = _1523 ? _1526 : _1521;
    assign _1528 = _1527[62:0];
    assign _1530 = { _1528,
                     _1529 };
    assign _1531 = _1530 < _1359;
    assign _1532 = ~ _1531;
    assign _1520 = _1356[45:45];
    assign _1517 = _1512 - _1359;
    assign _1518 = _1514 ? _1517 : _1512;
    assign _1519 = _1518[62:0];
    assign _1521 = { _1519,
                     _1520 };
    assign _1522 = _1521 < _1359;
    assign _1523 = ~ _1522;
    assign _1511 = _1356[46:46];
    assign _1508 = _1503 - _1359;
    assign _1509 = _1505 ? _1508 : _1503;
    assign _1510 = _1509[62:0];
    assign _1512 = { _1510,
                     _1511 };
    assign _1513 = _1512 < _1359;
    assign _1514 = ~ _1513;
    assign _1502 = _1356[47:47];
    assign _1499 = _1494 - _1359;
    assign _1500 = _1496 ? _1499 : _1494;
    assign _1501 = _1500[62:0];
    assign _1503 = { _1501,
                     _1502 };
    assign _1504 = _1503 < _1359;
    assign _1505 = ~ _1504;
    assign _1493 = _1356[48:48];
    assign _1490 = _1485 - _1359;
    assign _1491 = _1487 ? _1490 : _1485;
    assign _1492 = _1491[62:0];
    assign _1494 = { _1492,
                     _1493 };
    assign _1495 = _1494 < _1359;
    assign _1496 = ~ _1495;
    assign _1484 = _1356[49:49];
    assign _1481 = _1476 - _1359;
    assign _1482 = _1478 ? _1481 : _1476;
    assign _1483 = _1482[62:0];
    assign _1485 = { _1483,
                     _1484 };
    assign _1486 = _1485 < _1359;
    assign _1487 = ~ _1486;
    assign _1475 = _1356[50:50];
    assign _1472 = _1467 - _1359;
    assign _1473 = _1469 ? _1472 : _1467;
    assign _1474 = _1473[62:0];
    assign _1476 = { _1474,
                     _1475 };
    assign _1477 = _1476 < _1359;
    assign _1478 = ~ _1477;
    assign _1466 = _1356[51:51];
    assign _1463 = _1458 - _1359;
    assign _1464 = _1460 ? _1463 : _1458;
    assign _1465 = _1464[62:0];
    assign _1467 = { _1465,
                     _1466 };
    assign _1468 = _1467 < _1359;
    assign _1469 = ~ _1468;
    assign _1457 = _1356[52:52];
    assign _1454 = _1449 - _1359;
    assign _1455 = _1451 ? _1454 : _1449;
    assign _1456 = _1455[62:0];
    assign _1458 = { _1456,
                     _1457 };
    assign _1459 = _1458 < _1359;
    assign _1460 = ~ _1459;
    assign _1448 = _1356[53:53];
    assign _1445 = _1440 - _1359;
    assign _1446 = _1442 ? _1445 : _1440;
    assign _1447 = _1446[62:0];
    assign _1449 = { _1447,
                     _1448 };
    assign _1450 = _1449 < _1359;
    assign _1451 = ~ _1450;
    assign _1439 = _1356[54:54];
    assign _1436 = _1431 - _1359;
    assign _1437 = _1433 ? _1436 : _1431;
    assign _1438 = _1437[62:0];
    assign _1440 = { _1438,
                     _1439 };
    assign _1441 = _1440 < _1359;
    assign _1442 = ~ _1441;
    assign _1430 = _1356[55:55];
    assign _1427 = _1422 - _1359;
    assign _1428 = _1424 ? _1427 : _1422;
    assign _1429 = _1428[62:0];
    assign _1431 = { _1429,
                     _1430 };
    assign _1432 = _1431 < _1359;
    assign _1433 = ~ _1432;
    assign _1421 = _1356[56:56];
    assign _1418 = _1413 - _1359;
    assign _1419 = _1415 ? _1418 : _1413;
    assign _1420 = _1419[62:0];
    assign _1422 = { _1420,
                     _1421 };
    assign _1423 = _1422 < _1359;
    assign _1424 = ~ _1423;
    assign _1412 = _1356[57:57];
    assign _1409 = _1404 - _1359;
    assign _1410 = _1406 ? _1409 : _1404;
    assign _1411 = _1410[62:0];
    assign _1413 = { _1411,
                     _1412 };
    assign _1414 = _1413 < _1359;
    assign _1415 = ~ _1414;
    assign _1403 = _1356[58:58];
    assign _1400 = _1395 - _1359;
    assign _1401 = _1397 ? _1400 : _1395;
    assign _1402 = _1401[62:0];
    assign _1404 = { _1402,
                     _1403 };
    assign _1405 = _1404 < _1359;
    assign _1406 = ~ _1405;
    assign _1394 = _1356[59:59];
    assign _1391 = _1386 - _1359;
    assign _1392 = _1388 ? _1391 : _1386;
    assign _1393 = _1392[62:0];
    assign _1395 = { _1393,
                     _1394 };
    assign _1396 = _1395 < _1359;
    assign _1397 = ~ _1396;
    assign _1385 = _1356[60:60];
    assign _1382 = _1377 - _1359;
    assign _1383 = _1379 ? _1382 : _1377;
    assign _1384 = _1383[62:0];
    assign _1386 = { _1384,
                     _1385 };
    assign _1387 = _1386 < _1359;
    assign _1388 = ~ _1387;
    assign _1376 = _1356[61:61];
    assign _1373 = _1368 - _1359;
    assign _1374 = _1370 ? _1373 : _1368;
    assign _1375 = _1374[62:0];
    assign _1377 = { _1375,
                     _1376 };
    assign _1378 = _1377 < _1359;
    assign _1379 = ~ _1378;
    assign _1367 = _1356[62:62];
    assign _1364 = _1358 - _1359;
    assign _1365 = _1361 ? _1364 : _1358;
    assign _1366 = _1365[62:0];
    assign _1368 = { _1366,
                     _1367 };
    assign _1369 = _1368 < _1359;
    assign _1370 = ~ _1369;
    assign _1359 = 64'b0000000000000000000000000000000000000000000000000000000000000010;
    assign _1353 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    assign _1354 = _1346 + _1353;
    assign _1355 = _1346 * _1354;
    assign _1356 = _1355[63:0];
    assign _1357 = _1356[63:63];
    assign _1352 = 63'b000000000000000000000000000000000000000000000000000000000000000;
    assign _1358 = { _1352,
                     _1357 };
    assign _1360 = _1358 < _1359;
    assign _1361 = ~ _1360;
    assign _1362 = { _1352,
                     _1361 };
    assign _1363 = _1362[62:0];
    assign _1371 = { _1363,
                     _1370 };
    assign _1372 = _1371[62:0];
    assign _1380 = { _1372,
                     _1379 };
    assign _1381 = _1380[62:0];
    assign _1389 = { _1381,
                     _1388 };
    assign _1390 = _1389[62:0];
    assign _1398 = { _1390,
                     _1397 };
    assign _1399 = _1398[62:0];
    assign _1407 = { _1399,
                     _1406 };
    assign _1408 = _1407[62:0];
    assign _1416 = { _1408,
                     _1415 };
    assign _1417 = _1416[62:0];
    assign _1425 = { _1417,
                     _1424 };
    assign _1426 = _1425[62:0];
    assign _1434 = { _1426,
                     _1433 };
    assign _1435 = _1434[62:0];
    assign _1443 = { _1435,
                     _1442 };
    assign _1444 = _1443[62:0];
    assign _1452 = { _1444,
                     _1451 };
    assign _1453 = _1452[62:0];
    assign _1461 = { _1453,
                     _1460 };
    assign _1462 = _1461[62:0];
    assign _1470 = { _1462,
                     _1469 };
    assign _1471 = _1470[62:0];
    assign _1479 = { _1471,
                     _1478 };
    assign _1480 = _1479[62:0];
    assign _1488 = { _1480,
                     _1487 };
    assign _1489 = _1488[62:0];
    assign _1497 = { _1489,
                     _1496 };
    assign _1498 = _1497[62:0];
    assign _1506 = { _1498,
                     _1505 };
    assign _1507 = _1506[62:0];
    assign _1515 = { _1507,
                     _1514 };
    assign _1516 = _1515[62:0];
    assign _1524 = { _1516,
                     _1523 };
    assign _1525 = _1524[62:0];
    assign _1533 = { _1525,
                     _1532 };
    assign _1534 = _1533[62:0];
    assign _1542 = { _1534,
                     _1541 };
    assign _1543 = _1542[62:0];
    assign _1551 = { _1543,
                     _1550 };
    assign _1552 = _1551[62:0];
    assign _1560 = { _1552,
                     _1559 };
    assign _1561 = _1560[62:0];
    assign _1569 = { _1561,
                     _1568 };
    assign _1570 = _1569[62:0];
    assign _1578 = { _1570,
                     _1577 };
    assign _1579 = _1578[62:0];
    assign _1587 = { _1579,
                     _1586 };
    assign _1588 = _1587[62:0];
    assign _1596 = { _1588,
                     _1595 };
    assign _1597 = _1596[62:0];
    assign _1605 = { _1597,
                     _1604 };
    assign _1606 = _1605[62:0];
    assign _1614 = { _1606,
                     _1613 };
    assign _1615 = _1614[62:0];
    assign _1623 = { _1615,
                     _1622 };
    assign _1624 = _1623[62:0];
    assign _1632 = { _1624,
                     _1631 };
    assign _1633 = _1632[62:0];
    assign _1641 = { _1633,
                     _1640 };
    assign _1642 = _1641[62:0];
    assign _1650 = { _1642,
                     _1649 };
    assign _1651 = _1650[62:0];
    assign _1659 = { _1651,
                     _1658 };
    assign _1660 = _1659[62:0];
    assign _1668 = { _1660,
                     _1667 };
    assign _1669 = _1668[62:0];
    assign _1677 = { _1669,
                     _1676 };
    assign _1678 = _1677[62:0];
    assign _1686 = { _1678,
                     _1685 };
    assign _1687 = _1686[62:0];
    assign _1695 = { _1687,
                     _1694 };
    assign _1696 = _1695[62:0];
    assign _1704 = { _1696,
                     _1703 };
    assign _1705 = _1704[62:0];
    assign _1713 = { _1705,
                     _1712 };
    assign _1714 = _1713[62:0];
    assign _1722 = { _1714,
                     _1721 };
    assign _1723 = _1722[62:0];
    assign _1731 = { _1723,
                     _1730 };
    assign _1732 = _1731[62:0];
    assign _1740 = { _1732,
                     _1739 };
    assign _1741 = _1740[62:0];
    assign _1749 = { _1741,
                     _1748 };
    assign _1750 = _1749[62:0];
    assign _1758 = { _1750,
                     _1757 };
    assign _1759 = _1758[62:0];
    assign _1767 = { _1759,
                     _1766 };
    assign _1768 = _1767[62:0];
    assign _1776 = { _1768,
                     _1775 };
    assign _1777 = _1776[62:0];
    assign _1785 = { _1777,
                     _1784 };
    assign _1786 = _1785[62:0];
    assign _1794 = { _1786,
                     _1793 };
    assign _1795 = _1794[62:0];
    assign _1803 = { _1795,
                     _1802 };
    assign _1804 = _1803[62:0];
    assign _1812 = { _1804,
                     _1811 };
    assign _1813 = _1812[62:0];
    assign _1821 = { _1813,
                     _1820 };
    assign _1822 = _1821[62:0];
    assign _1830 = { _1822,
                     _1829 };
    assign _1831 = _1830[62:0];
    assign _1839 = { _1831,
                     _1838 };
    assign _1840 = _1839[62:0];
    assign _1848 = { _1840,
                     _1847 };
    assign _1849 = _1848[62:0];
    assign _1857 = { _1849,
                     _1856 };
    assign _1858 = _1857[62:0];
    assign _1866 = { _1858,
                     _1865 };
    assign _1867 = _1866[62:0];
    assign _1875 = { _1867,
                     _1874 };
    assign _1876 = _1875[62:0];
    assign _1884 = { _1876,
                     _1883 };
    assign _1885 = _1884[62:0];
    assign _1893 = { _1885,
                     _1892 };
    assign _1894 = _1893[62:0];
    assign _1902 = { _1894,
                     _1901 };
    assign _1903 = _1902[62:0];
    assign _1911 = { _1903,
                     _1910 };
    assign _1912 = _1911[62:0];
    assign _1920 = { _1912,
                     _1919 };
    assign _1921 = _1920[62:0];
    assign _1929 = { _1921,
                     _1928 };
    assign _1930 = _163 * _1929;
    assign _1931 = _1930[63:0];
    assign _1342 = _774[0:0];
    assign _1339 = _1334 - _163;
    assign _1340 = _1336 ? _1339 : _1334;
    assign _1341 = _1340[62:0];
    assign _1343 = { _1341,
                     _1342 };
    assign _1344 = _1343 < _163;
    assign _1345 = ~ _1344;
    assign _1333 = _774[1:1];
    assign _1330 = _1325 - _163;
    assign _1331 = _1327 ? _1330 : _1325;
    assign _1332 = _1331[62:0];
    assign _1334 = { _1332,
                     _1333 };
    assign _1335 = _1334 < _163;
    assign _1336 = ~ _1335;
    assign _1324 = _774[2:2];
    assign _1321 = _1316 - _163;
    assign _1322 = _1318 ? _1321 : _1316;
    assign _1323 = _1322[62:0];
    assign _1325 = { _1323,
                     _1324 };
    assign _1326 = _1325 < _163;
    assign _1327 = ~ _1326;
    assign _1315 = _774[3:3];
    assign _1312 = _1307 - _163;
    assign _1313 = _1309 ? _1312 : _1307;
    assign _1314 = _1313[62:0];
    assign _1316 = { _1314,
                     _1315 };
    assign _1317 = _1316 < _163;
    assign _1318 = ~ _1317;
    assign _1306 = _774[4:4];
    assign _1303 = _1298 - _163;
    assign _1304 = _1300 ? _1303 : _1298;
    assign _1305 = _1304[62:0];
    assign _1307 = { _1305,
                     _1306 };
    assign _1308 = _1307 < _163;
    assign _1309 = ~ _1308;
    assign _1297 = _774[5:5];
    assign _1294 = _1289 - _163;
    assign _1295 = _1291 ? _1294 : _1289;
    assign _1296 = _1295[62:0];
    assign _1298 = { _1296,
                     _1297 };
    assign _1299 = _1298 < _163;
    assign _1300 = ~ _1299;
    assign _1288 = _774[6:6];
    assign _1285 = _1280 - _163;
    assign _1286 = _1282 ? _1285 : _1280;
    assign _1287 = _1286[62:0];
    assign _1289 = { _1287,
                     _1288 };
    assign _1290 = _1289 < _163;
    assign _1291 = ~ _1290;
    assign _1279 = _774[7:7];
    assign _1276 = _1271 - _163;
    assign _1277 = _1273 ? _1276 : _1271;
    assign _1278 = _1277[62:0];
    assign _1280 = { _1278,
                     _1279 };
    assign _1281 = _1280 < _163;
    assign _1282 = ~ _1281;
    assign _1270 = _774[8:8];
    assign _1267 = _1262 - _163;
    assign _1268 = _1264 ? _1267 : _1262;
    assign _1269 = _1268[62:0];
    assign _1271 = { _1269,
                     _1270 };
    assign _1272 = _1271 < _163;
    assign _1273 = ~ _1272;
    assign _1261 = _774[9:9];
    assign _1258 = _1253 - _163;
    assign _1259 = _1255 ? _1258 : _1253;
    assign _1260 = _1259[62:0];
    assign _1262 = { _1260,
                     _1261 };
    assign _1263 = _1262 < _163;
    assign _1264 = ~ _1263;
    assign _1252 = _774[10:10];
    assign _1249 = _1244 - _163;
    assign _1250 = _1246 ? _1249 : _1244;
    assign _1251 = _1250[62:0];
    assign _1253 = { _1251,
                     _1252 };
    assign _1254 = _1253 < _163;
    assign _1255 = ~ _1254;
    assign _1243 = _774[11:11];
    assign _1240 = _1235 - _163;
    assign _1241 = _1237 ? _1240 : _1235;
    assign _1242 = _1241[62:0];
    assign _1244 = { _1242,
                     _1243 };
    assign _1245 = _1244 < _163;
    assign _1246 = ~ _1245;
    assign _1234 = _774[12:12];
    assign _1231 = _1226 - _163;
    assign _1232 = _1228 ? _1231 : _1226;
    assign _1233 = _1232[62:0];
    assign _1235 = { _1233,
                     _1234 };
    assign _1236 = _1235 < _163;
    assign _1237 = ~ _1236;
    assign _1225 = _774[13:13];
    assign _1222 = _1217 - _163;
    assign _1223 = _1219 ? _1222 : _1217;
    assign _1224 = _1223[62:0];
    assign _1226 = { _1224,
                     _1225 };
    assign _1227 = _1226 < _163;
    assign _1228 = ~ _1227;
    assign _1216 = _774[14:14];
    assign _1213 = _1208 - _163;
    assign _1214 = _1210 ? _1213 : _1208;
    assign _1215 = _1214[62:0];
    assign _1217 = { _1215,
                     _1216 };
    assign _1218 = _1217 < _163;
    assign _1219 = ~ _1218;
    assign _1207 = _774[15:15];
    assign _1204 = _1199 - _163;
    assign _1205 = _1201 ? _1204 : _1199;
    assign _1206 = _1205[62:0];
    assign _1208 = { _1206,
                     _1207 };
    assign _1209 = _1208 < _163;
    assign _1210 = ~ _1209;
    assign _1198 = _774[16:16];
    assign _1195 = _1190 - _163;
    assign _1196 = _1192 ? _1195 : _1190;
    assign _1197 = _1196[62:0];
    assign _1199 = { _1197,
                     _1198 };
    assign _1200 = _1199 < _163;
    assign _1201 = ~ _1200;
    assign _1189 = _774[17:17];
    assign _1186 = _1181 - _163;
    assign _1187 = _1183 ? _1186 : _1181;
    assign _1188 = _1187[62:0];
    assign _1190 = { _1188,
                     _1189 };
    assign _1191 = _1190 < _163;
    assign _1192 = ~ _1191;
    assign _1180 = _774[18:18];
    assign _1177 = _1172 - _163;
    assign _1178 = _1174 ? _1177 : _1172;
    assign _1179 = _1178[62:0];
    assign _1181 = { _1179,
                     _1180 };
    assign _1182 = _1181 < _163;
    assign _1183 = ~ _1182;
    assign _1171 = _774[19:19];
    assign _1168 = _1163 - _163;
    assign _1169 = _1165 ? _1168 : _1163;
    assign _1170 = _1169[62:0];
    assign _1172 = { _1170,
                     _1171 };
    assign _1173 = _1172 < _163;
    assign _1174 = ~ _1173;
    assign _1162 = _774[20:20];
    assign _1159 = _1154 - _163;
    assign _1160 = _1156 ? _1159 : _1154;
    assign _1161 = _1160[62:0];
    assign _1163 = { _1161,
                     _1162 };
    assign _1164 = _1163 < _163;
    assign _1165 = ~ _1164;
    assign _1153 = _774[21:21];
    assign _1150 = _1145 - _163;
    assign _1151 = _1147 ? _1150 : _1145;
    assign _1152 = _1151[62:0];
    assign _1154 = { _1152,
                     _1153 };
    assign _1155 = _1154 < _163;
    assign _1156 = ~ _1155;
    assign _1144 = _774[22:22];
    assign _1141 = _1136 - _163;
    assign _1142 = _1138 ? _1141 : _1136;
    assign _1143 = _1142[62:0];
    assign _1145 = { _1143,
                     _1144 };
    assign _1146 = _1145 < _163;
    assign _1147 = ~ _1146;
    assign _1135 = _774[23:23];
    assign _1132 = _1127 - _163;
    assign _1133 = _1129 ? _1132 : _1127;
    assign _1134 = _1133[62:0];
    assign _1136 = { _1134,
                     _1135 };
    assign _1137 = _1136 < _163;
    assign _1138 = ~ _1137;
    assign _1126 = _774[24:24];
    assign _1123 = _1118 - _163;
    assign _1124 = _1120 ? _1123 : _1118;
    assign _1125 = _1124[62:0];
    assign _1127 = { _1125,
                     _1126 };
    assign _1128 = _1127 < _163;
    assign _1129 = ~ _1128;
    assign _1117 = _774[25:25];
    assign _1114 = _1109 - _163;
    assign _1115 = _1111 ? _1114 : _1109;
    assign _1116 = _1115[62:0];
    assign _1118 = { _1116,
                     _1117 };
    assign _1119 = _1118 < _163;
    assign _1120 = ~ _1119;
    assign _1108 = _774[26:26];
    assign _1105 = _1100 - _163;
    assign _1106 = _1102 ? _1105 : _1100;
    assign _1107 = _1106[62:0];
    assign _1109 = { _1107,
                     _1108 };
    assign _1110 = _1109 < _163;
    assign _1111 = ~ _1110;
    assign _1099 = _774[27:27];
    assign _1096 = _1091 - _163;
    assign _1097 = _1093 ? _1096 : _1091;
    assign _1098 = _1097[62:0];
    assign _1100 = { _1098,
                     _1099 };
    assign _1101 = _1100 < _163;
    assign _1102 = ~ _1101;
    assign _1090 = _774[28:28];
    assign _1087 = _1082 - _163;
    assign _1088 = _1084 ? _1087 : _1082;
    assign _1089 = _1088[62:0];
    assign _1091 = { _1089,
                     _1090 };
    assign _1092 = _1091 < _163;
    assign _1093 = ~ _1092;
    assign _1081 = _774[29:29];
    assign _1078 = _1073 - _163;
    assign _1079 = _1075 ? _1078 : _1073;
    assign _1080 = _1079[62:0];
    assign _1082 = { _1080,
                     _1081 };
    assign _1083 = _1082 < _163;
    assign _1084 = ~ _1083;
    assign _1072 = _774[30:30];
    assign _1069 = _1064 - _163;
    assign _1070 = _1066 ? _1069 : _1064;
    assign _1071 = _1070[62:0];
    assign _1073 = { _1071,
                     _1072 };
    assign _1074 = _1073 < _163;
    assign _1075 = ~ _1074;
    assign _1063 = _774[31:31];
    assign _1060 = _1055 - _163;
    assign _1061 = _1057 ? _1060 : _1055;
    assign _1062 = _1061[62:0];
    assign _1064 = { _1062,
                     _1063 };
    assign _1065 = _1064 < _163;
    assign _1066 = ~ _1065;
    assign _1054 = _774[32:32];
    assign _1051 = _1046 - _163;
    assign _1052 = _1048 ? _1051 : _1046;
    assign _1053 = _1052[62:0];
    assign _1055 = { _1053,
                     _1054 };
    assign _1056 = _1055 < _163;
    assign _1057 = ~ _1056;
    assign _1045 = _774[33:33];
    assign _1042 = _1037 - _163;
    assign _1043 = _1039 ? _1042 : _1037;
    assign _1044 = _1043[62:0];
    assign _1046 = { _1044,
                     _1045 };
    assign _1047 = _1046 < _163;
    assign _1048 = ~ _1047;
    assign _1036 = _774[34:34];
    assign _1033 = _1028 - _163;
    assign _1034 = _1030 ? _1033 : _1028;
    assign _1035 = _1034[62:0];
    assign _1037 = { _1035,
                     _1036 };
    assign _1038 = _1037 < _163;
    assign _1039 = ~ _1038;
    assign _1027 = _774[35:35];
    assign _1024 = _1019 - _163;
    assign _1025 = _1021 ? _1024 : _1019;
    assign _1026 = _1025[62:0];
    assign _1028 = { _1026,
                     _1027 };
    assign _1029 = _1028 < _163;
    assign _1030 = ~ _1029;
    assign _1018 = _774[36:36];
    assign _1015 = _1010 - _163;
    assign _1016 = _1012 ? _1015 : _1010;
    assign _1017 = _1016[62:0];
    assign _1019 = { _1017,
                     _1018 };
    assign _1020 = _1019 < _163;
    assign _1021 = ~ _1020;
    assign _1009 = _774[37:37];
    assign _1006 = _1001 - _163;
    assign _1007 = _1003 ? _1006 : _1001;
    assign _1008 = _1007[62:0];
    assign _1010 = { _1008,
                     _1009 };
    assign _1011 = _1010 < _163;
    assign _1012 = ~ _1011;
    assign _1000 = _774[38:38];
    assign _997 = _992 - _163;
    assign _998 = _994 ? _997 : _992;
    assign _999 = _998[62:0];
    assign _1001 = { _999,
                     _1000 };
    assign _1002 = _1001 < _163;
    assign _1003 = ~ _1002;
    assign _991 = _774[39:39];
    assign _988 = _983 - _163;
    assign _989 = _985 ? _988 : _983;
    assign _990 = _989[62:0];
    assign _992 = { _990,
                    _991 };
    assign _993 = _992 < _163;
    assign _994 = ~ _993;
    assign _982 = _774[40:40];
    assign _979 = _974 - _163;
    assign _980 = _976 ? _979 : _974;
    assign _981 = _980[62:0];
    assign _983 = { _981,
                    _982 };
    assign _984 = _983 < _163;
    assign _985 = ~ _984;
    assign _973 = _774[41:41];
    assign _970 = _965 - _163;
    assign _971 = _967 ? _970 : _965;
    assign _972 = _971[62:0];
    assign _974 = { _972,
                    _973 };
    assign _975 = _974 < _163;
    assign _976 = ~ _975;
    assign _964 = _774[42:42];
    assign _961 = _956 - _163;
    assign _962 = _958 ? _961 : _956;
    assign _963 = _962[62:0];
    assign _965 = { _963,
                    _964 };
    assign _966 = _965 < _163;
    assign _967 = ~ _966;
    assign _955 = _774[43:43];
    assign _952 = _947 - _163;
    assign _953 = _949 ? _952 : _947;
    assign _954 = _953[62:0];
    assign _956 = { _954,
                    _955 };
    assign _957 = _956 < _163;
    assign _958 = ~ _957;
    assign _946 = _774[44:44];
    assign _943 = _938 - _163;
    assign _944 = _940 ? _943 : _938;
    assign _945 = _944[62:0];
    assign _947 = { _945,
                    _946 };
    assign _948 = _947 < _163;
    assign _949 = ~ _948;
    assign _937 = _774[45:45];
    assign _934 = _929 - _163;
    assign _935 = _931 ? _934 : _929;
    assign _936 = _935[62:0];
    assign _938 = { _936,
                    _937 };
    assign _939 = _938 < _163;
    assign _940 = ~ _939;
    assign _928 = _774[46:46];
    assign _925 = _920 - _163;
    assign _926 = _922 ? _925 : _920;
    assign _927 = _926[62:0];
    assign _929 = { _927,
                    _928 };
    assign _930 = _929 < _163;
    assign _931 = ~ _930;
    assign _919 = _774[47:47];
    assign _916 = _911 - _163;
    assign _917 = _913 ? _916 : _911;
    assign _918 = _917[62:0];
    assign _920 = { _918,
                    _919 };
    assign _921 = _920 < _163;
    assign _922 = ~ _921;
    assign _910 = _774[48:48];
    assign _907 = _902 - _163;
    assign _908 = _904 ? _907 : _902;
    assign _909 = _908[62:0];
    assign _911 = { _909,
                    _910 };
    assign _912 = _911 < _163;
    assign _913 = ~ _912;
    assign _901 = _774[49:49];
    assign _898 = _893 - _163;
    assign _899 = _895 ? _898 : _893;
    assign _900 = _899[62:0];
    assign _902 = { _900,
                    _901 };
    assign _903 = _902 < _163;
    assign _904 = ~ _903;
    assign _892 = _774[50:50];
    assign _889 = _884 - _163;
    assign _890 = _886 ? _889 : _884;
    assign _891 = _890[62:0];
    assign _893 = { _891,
                    _892 };
    assign _894 = _893 < _163;
    assign _895 = ~ _894;
    assign _883 = _774[51:51];
    assign _880 = _875 - _163;
    assign _881 = _877 ? _880 : _875;
    assign _882 = _881[62:0];
    assign _884 = { _882,
                    _883 };
    assign _885 = _884 < _163;
    assign _886 = ~ _885;
    assign _874 = _774[52:52];
    assign _871 = _866 - _163;
    assign _872 = _868 ? _871 : _866;
    assign _873 = _872[62:0];
    assign _875 = { _873,
                    _874 };
    assign _876 = _875 < _163;
    assign _877 = ~ _876;
    assign _865 = _774[53:53];
    assign _862 = _857 - _163;
    assign _863 = _859 ? _862 : _857;
    assign _864 = _863[62:0];
    assign _866 = { _864,
                    _865 };
    assign _867 = _866 < _163;
    assign _868 = ~ _867;
    assign _856 = _774[54:54];
    assign _853 = _848 - _163;
    assign _854 = _850 ? _853 : _848;
    assign _855 = _854[62:0];
    assign _857 = { _855,
                    _856 };
    assign _858 = _857 < _163;
    assign _859 = ~ _858;
    assign _847 = _774[55:55];
    assign _844 = _839 - _163;
    assign _845 = _841 ? _844 : _839;
    assign _846 = _845[62:0];
    assign _848 = { _846,
                    _847 };
    assign _849 = _848 < _163;
    assign _850 = ~ _849;
    assign _838 = _774[56:56];
    assign _835 = _830 - _163;
    assign _836 = _832 ? _835 : _830;
    assign _837 = _836[62:0];
    assign _839 = { _837,
                    _838 };
    assign _840 = _839 < _163;
    assign _841 = ~ _840;
    assign _829 = _774[57:57];
    assign _826 = _821 - _163;
    assign _827 = _823 ? _826 : _821;
    assign _828 = _827[62:0];
    assign _830 = { _828,
                    _829 };
    assign _831 = _830 < _163;
    assign _832 = ~ _831;
    assign _820 = _774[58:58];
    assign _817 = _812 - _163;
    assign _818 = _814 ? _817 : _812;
    assign _819 = _818[62:0];
    assign _821 = { _819,
                    _820 };
    assign _822 = _821 < _163;
    assign _823 = ~ _822;
    assign _811 = _774[59:59];
    assign _808 = _803 - _163;
    assign _809 = _805 ? _808 : _803;
    assign _810 = _809[62:0];
    assign _812 = { _810,
                    _811 };
    assign _813 = _812 < _163;
    assign _814 = ~ _813;
    assign _802 = _774[60:60];
    assign _799 = _794 - _163;
    assign _800 = _796 ? _799 : _794;
    assign _801 = _800[62:0];
    assign _803 = { _801,
                    _802 };
    assign _804 = _803 < _163;
    assign _805 = ~ _804;
    assign _793 = _774[61:61];
    assign _790 = _785 - _163;
    assign _791 = _787 ? _790 : _785;
    assign _792 = _791[62:0];
    assign _794 = { _792,
                    _793 };
    assign _795 = _794 < _163;
    assign _796 = ~ _795;
    assign _784 = _774[62:62];
    assign _781 = _776 - _163;
    assign _782 = _778 ? _781 : _776;
    assign _783 = _782[62:0];
    assign _785 = { _783,
                    _784 };
    assign _786 = _785 < _163;
    assign _787 = ~ _786;
    assign _774 = _104 - _742;
    assign _775 = _774[63:63];
    assign _776 = { _1352,
                    _775 };
    assign _777 = _776 < _163;
    assign _778 = ~ _777;
    assign _779 = { _1352,
                    _778 };
    assign _780 = _779[62:0];
    assign _788 = { _780,
                    _787 };
    assign _789 = _788[62:0];
    assign _797 = { _789,
                    _796 };
    assign _798 = _797[62:0];
    assign _806 = { _798,
                    _805 };
    assign _807 = _806[62:0];
    assign _815 = { _807,
                    _814 };
    assign _816 = _815[62:0];
    assign _824 = { _816,
                    _823 };
    assign _825 = _824[62:0];
    assign _833 = { _825,
                    _832 };
    assign _834 = _833[62:0];
    assign _842 = { _834,
                    _841 };
    assign _843 = _842[62:0];
    assign _851 = { _843,
                    _850 };
    assign _852 = _851[62:0];
    assign _860 = { _852,
                    _859 };
    assign _861 = _860[62:0];
    assign _869 = { _861,
                    _868 };
    assign _870 = _869[62:0];
    assign _878 = { _870,
                    _877 };
    assign _879 = _878[62:0];
    assign _887 = { _879,
                    _886 };
    assign _888 = _887[62:0];
    assign _896 = { _888,
                    _895 };
    assign _897 = _896[62:0];
    assign _905 = { _897,
                    _904 };
    assign _906 = _905[62:0];
    assign _914 = { _906,
                    _913 };
    assign _915 = _914[62:0];
    assign _923 = { _915,
                    _922 };
    assign _924 = _923[62:0];
    assign _932 = { _924,
                    _931 };
    assign _933 = _932[62:0];
    assign _941 = { _933,
                    _940 };
    assign _942 = _941[62:0];
    assign _950 = { _942,
                    _949 };
    assign _951 = _950[62:0];
    assign _959 = { _951,
                    _958 };
    assign _960 = _959[62:0];
    assign _968 = { _960,
                    _967 };
    assign _969 = _968[62:0];
    assign _977 = { _969,
                    _976 };
    assign _978 = _977[62:0];
    assign _986 = { _978,
                    _985 };
    assign _987 = _986[62:0];
    assign _995 = { _987,
                    _994 };
    assign _996 = _995[62:0];
    assign _1004 = { _996,
                     _1003 };
    assign _1005 = _1004[62:0];
    assign _1013 = { _1005,
                     _1012 };
    assign _1014 = _1013[62:0];
    assign _1022 = { _1014,
                     _1021 };
    assign _1023 = _1022[62:0];
    assign _1031 = { _1023,
                     _1030 };
    assign _1032 = _1031[62:0];
    assign _1040 = { _1032,
                     _1039 };
    assign _1041 = _1040[62:0];
    assign _1049 = { _1041,
                     _1048 };
    assign _1050 = _1049[62:0];
    assign _1058 = { _1050,
                     _1057 };
    assign _1059 = _1058[62:0];
    assign _1067 = { _1059,
                     _1066 };
    assign _1068 = _1067[62:0];
    assign _1076 = { _1068,
                     _1075 };
    assign _1077 = _1076[62:0];
    assign _1085 = { _1077,
                     _1084 };
    assign _1086 = _1085[62:0];
    assign _1094 = { _1086,
                     _1093 };
    assign _1095 = _1094[62:0];
    assign _1103 = { _1095,
                     _1102 };
    assign _1104 = _1103[62:0];
    assign _1112 = { _1104,
                     _1111 };
    assign _1113 = _1112[62:0];
    assign _1121 = { _1113,
                     _1120 };
    assign _1122 = _1121[62:0];
    assign _1130 = { _1122,
                     _1129 };
    assign _1131 = _1130[62:0];
    assign _1139 = { _1131,
                     _1138 };
    assign _1140 = _1139[62:0];
    assign _1148 = { _1140,
                     _1147 };
    assign _1149 = _1148[62:0];
    assign _1157 = { _1149,
                     _1156 };
    assign _1158 = _1157[62:0];
    assign _1166 = { _1158,
                     _1165 };
    assign _1167 = _1166[62:0];
    assign _1175 = { _1167,
                     _1174 };
    assign _1176 = _1175[62:0];
    assign _1184 = { _1176,
                     _1183 };
    assign _1185 = _1184[62:0];
    assign _1193 = { _1185,
                     _1192 };
    assign _1194 = _1193[62:0];
    assign _1202 = { _1194,
                     _1201 };
    assign _1203 = _1202[62:0];
    assign _1211 = { _1203,
                     _1210 };
    assign _1212 = _1211[62:0];
    assign _1220 = { _1212,
                     _1219 };
    assign _1221 = _1220[62:0];
    assign _1229 = { _1221,
                     _1228 };
    assign _1230 = _1229[62:0];
    assign _1238 = { _1230,
                     _1237 };
    assign _1239 = _1238[62:0];
    assign _1247 = { _1239,
                     _1246 };
    assign _1248 = _1247[62:0];
    assign _1256 = { _1248,
                     _1255 };
    assign _1257 = _1256[62:0];
    assign _1265 = { _1257,
                     _1264 };
    assign _1266 = _1265[62:0];
    assign _1274 = { _1266,
                     _1273 };
    assign _1275 = _1274[62:0];
    assign _1283 = { _1275,
                     _1282 };
    assign _1284 = _1283[62:0];
    assign _1292 = { _1284,
                     _1291 };
    assign _1293 = _1292[62:0];
    assign _1301 = { _1293,
                     _1300 };
    assign _1302 = _1301[62:0];
    assign _1310 = { _1302,
                     _1309 };
    assign _1311 = _1310[62:0];
    assign _1319 = { _1311,
                     _1318 };
    assign _1320 = _1319[62:0];
    assign _1328 = { _1320,
                     _1327 };
    assign _1329 = _1328[62:0];
    assign _1337 = { _1329,
                     _1336 };
    assign _1338 = _1337[62:0];
    assign _1346 = { _1338,
                     _1345 };
    assign _1348 = _1346 + _1353;
    assign _1349 = _742 * _1348;
    assign _1350 = _1349[63:0];
    assign _1932 = _1350 + _1931;
    assign _2010 = _75 ? vdd : vdd;
    assign _2011 = _73 ? vdd : _2010;
    assign _2012 = _71 ? vdd : _2011;
    assign _2013 = _69 ? vdd : _2012;
    assign _2014 = _67 ? vdd : _2013;
    assign _2016 = _65 ? _766 : _2014;
    assign _2018 = _63 ? _766 : _2016;
    assign _2020 = _61 ? _766 : _2018;
    assign _2022 = _59 ? _766 : _2020;
    assign _2024 = _57 ? _766 : _2022;
    assign _2026 = _55 ? _766 : _2024;
    assign _2028 = _53 ? _766 : _2026;
    assign _2030 = _51 ? _766 : _2028;
    assign _734 = _166[0:0];
    assign _731 = _726 - _163;
    assign _732 = _728 ? _731 : _726;
    assign _733 = _732[62:0];
    assign _735 = { _733,
                    _734 };
    assign _736 = _735 < _163;
    assign _737 = ~ _736;
    assign _725 = _166[1:1];
    assign _722 = _717 - _163;
    assign _723 = _719 ? _722 : _717;
    assign _724 = _723[62:0];
    assign _726 = { _724,
                    _725 };
    assign _727 = _726 < _163;
    assign _728 = ~ _727;
    assign _716 = _166[2:2];
    assign _713 = _708 - _163;
    assign _714 = _710 ? _713 : _708;
    assign _715 = _714[62:0];
    assign _717 = { _715,
                    _716 };
    assign _718 = _717 < _163;
    assign _719 = ~ _718;
    assign _707 = _166[3:3];
    assign _704 = _699 - _163;
    assign _705 = _701 ? _704 : _699;
    assign _706 = _705[62:0];
    assign _708 = { _706,
                    _707 };
    assign _709 = _708 < _163;
    assign _710 = ~ _709;
    assign _698 = _166[4:4];
    assign _695 = _690 - _163;
    assign _696 = _692 ? _695 : _690;
    assign _697 = _696[62:0];
    assign _699 = { _697,
                    _698 };
    assign _700 = _699 < _163;
    assign _701 = ~ _700;
    assign _689 = _166[5:5];
    assign _686 = _681 - _163;
    assign _687 = _683 ? _686 : _681;
    assign _688 = _687[62:0];
    assign _690 = { _688,
                    _689 };
    assign _691 = _690 < _163;
    assign _692 = ~ _691;
    assign _680 = _166[6:6];
    assign _677 = _672 - _163;
    assign _678 = _674 ? _677 : _672;
    assign _679 = _678[62:0];
    assign _681 = { _679,
                    _680 };
    assign _682 = _681 < _163;
    assign _683 = ~ _682;
    assign _671 = _166[7:7];
    assign _668 = _663 - _163;
    assign _669 = _665 ? _668 : _663;
    assign _670 = _669[62:0];
    assign _672 = { _670,
                    _671 };
    assign _673 = _672 < _163;
    assign _674 = ~ _673;
    assign _662 = _166[8:8];
    assign _659 = _654 - _163;
    assign _660 = _656 ? _659 : _654;
    assign _661 = _660[62:0];
    assign _663 = { _661,
                    _662 };
    assign _664 = _663 < _163;
    assign _665 = ~ _664;
    assign _653 = _166[9:9];
    assign _650 = _645 - _163;
    assign _651 = _647 ? _650 : _645;
    assign _652 = _651[62:0];
    assign _654 = { _652,
                    _653 };
    assign _655 = _654 < _163;
    assign _656 = ~ _655;
    assign _644 = _166[10:10];
    assign _641 = _636 - _163;
    assign _642 = _638 ? _641 : _636;
    assign _643 = _642[62:0];
    assign _645 = { _643,
                    _644 };
    assign _646 = _645 < _163;
    assign _647 = ~ _646;
    assign _635 = _166[11:11];
    assign _632 = _627 - _163;
    assign _633 = _629 ? _632 : _627;
    assign _634 = _633[62:0];
    assign _636 = { _634,
                    _635 };
    assign _637 = _636 < _163;
    assign _638 = ~ _637;
    assign _626 = _166[12:12];
    assign _623 = _618 - _163;
    assign _624 = _620 ? _623 : _618;
    assign _625 = _624[62:0];
    assign _627 = { _625,
                    _626 };
    assign _628 = _627 < _163;
    assign _629 = ~ _628;
    assign _617 = _166[13:13];
    assign _614 = _609 - _163;
    assign _615 = _611 ? _614 : _609;
    assign _616 = _615[62:0];
    assign _618 = { _616,
                    _617 };
    assign _619 = _618 < _163;
    assign _620 = ~ _619;
    assign _608 = _166[14:14];
    assign _605 = _600 - _163;
    assign _606 = _602 ? _605 : _600;
    assign _607 = _606[62:0];
    assign _609 = { _607,
                    _608 };
    assign _610 = _609 < _163;
    assign _611 = ~ _610;
    assign _599 = _166[15:15];
    assign _596 = _591 - _163;
    assign _597 = _593 ? _596 : _591;
    assign _598 = _597[62:0];
    assign _600 = { _598,
                    _599 };
    assign _601 = _600 < _163;
    assign _602 = ~ _601;
    assign _590 = _166[16:16];
    assign _587 = _582 - _163;
    assign _588 = _584 ? _587 : _582;
    assign _589 = _588[62:0];
    assign _591 = { _589,
                    _590 };
    assign _592 = _591 < _163;
    assign _593 = ~ _592;
    assign _581 = _166[17:17];
    assign _578 = _573 - _163;
    assign _579 = _575 ? _578 : _573;
    assign _580 = _579[62:0];
    assign _582 = { _580,
                    _581 };
    assign _583 = _582 < _163;
    assign _584 = ~ _583;
    assign _572 = _166[18:18];
    assign _569 = _564 - _163;
    assign _570 = _566 ? _569 : _564;
    assign _571 = _570[62:0];
    assign _573 = { _571,
                    _572 };
    assign _574 = _573 < _163;
    assign _575 = ~ _574;
    assign _563 = _166[19:19];
    assign _560 = _555 - _163;
    assign _561 = _557 ? _560 : _555;
    assign _562 = _561[62:0];
    assign _564 = { _562,
                    _563 };
    assign _565 = _564 < _163;
    assign _566 = ~ _565;
    assign _554 = _166[20:20];
    assign _551 = _546 - _163;
    assign _552 = _548 ? _551 : _546;
    assign _553 = _552[62:0];
    assign _555 = { _553,
                    _554 };
    assign _556 = _555 < _163;
    assign _557 = ~ _556;
    assign _545 = _166[21:21];
    assign _542 = _537 - _163;
    assign _543 = _539 ? _542 : _537;
    assign _544 = _543[62:0];
    assign _546 = { _544,
                    _545 };
    assign _547 = _546 < _163;
    assign _548 = ~ _547;
    assign _536 = _166[22:22];
    assign _533 = _528 - _163;
    assign _534 = _530 ? _533 : _528;
    assign _535 = _534[62:0];
    assign _537 = { _535,
                    _536 };
    assign _538 = _537 < _163;
    assign _539 = ~ _538;
    assign _527 = _166[23:23];
    assign _524 = _519 - _163;
    assign _525 = _521 ? _524 : _519;
    assign _526 = _525[62:0];
    assign _528 = { _526,
                    _527 };
    assign _529 = _528 < _163;
    assign _530 = ~ _529;
    assign _518 = _166[24:24];
    assign _515 = _510 - _163;
    assign _516 = _512 ? _515 : _510;
    assign _517 = _516[62:0];
    assign _519 = { _517,
                    _518 };
    assign _520 = _519 < _163;
    assign _521 = ~ _520;
    assign _509 = _166[25:25];
    assign _506 = _501 - _163;
    assign _507 = _503 ? _506 : _501;
    assign _508 = _507[62:0];
    assign _510 = { _508,
                    _509 };
    assign _511 = _510 < _163;
    assign _512 = ~ _511;
    assign _500 = _166[26:26];
    assign _497 = _492 - _163;
    assign _498 = _494 ? _497 : _492;
    assign _499 = _498[62:0];
    assign _501 = { _499,
                    _500 };
    assign _502 = _501 < _163;
    assign _503 = ~ _502;
    assign _491 = _166[27:27];
    assign _488 = _483 - _163;
    assign _489 = _485 ? _488 : _483;
    assign _490 = _489[62:0];
    assign _492 = { _490,
                    _491 };
    assign _493 = _492 < _163;
    assign _494 = ~ _493;
    assign _482 = _166[28:28];
    assign _479 = _474 - _163;
    assign _480 = _476 ? _479 : _474;
    assign _481 = _480[62:0];
    assign _483 = { _481,
                    _482 };
    assign _484 = _483 < _163;
    assign _485 = ~ _484;
    assign _473 = _166[29:29];
    assign _470 = _465 - _163;
    assign _471 = _467 ? _470 : _465;
    assign _472 = _471[62:0];
    assign _474 = { _472,
                    _473 };
    assign _475 = _474 < _163;
    assign _476 = ~ _475;
    assign _464 = _166[30:30];
    assign _461 = _456 - _163;
    assign _462 = _458 ? _461 : _456;
    assign _463 = _462[62:0];
    assign _465 = { _463,
                    _464 };
    assign _466 = _465 < _163;
    assign _467 = ~ _466;
    assign _455 = _166[31:31];
    assign _452 = _447 - _163;
    assign _453 = _449 ? _452 : _447;
    assign _454 = _453[62:0];
    assign _456 = { _454,
                    _455 };
    assign _457 = _456 < _163;
    assign _458 = ~ _457;
    assign _446 = _166[32:32];
    assign _443 = _438 - _163;
    assign _444 = _440 ? _443 : _438;
    assign _445 = _444[62:0];
    assign _447 = { _445,
                    _446 };
    assign _448 = _447 < _163;
    assign _449 = ~ _448;
    assign _437 = _166[33:33];
    assign _434 = _429 - _163;
    assign _435 = _431 ? _434 : _429;
    assign _436 = _435[62:0];
    assign _438 = { _436,
                    _437 };
    assign _439 = _438 < _163;
    assign _440 = ~ _439;
    assign _428 = _166[34:34];
    assign _425 = _420 - _163;
    assign _426 = _422 ? _425 : _420;
    assign _427 = _426[62:0];
    assign _429 = { _427,
                    _428 };
    assign _430 = _429 < _163;
    assign _431 = ~ _430;
    assign _419 = _166[35:35];
    assign _416 = _411 - _163;
    assign _417 = _413 ? _416 : _411;
    assign _418 = _417[62:0];
    assign _420 = { _418,
                    _419 };
    assign _421 = _420 < _163;
    assign _422 = ~ _421;
    assign _410 = _166[36:36];
    assign _407 = _402 - _163;
    assign _408 = _404 ? _407 : _402;
    assign _409 = _408[62:0];
    assign _411 = { _409,
                    _410 };
    assign _412 = _411 < _163;
    assign _413 = ~ _412;
    assign _401 = _166[37:37];
    assign _398 = _393 - _163;
    assign _399 = _395 ? _398 : _393;
    assign _400 = _399[62:0];
    assign _402 = { _400,
                    _401 };
    assign _403 = _402 < _163;
    assign _404 = ~ _403;
    assign _392 = _166[38:38];
    assign _389 = _384 - _163;
    assign _390 = _386 ? _389 : _384;
    assign _391 = _390[62:0];
    assign _393 = { _391,
                    _392 };
    assign _394 = _393 < _163;
    assign _395 = ~ _394;
    assign _383 = _166[39:39];
    assign _380 = _375 - _163;
    assign _381 = _377 ? _380 : _375;
    assign _382 = _381[62:0];
    assign _384 = { _382,
                    _383 };
    assign _385 = _384 < _163;
    assign _386 = ~ _385;
    assign _374 = _166[40:40];
    assign _371 = _366 - _163;
    assign _372 = _368 ? _371 : _366;
    assign _373 = _372[62:0];
    assign _375 = { _373,
                    _374 };
    assign _376 = _375 < _163;
    assign _377 = ~ _376;
    assign _365 = _166[41:41];
    assign _362 = _357 - _163;
    assign _363 = _359 ? _362 : _357;
    assign _364 = _363[62:0];
    assign _366 = { _364,
                    _365 };
    assign _367 = _366 < _163;
    assign _368 = ~ _367;
    assign _356 = _166[42:42];
    assign _353 = _348 - _163;
    assign _354 = _350 ? _353 : _348;
    assign _355 = _354[62:0];
    assign _357 = { _355,
                    _356 };
    assign _358 = _357 < _163;
    assign _359 = ~ _358;
    assign _347 = _166[43:43];
    assign _344 = _339 - _163;
    assign _345 = _341 ? _344 : _339;
    assign _346 = _345[62:0];
    assign _348 = { _346,
                    _347 };
    assign _349 = _348 < _163;
    assign _350 = ~ _349;
    assign _338 = _166[44:44];
    assign _335 = _330 - _163;
    assign _336 = _332 ? _335 : _330;
    assign _337 = _336[62:0];
    assign _339 = { _337,
                    _338 };
    assign _340 = _339 < _163;
    assign _341 = ~ _340;
    assign _329 = _166[45:45];
    assign _326 = _321 - _163;
    assign _327 = _323 ? _326 : _321;
    assign _328 = _327[62:0];
    assign _330 = { _328,
                    _329 };
    assign _331 = _330 < _163;
    assign _332 = ~ _331;
    assign _320 = _166[46:46];
    assign _317 = _312 - _163;
    assign _318 = _314 ? _317 : _312;
    assign _319 = _318[62:0];
    assign _321 = { _319,
                    _320 };
    assign _322 = _321 < _163;
    assign _323 = ~ _322;
    assign _311 = _166[47:47];
    assign _308 = _303 - _163;
    assign _309 = _305 ? _308 : _303;
    assign _310 = _309[62:0];
    assign _312 = { _310,
                    _311 };
    assign _313 = _312 < _163;
    assign _314 = ~ _313;
    assign _302 = _166[48:48];
    assign _299 = _294 - _163;
    assign _300 = _296 ? _299 : _294;
    assign _301 = _300[62:0];
    assign _303 = { _301,
                    _302 };
    assign _304 = _303 < _163;
    assign _305 = ~ _304;
    assign _293 = _166[49:49];
    assign _290 = _285 - _163;
    assign _291 = _287 ? _290 : _285;
    assign _292 = _291[62:0];
    assign _294 = { _292,
                    _293 };
    assign _295 = _294 < _163;
    assign _296 = ~ _295;
    assign _284 = _166[50:50];
    assign _281 = _276 - _163;
    assign _282 = _278 ? _281 : _276;
    assign _283 = _282[62:0];
    assign _285 = { _283,
                    _284 };
    assign _286 = _285 < _163;
    assign _287 = ~ _286;
    assign _275 = _166[51:51];
    assign _272 = _267 - _163;
    assign _273 = _269 ? _272 : _267;
    assign _274 = _273[62:0];
    assign _276 = { _274,
                    _275 };
    assign _277 = _276 < _163;
    assign _278 = ~ _277;
    assign _266 = _166[52:52];
    assign _263 = _258 - _163;
    assign _264 = _260 ? _263 : _258;
    assign _265 = _264[62:0];
    assign _267 = { _265,
                    _266 };
    assign _268 = _267 < _163;
    assign _269 = ~ _268;
    assign _257 = _166[53:53];
    assign _254 = _249 - _163;
    assign _255 = _251 ? _254 : _249;
    assign _256 = _255[62:0];
    assign _258 = { _256,
                    _257 };
    assign _259 = _258 < _163;
    assign _260 = ~ _259;
    assign _248 = _166[54:54];
    assign _245 = _240 - _163;
    assign _246 = _242 ? _245 : _240;
    assign _247 = _246[62:0];
    assign _249 = { _247,
                    _248 };
    assign _250 = _249 < _163;
    assign _251 = ~ _250;
    assign _239 = _166[55:55];
    assign _236 = _231 - _163;
    assign _237 = _233 ? _236 : _231;
    assign _238 = _237[62:0];
    assign _240 = { _238,
                    _239 };
    assign _241 = _240 < _163;
    assign _242 = ~ _241;
    assign _230 = _166[56:56];
    assign _227 = _222 - _163;
    assign _228 = _224 ? _227 : _222;
    assign _229 = _228[62:0];
    assign _231 = { _229,
                    _230 };
    assign _232 = _231 < _163;
    assign _233 = ~ _232;
    assign _221 = _166[57:57];
    assign _218 = _213 - _163;
    assign _219 = _215 ? _218 : _213;
    assign _220 = _219[62:0];
    assign _222 = { _220,
                    _221 };
    assign _223 = _222 < _163;
    assign _224 = ~ _223;
    assign _212 = _166[58:58];
    assign _209 = _204 - _163;
    assign _210 = _206 ? _209 : _204;
    assign _211 = _210[62:0];
    assign _213 = { _211,
                    _212 };
    assign _214 = _213 < _163;
    assign _215 = ~ _214;
    assign _203 = _166[59:59];
    assign _200 = _195 - _163;
    assign _201 = _197 ? _200 : _195;
    assign _202 = _201[62:0];
    assign _204 = { _202,
                    _203 };
    assign _205 = _204 < _163;
    assign _206 = ~ _205;
    assign _194 = _166[60:60];
    assign _191 = _186 - _163;
    assign _192 = _188 ? _191 : _186;
    assign _193 = _192[62:0];
    assign _195 = { _193,
                    _194 };
    assign _196 = _195 < _163;
    assign _197 = ~ _196;
    assign _185 = _166[61:61];
    assign _182 = _177 - _163;
    assign _183 = _179 ? _182 : _177;
    assign _184 = _183[62:0];
    assign _186 = { _184,
                    _185 };
    assign _187 = _186 < _163;
    assign _188 = ~ _187;
    assign _176 = _166[62:62];
    assign _173 = _168 - _163;
    assign _174 = _170 ? _173 : _168;
    assign _175 = _174[62:0];
    assign _177 = { _175,
                    _176 };
    assign _178 = _177 < _163;
    assign _179 = ~ _178;
    assign _162 = 64'b0000000000000000000000000000000001000010001110100011010111000111;
    assign _160 = 64'b0000000000000000000000000000000000000000000000011011001000000111;
    assign _158 = 64'b0000000000000000000000000000000000000110000001010100101010110101;
    assign _156 = 64'b0000000000000000000000000000000000000000000011110100011000101001;
    assign _154 = 64'b0000000000000000000000000000000000000000000100001111010001000111;
    assign _152 = 64'b0000000000000000000000000000000000000000000000000010011101110101;
    assign _150 = 64'b0000000000000000000000000000000000000000000000000010101101100111;
    assign _148 = 64'b0000000000000000000000000000000000000000000000000000000001101111;
    assign _146 = 64'b0000000000000000000000000000000000000000000000011000011010100001;
    assign _144 = 64'b0000000000000000000000000000000000000000000000000010011100010001;
    assign _142 = 64'b0000000000000000000000000000000000000000000000000000001111101001;
    assign _140 = 64'b0000000000000000000000000000000000000000000000000000000001100101;
    assign _138 = 64'b0000000000000000000000000000000000000000000000000000000000001011;
    assign _139 = _75 ? _138 : _138;
    assign _141 = _73 ? _140 : _139;
    assign _143 = _71 ? _142 : _141;
    assign _145 = _69 ? _144 : _143;
    assign _147 = _67 ? _146 : _145;
    assign _149 = _65 ? _148 : _147;
    assign _151 = _63 ? _150 : _149;
    assign _153 = _61 ? _152 : _151;
    assign _155 = _59 ? _154 : _153;
    assign _157 = _57 ? _156 : _155;
    assign _159 = _55 ? _158 : _157;
    assign _161 = _53 ? _160 : _159;
    assign _163 = _51 ? _162 : _161;
    assign _165 = _163 - _1353;
    assign _8 = from_;
    assign _1977 = _1976 ? _8 : _136;
    assign _1979 = _26 ? _45 : _1977;
    assign _9 = _1979;
    always @(posedge _19) begin
        if (_17)
            _136 <= _45;
        else
            _136 <= _9;
    end
    assign _166 = _136 + _165;
    assign _167 = _166[63:63];
    assign _168 = { _1352,
                    _167 };
    assign _169 = _168 < _163;
    assign _170 = ~ _169;
    assign _171 = { _1352,
                    _170 };
    assign _172 = _171[62:0];
    assign _180 = { _172,
                    _179 };
    assign _181 = _180[62:0];
    assign _189 = { _181,
                    _188 };
    assign _190 = _189[62:0];
    assign _198 = { _190,
                    _197 };
    assign _199 = _198[62:0];
    assign _207 = { _199,
                    _206 };
    assign _208 = _207[62:0];
    assign _216 = { _208,
                    _215 };
    assign _217 = _216[62:0];
    assign _225 = { _217,
                    _224 };
    assign _226 = _225[62:0];
    assign _234 = { _226,
                    _233 };
    assign _235 = _234[62:0];
    assign _243 = { _235,
                    _242 };
    assign _244 = _243[62:0];
    assign _252 = { _244,
                    _251 };
    assign _253 = _252[62:0];
    assign _261 = { _253,
                    _260 };
    assign _262 = _261[62:0];
    assign _270 = { _262,
                    _269 };
    assign _271 = _270[62:0];
    assign _279 = { _271,
                    _278 };
    assign _280 = _279[62:0];
    assign _288 = { _280,
                    _287 };
    assign _289 = _288[62:0];
    assign _297 = { _289,
                    _296 };
    assign _298 = _297[62:0];
    assign _306 = { _298,
                    _305 };
    assign _307 = _306[62:0];
    assign _315 = { _307,
                    _314 };
    assign _316 = _315[62:0];
    assign _324 = { _316,
                    _323 };
    assign _325 = _324[62:0];
    assign _333 = { _325,
                    _332 };
    assign _334 = _333[62:0];
    assign _342 = { _334,
                    _341 };
    assign _343 = _342[62:0];
    assign _351 = { _343,
                    _350 };
    assign _352 = _351[62:0];
    assign _360 = { _352,
                    _359 };
    assign _361 = _360[62:0];
    assign _369 = { _361,
                    _368 };
    assign _370 = _369[62:0];
    assign _378 = { _370,
                    _377 };
    assign _379 = _378[62:0];
    assign _387 = { _379,
                    _386 };
    assign _388 = _387[62:0];
    assign _396 = { _388,
                    _395 };
    assign _397 = _396[62:0];
    assign _405 = { _397,
                    _404 };
    assign _406 = _405[62:0];
    assign _414 = { _406,
                    _413 };
    assign _415 = _414[62:0];
    assign _423 = { _415,
                    _422 };
    assign _424 = _423[62:0];
    assign _432 = { _424,
                    _431 };
    assign _433 = _432[62:0];
    assign _441 = { _433,
                    _440 };
    assign _442 = _441[62:0];
    assign _450 = { _442,
                    _449 };
    assign _451 = _450[62:0];
    assign _459 = { _451,
                    _458 };
    assign _460 = _459[62:0];
    assign _468 = { _460,
                    _467 };
    assign _469 = _468[62:0];
    assign _477 = { _469,
                    _476 };
    assign _478 = _477[62:0];
    assign _486 = { _478,
                    _485 };
    assign _487 = _486[62:0];
    assign _495 = { _487,
                    _494 };
    assign _496 = _495[62:0];
    assign _504 = { _496,
                    _503 };
    assign _505 = _504[62:0];
    assign _513 = { _505,
                    _512 };
    assign _514 = _513[62:0];
    assign _522 = { _514,
                    _521 };
    assign _523 = _522[62:0];
    assign _531 = { _523,
                    _530 };
    assign _532 = _531[62:0];
    assign _540 = { _532,
                    _539 };
    assign _541 = _540[62:0];
    assign _549 = { _541,
                    _548 };
    assign _550 = _549[62:0];
    assign _558 = { _550,
                    _557 };
    assign _559 = _558[62:0];
    assign _567 = { _559,
                    _566 };
    assign _568 = _567[62:0];
    assign _576 = { _568,
                    _575 };
    assign _577 = _576[62:0];
    assign _585 = { _577,
                    _584 };
    assign _586 = _585[62:0];
    assign _594 = { _586,
                    _593 };
    assign _595 = _594[62:0];
    assign _603 = { _595,
                    _602 };
    assign _604 = _603[62:0];
    assign _612 = { _604,
                    _611 };
    assign _613 = _612[62:0];
    assign _621 = { _613,
                    _620 };
    assign _622 = _621[62:0];
    assign _630 = { _622,
                    _629 };
    assign _631 = _630[62:0];
    assign _639 = { _631,
                    _638 };
    assign _640 = _639[62:0];
    assign _648 = { _640,
                    _647 };
    assign _649 = _648[62:0];
    assign _657 = { _649,
                    _656 };
    assign _658 = _657[62:0];
    assign _666 = { _658,
                    _665 };
    assign _667 = _666[62:0];
    assign _675 = { _667,
                    _674 };
    assign _676 = _675[62:0];
    assign _684 = { _676,
                    _683 };
    assign _685 = _684[62:0];
    assign _693 = { _685,
                    _692 };
    assign _694 = _693[62:0];
    assign _702 = { _694,
                    _701 };
    assign _703 = _702[62:0];
    assign _711 = { _703,
                    _710 };
    assign _712 = _711[62:0];
    assign _720 = { _712,
                    _719 };
    assign _721 = _720[62:0];
    assign _729 = { _721,
                    _728 };
    assign _730 = _729[62:0];
    assign _738 = { _730,
                    _737 };
    assign _739 = _738 * _163;
    assign _740 = _739[63:0];
    assign _126 = 64'b0000000000000000000000000000000000111100001101001110101100010010;
    assign _124 = 64'b0000000000000000000000000000000000000101111101110110100000000100;
    assign _120 = 64'b0000000000000000000000000000000000000000000000011000101010010010;
    assign _114 = 64'b0000000000000000000000000000000000111011100110101111000100010000;
    assign _112 = 64'b0000000000000000000000000000000000000000100110001001101001101000;
    assign _110 = 64'b0000000000000000000000000000000000000000000000011000011100000100;
    assign _108 = 64'b0000000000000000000000000000000000000000000000000000001111110010;
    assign _107 = _75 ? _138 : _138;
    assign _109 = _73 ? _108 : _107;
    assign _111 = _71 ? _110 : _109;
    assign _113 = _69 ? _112 : _111;
    assign _115 = _67 ? _114 : _113;
    assign _117 = _65 ? _148 : _115;
    assign _119 = _63 ? _150 : _117;
    assign _121 = _61 ? _120 : _119;
    assign _123 = _59 ? _154 : _121;
    assign _125 = _57 ? _124 : _123;
    assign _127 = _55 ? _126 : _125;
    assign _129 = _53 ? _160 : _127;
    assign _131 = _51 ? _162 : _129;
    assign _741 = _131 < _740;
    assign _742 = _741 ? _740 : _131;
    assign _101 = 64'b0000000000000000000000000000001001010100000010111110001111111111;
    assign _99 = 64'b0000000000000000000000000000000000000000000011110100001000111111;
    assign _95 = 64'b0000000000000000000000000000000000111011100110101100100111111111;
    assign _93 = 64'b0000000000000000000000000000000000000000100110001001011001111111;
    assign _89 = 64'b0000000000000000000000000000000000000000000000011000011010011111;
    assign _87 = 64'b0000000000000000000000000000000000000000000000000000001111100111;
    assign _83 = 64'b0000000000000000000000000000000000000101111101011110000011111111;
    assign _79 = 64'b0000000000000000000000000000000000000000000000000010011100001111;
    assign _77 = 64'b0000000000000000000000000000000000000000000000000000000001100011;
    assign _74 = 4'b0000;
    assign _75 = _32 == _74;
    assign _78 = _75 ? _77 : _77;
    assign _72 = 4'b0001;
    assign _73 = _32 == _72;
    assign _80 = _73 ? _79 : _78;
    assign _70 = 4'b0010;
    assign _71 = _32 == _70;
    assign _82 = _71 ? _99 : _80;
    assign _68 = 4'b0011;
    assign _69 = _32 == _68;
    assign _84 = _69 ? _83 : _82;
    assign _66 = 4'b0100;
    assign _67 = _32 == _66;
    assign _86 = _67 ? _101 : _84;
    assign _64 = 4'b0101;
    assign _65 = _32 == _64;
    assign _88 = _65 ? _87 : _86;
    assign _62 = 4'b0110;
    assign _63 = _32 == _62;
    assign _90 = _63 ? _89 : _88;
    assign _60 = 4'b0111;
    assign _61 = _32 == _60;
    assign _92 = _61 ? _99 : _90;
    assign _58 = 4'b1000;
    assign _59 = _32 == _58;
    assign _94 = _59 ? _93 : _92;
    assign _56 = 4'b1001;
    assign _57 = _32 == _56;
    assign _96 = _57 ? _95 : _94;
    assign _54 = 4'b1010;
    assign _55 = _32 == _54;
    assign _98 = _55 ? _101 : _96;
    assign _52 = 4'b1011;
    assign _53 = _32 == _52;
    assign _100 = _53 ? _99 : _98;
    assign _50 = 4'b1100;
    assign _51 = _32 == _50;
    assign _102 = _51 ? _101 : _100;
    assign _11 = to_;
    assign _1980 = _1976 ? _11 : _49;
    assign _1982 = _26 ? _45 : _1980;
    assign _12 = _1982;
    always @(posedge _19) begin
        if (_17)
            _49 <= _45;
        else
            _49 <= _12;
    end
    assign _103 = _49 < _102;
    assign _104 = _103 ? _49 : _102;
    assign _743 = _104 < _742;
    assign _744 = ~ _743;
    assign _2031 = _744 & _2030;
    assign _2033 = _2031 ? _1932 : _45;
    assign _2034 = _1973 + _2033;
    assign _2008 = ~ _35;
    assign _2004 = _1997 ? _766 : _38;
    assign _14 = last;
    assign _1986 = _1976 ? _14 : _1985;
    assign _1988 = _26 ? _766 : _1986;
    assign _15 = _1988;
    always @(posedge _19) begin
        if (_17)
            _1985 <= _766;
        else
            _1985 <= _15;
    end
    assign vdd = 1'b1;
    assign _17 = clear;
    assign _19 = clock;
    assign _1990 = _32 + _72;
    assign _1991 = _38 ? _1990 : _32;
    assign _1993 = _1976 ? _74 : _1991;
    assign _1995 = _26 ? _74 : _1993;
    assign _20 = _1995;
    always @(posedge _19) begin
        if (_17)
            _32 <= _74;
        else
            _32 <= _20;
    end
    assign _1997 = _32 == _50;
    assign _1998 = _38 & _1997;
    assign _1999 = _1998 & _1985;
    assign _2000 = _1999 ? vdd : _35;
    assign _2002 = _26 ? _766 : _2000;
    assign _21 = _2002;
    always @(posedge _19) begin
        if (_17)
            _35 <= _766;
        else
            _35 <= _21;
    end
    assign _40 = ~ _35;
    assign _39 = ~ _38;
    assign _41 = _39 & _40;
    assign _23 = pair_valid;
    assign _1976 = _23 & _41;
    assign _2005 = _1976 ? vdd : _2004;
    assign _2007 = _26 ? _766 : _2005;
    assign _24 = _2007;
    always @(posedge _19) begin
        if (_17)
            _38 <= _766;
        else
            _38 <= _24;
    end
    assign _2009 = _38 & _2008;
    assign _2035 = _2009 ? _2034 : _1973;
    assign _26 = load;
    assign _2037 = _26 ? _45 : _2035;
    assign _27 = _2037;
    always @(posedge _19) begin
        if (_17)
            _1973 <= _45;
        else
            _1973 <= _27;
    end
    assign sum_p1 = _1973;
    assign sum_p2 = _1975;
    assign ready = _41;
    assign done_ = _35;
    assign family_index = _32;

endmodule
