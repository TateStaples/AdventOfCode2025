module day2_opt_c_family_unroll (
    from_,
    to_,
    sum_p1,
    sum_p2
);

    input [63:0] from_;
    input [63:0] to_;
    output [63:0] sum_p1;
    output [63:0] sum_p2;

    wire _22758;
    wire [63:0] _22755;
    wire [63:0] _22756;
    wire [62:0] _22757;
    wire [63:0] _22759;
    wire _22760;
    wire _22761;
    wire _22749;
    wire [63:0] _22746;
    wire [63:0] _22747;
    wire [62:0] _22748;
    wire [63:0] _22750;
    wire _22751;
    wire _22752;
    wire _22740;
    wire [63:0] _22737;
    wire [63:0] _22738;
    wire [62:0] _22739;
    wire [63:0] _22741;
    wire _22742;
    wire _22743;
    wire _22731;
    wire [63:0] _22728;
    wire [63:0] _22729;
    wire [62:0] _22730;
    wire [63:0] _22732;
    wire _22733;
    wire _22734;
    wire _22722;
    wire [63:0] _22719;
    wire [63:0] _22720;
    wire [62:0] _22721;
    wire [63:0] _22723;
    wire _22724;
    wire _22725;
    wire _22713;
    wire [63:0] _22710;
    wire [63:0] _22711;
    wire [62:0] _22712;
    wire [63:0] _22714;
    wire _22715;
    wire _22716;
    wire _22704;
    wire [63:0] _22701;
    wire [63:0] _22702;
    wire [62:0] _22703;
    wire [63:0] _22705;
    wire _22706;
    wire _22707;
    wire _22695;
    wire [63:0] _22692;
    wire [63:0] _22693;
    wire [62:0] _22694;
    wire [63:0] _22696;
    wire _22697;
    wire _22698;
    wire _22686;
    wire [63:0] _22683;
    wire [63:0] _22684;
    wire [62:0] _22685;
    wire [63:0] _22687;
    wire _22688;
    wire _22689;
    wire _22677;
    wire [63:0] _22674;
    wire [63:0] _22675;
    wire [62:0] _22676;
    wire [63:0] _22678;
    wire _22679;
    wire _22680;
    wire _22668;
    wire [63:0] _22665;
    wire [63:0] _22666;
    wire [62:0] _22667;
    wire [63:0] _22669;
    wire _22670;
    wire _22671;
    wire _22659;
    wire [63:0] _22656;
    wire [63:0] _22657;
    wire [62:0] _22658;
    wire [63:0] _22660;
    wire _22661;
    wire _22662;
    wire _22650;
    wire [63:0] _22647;
    wire [63:0] _22648;
    wire [62:0] _22649;
    wire [63:0] _22651;
    wire _22652;
    wire _22653;
    wire _22641;
    wire [63:0] _22638;
    wire [63:0] _22639;
    wire [62:0] _22640;
    wire [63:0] _22642;
    wire _22643;
    wire _22644;
    wire _22632;
    wire [63:0] _22629;
    wire [63:0] _22630;
    wire [62:0] _22631;
    wire [63:0] _22633;
    wire _22634;
    wire _22635;
    wire _22623;
    wire [63:0] _22620;
    wire [63:0] _22621;
    wire [62:0] _22622;
    wire [63:0] _22624;
    wire _22625;
    wire _22626;
    wire _22614;
    wire [63:0] _22611;
    wire [63:0] _22612;
    wire [62:0] _22613;
    wire [63:0] _22615;
    wire _22616;
    wire _22617;
    wire _22605;
    wire [63:0] _22602;
    wire [63:0] _22603;
    wire [62:0] _22604;
    wire [63:0] _22606;
    wire _22607;
    wire _22608;
    wire _22596;
    wire [63:0] _22593;
    wire [63:0] _22594;
    wire [62:0] _22595;
    wire [63:0] _22597;
    wire _22598;
    wire _22599;
    wire _22587;
    wire [63:0] _22584;
    wire [63:0] _22585;
    wire [62:0] _22586;
    wire [63:0] _22588;
    wire _22589;
    wire _22590;
    wire _22578;
    wire [63:0] _22575;
    wire [63:0] _22576;
    wire [62:0] _22577;
    wire [63:0] _22579;
    wire _22580;
    wire _22581;
    wire _22569;
    wire [63:0] _22566;
    wire [63:0] _22567;
    wire [62:0] _22568;
    wire [63:0] _22570;
    wire _22571;
    wire _22572;
    wire _22560;
    wire [63:0] _22557;
    wire [63:0] _22558;
    wire [62:0] _22559;
    wire [63:0] _22561;
    wire _22562;
    wire _22563;
    wire _22551;
    wire [63:0] _22548;
    wire [63:0] _22549;
    wire [62:0] _22550;
    wire [63:0] _22552;
    wire _22553;
    wire _22554;
    wire _22542;
    wire [63:0] _22539;
    wire [63:0] _22540;
    wire [62:0] _22541;
    wire [63:0] _22543;
    wire _22544;
    wire _22545;
    wire _22533;
    wire [63:0] _22530;
    wire [63:0] _22531;
    wire [62:0] _22532;
    wire [63:0] _22534;
    wire _22535;
    wire _22536;
    wire _22524;
    wire [63:0] _22521;
    wire [63:0] _22522;
    wire [62:0] _22523;
    wire [63:0] _22525;
    wire _22526;
    wire _22527;
    wire _22515;
    wire [63:0] _22512;
    wire [63:0] _22513;
    wire [62:0] _22514;
    wire [63:0] _22516;
    wire _22517;
    wire _22518;
    wire _22506;
    wire [63:0] _22503;
    wire [63:0] _22504;
    wire [62:0] _22505;
    wire [63:0] _22507;
    wire _22508;
    wire _22509;
    wire _22497;
    wire [63:0] _22494;
    wire [63:0] _22495;
    wire [62:0] _22496;
    wire [63:0] _22498;
    wire _22499;
    wire _22500;
    wire _22488;
    wire [63:0] _22485;
    wire [63:0] _22486;
    wire [62:0] _22487;
    wire [63:0] _22489;
    wire _22490;
    wire _22491;
    wire _22479;
    wire [63:0] _22476;
    wire [63:0] _22477;
    wire [62:0] _22478;
    wire [63:0] _22480;
    wire _22481;
    wire _22482;
    wire _22470;
    wire [63:0] _22467;
    wire [63:0] _22468;
    wire [62:0] _22469;
    wire [63:0] _22471;
    wire _22472;
    wire _22473;
    wire _22461;
    wire [63:0] _22458;
    wire [63:0] _22459;
    wire [62:0] _22460;
    wire [63:0] _22462;
    wire _22463;
    wire _22464;
    wire _22452;
    wire [63:0] _22449;
    wire [63:0] _22450;
    wire [62:0] _22451;
    wire [63:0] _22453;
    wire _22454;
    wire _22455;
    wire _22443;
    wire [63:0] _22440;
    wire [63:0] _22441;
    wire [62:0] _22442;
    wire [63:0] _22444;
    wire _22445;
    wire _22446;
    wire _22434;
    wire [63:0] _22431;
    wire [63:0] _22432;
    wire [62:0] _22433;
    wire [63:0] _22435;
    wire _22436;
    wire _22437;
    wire _22425;
    wire [63:0] _22422;
    wire [63:0] _22423;
    wire [62:0] _22424;
    wire [63:0] _22426;
    wire _22427;
    wire _22428;
    wire _22416;
    wire [63:0] _22413;
    wire [63:0] _22414;
    wire [62:0] _22415;
    wire [63:0] _22417;
    wire _22418;
    wire _22419;
    wire _22407;
    wire [63:0] _22404;
    wire [63:0] _22405;
    wire [62:0] _22406;
    wire [63:0] _22408;
    wire _22409;
    wire _22410;
    wire _22398;
    wire [63:0] _22395;
    wire [63:0] _22396;
    wire [62:0] _22397;
    wire [63:0] _22399;
    wire _22400;
    wire _22401;
    wire _22389;
    wire [63:0] _22386;
    wire [63:0] _22387;
    wire [62:0] _22388;
    wire [63:0] _22390;
    wire _22391;
    wire _22392;
    wire _22380;
    wire [63:0] _22377;
    wire [63:0] _22378;
    wire [62:0] _22379;
    wire [63:0] _22381;
    wire _22382;
    wire _22383;
    wire _22371;
    wire [63:0] _22368;
    wire [63:0] _22369;
    wire [62:0] _22370;
    wire [63:0] _22372;
    wire _22373;
    wire _22374;
    wire _22362;
    wire [63:0] _22359;
    wire [63:0] _22360;
    wire [62:0] _22361;
    wire [63:0] _22363;
    wire _22364;
    wire _22365;
    wire _22353;
    wire [63:0] _22350;
    wire [63:0] _22351;
    wire [62:0] _22352;
    wire [63:0] _22354;
    wire _22355;
    wire _22356;
    wire _22344;
    wire [63:0] _22341;
    wire [63:0] _22342;
    wire [62:0] _22343;
    wire [63:0] _22345;
    wire _22346;
    wire _22347;
    wire _22335;
    wire [63:0] _22332;
    wire [63:0] _22333;
    wire [62:0] _22334;
    wire [63:0] _22336;
    wire _22337;
    wire _22338;
    wire _22326;
    wire [63:0] _22323;
    wire [63:0] _22324;
    wire [62:0] _22325;
    wire [63:0] _22327;
    wire _22328;
    wire _22329;
    wire _22317;
    wire [63:0] _22314;
    wire [63:0] _22315;
    wire [62:0] _22316;
    wire [63:0] _22318;
    wire _22319;
    wire _22320;
    wire _22308;
    wire [63:0] _22305;
    wire [63:0] _22306;
    wire [62:0] _22307;
    wire [63:0] _22309;
    wire _22310;
    wire _22311;
    wire _22299;
    wire [63:0] _22296;
    wire [63:0] _22297;
    wire [62:0] _22298;
    wire [63:0] _22300;
    wire _22301;
    wire _22302;
    wire _22290;
    wire [63:0] _22287;
    wire [63:0] _22288;
    wire [62:0] _22289;
    wire [63:0] _22291;
    wire _22292;
    wire _22293;
    wire _22281;
    wire [63:0] _22278;
    wire [63:0] _22279;
    wire [62:0] _22280;
    wire [63:0] _22282;
    wire _22283;
    wire _22284;
    wire _22272;
    wire [63:0] _22269;
    wire [63:0] _22270;
    wire [62:0] _22271;
    wire [63:0] _22273;
    wire _22274;
    wire _22275;
    wire _22263;
    wire [63:0] _22260;
    wire [63:0] _22261;
    wire [62:0] _22262;
    wire [63:0] _22264;
    wire _22265;
    wire _22266;
    wire _22254;
    wire [63:0] _22251;
    wire [63:0] _22252;
    wire [62:0] _22253;
    wire [63:0] _22255;
    wire _22256;
    wire _22257;
    wire _22245;
    wire [63:0] _22242;
    wire [63:0] _22243;
    wire [62:0] _22244;
    wire [63:0] _22246;
    wire _22247;
    wire _22248;
    wire _22236;
    wire [63:0] _22233;
    wire [63:0] _22234;
    wire [62:0] _22235;
    wire [63:0] _22237;
    wire _22238;
    wire _22239;
    wire _22227;
    wire [63:0] _22224;
    wire [63:0] _22225;
    wire [62:0] _22226;
    wire [63:0] _22228;
    wire _22229;
    wire _22230;
    wire _22218;
    wire [63:0] _22215;
    wire [63:0] _22216;
    wire [62:0] _22217;
    wire [63:0] _22219;
    wire _22220;
    wire _22221;
    wire _22209;
    wire [63:0] _22206;
    wire [63:0] _22207;
    wire [62:0] _22208;
    wire [63:0] _22210;
    wire _22211;
    wire _22212;
    wire _22200;
    wire [63:0] _22197;
    wire [63:0] _22198;
    wire [62:0] _22199;
    wire [63:0] _22201;
    wire _22202;
    wire _22203;
    wire [63:0] _22192;
    wire [63:0] _22186;
    wire [63:0] _22187;
    wire [127:0] _22188;
    wire [63:0] _22189;
    wire _22190;
    wire [62:0] _22185;
    wire [63:0] _22191;
    wire _22193;
    wire _22194;
    wire [63:0] _22195;
    wire [62:0] _22196;
    wire [63:0] _22204;
    wire [62:0] _22205;
    wire [63:0] _22213;
    wire [62:0] _22214;
    wire [63:0] _22222;
    wire [62:0] _22223;
    wire [63:0] _22231;
    wire [62:0] _22232;
    wire [63:0] _22240;
    wire [62:0] _22241;
    wire [63:0] _22249;
    wire [62:0] _22250;
    wire [63:0] _22258;
    wire [62:0] _22259;
    wire [63:0] _22267;
    wire [62:0] _22268;
    wire [63:0] _22276;
    wire [62:0] _22277;
    wire [63:0] _22285;
    wire [62:0] _22286;
    wire [63:0] _22294;
    wire [62:0] _22295;
    wire [63:0] _22303;
    wire [62:0] _22304;
    wire [63:0] _22312;
    wire [62:0] _22313;
    wire [63:0] _22321;
    wire [62:0] _22322;
    wire [63:0] _22330;
    wire [62:0] _22331;
    wire [63:0] _22339;
    wire [62:0] _22340;
    wire [63:0] _22348;
    wire [62:0] _22349;
    wire [63:0] _22357;
    wire [62:0] _22358;
    wire [63:0] _22366;
    wire [62:0] _22367;
    wire [63:0] _22375;
    wire [62:0] _22376;
    wire [63:0] _22384;
    wire [62:0] _22385;
    wire [63:0] _22393;
    wire [62:0] _22394;
    wire [63:0] _22402;
    wire [62:0] _22403;
    wire [63:0] _22411;
    wire [62:0] _22412;
    wire [63:0] _22420;
    wire [62:0] _22421;
    wire [63:0] _22429;
    wire [62:0] _22430;
    wire [63:0] _22438;
    wire [62:0] _22439;
    wire [63:0] _22447;
    wire [62:0] _22448;
    wire [63:0] _22456;
    wire [62:0] _22457;
    wire [63:0] _22465;
    wire [62:0] _22466;
    wire [63:0] _22474;
    wire [62:0] _22475;
    wire [63:0] _22483;
    wire [62:0] _22484;
    wire [63:0] _22492;
    wire [62:0] _22493;
    wire [63:0] _22501;
    wire [62:0] _22502;
    wire [63:0] _22510;
    wire [62:0] _22511;
    wire [63:0] _22519;
    wire [62:0] _22520;
    wire [63:0] _22528;
    wire [62:0] _22529;
    wire [63:0] _22537;
    wire [62:0] _22538;
    wire [63:0] _22546;
    wire [62:0] _22547;
    wire [63:0] _22555;
    wire [62:0] _22556;
    wire [63:0] _22564;
    wire [62:0] _22565;
    wire [63:0] _22573;
    wire [62:0] _22574;
    wire [63:0] _22582;
    wire [62:0] _22583;
    wire [63:0] _22591;
    wire [62:0] _22592;
    wire [63:0] _22600;
    wire [62:0] _22601;
    wire [63:0] _22609;
    wire [62:0] _22610;
    wire [63:0] _22618;
    wire [62:0] _22619;
    wire [63:0] _22627;
    wire [62:0] _22628;
    wire [63:0] _22636;
    wire [62:0] _22637;
    wire [63:0] _22645;
    wire [62:0] _22646;
    wire [63:0] _22654;
    wire [62:0] _22655;
    wire [63:0] _22663;
    wire [62:0] _22664;
    wire [63:0] _22672;
    wire [62:0] _22673;
    wire [63:0] _22681;
    wire [62:0] _22682;
    wire [63:0] _22690;
    wire [62:0] _22691;
    wire [63:0] _22699;
    wire [62:0] _22700;
    wire [63:0] _22708;
    wire [62:0] _22709;
    wire [63:0] _22717;
    wire [62:0] _22718;
    wire [63:0] _22726;
    wire [62:0] _22727;
    wire [63:0] _22735;
    wire [62:0] _22736;
    wire [63:0] _22744;
    wire [62:0] _22745;
    wire [63:0] _22753;
    wire [62:0] _22754;
    wire [63:0] _22762;
    wire [127:0] _22763;
    wire [63:0] _22764;
    wire _22175;
    wire [63:0] _22172;
    wire [63:0] _22173;
    wire [62:0] _22174;
    wire [63:0] _22176;
    wire _22177;
    wire _22178;
    wire _22166;
    wire [63:0] _22163;
    wire [63:0] _22164;
    wire [62:0] _22165;
    wire [63:0] _22167;
    wire _22168;
    wire _22169;
    wire _22157;
    wire [63:0] _22154;
    wire [63:0] _22155;
    wire [62:0] _22156;
    wire [63:0] _22158;
    wire _22159;
    wire _22160;
    wire _22148;
    wire [63:0] _22145;
    wire [63:0] _22146;
    wire [62:0] _22147;
    wire [63:0] _22149;
    wire _22150;
    wire _22151;
    wire _22139;
    wire [63:0] _22136;
    wire [63:0] _22137;
    wire [62:0] _22138;
    wire [63:0] _22140;
    wire _22141;
    wire _22142;
    wire _22130;
    wire [63:0] _22127;
    wire [63:0] _22128;
    wire [62:0] _22129;
    wire [63:0] _22131;
    wire _22132;
    wire _22133;
    wire _22121;
    wire [63:0] _22118;
    wire [63:0] _22119;
    wire [62:0] _22120;
    wire [63:0] _22122;
    wire _22123;
    wire _22124;
    wire _22112;
    wire [63:0] _22109;
    wire [63:0] _22110;
    wire [62:0] _22111;
    wire [63:0] _22113;
    wire _22114;
    wire _22115;
    wire _22103;
    wire [63:0] _22100;
    wire [63:0] _22101;
    wire [62:0] _22102;
    wire [63:0] _22104;
    wire _22105;
    wire _22106;
    wire _22094;
    wire [63:0] _22091;
    wire [63:0] _22092;
    wire [62:0] _22093;
    wire [63:0] _22095;
    wire _22096;
    wire _22097;
    wire _22085;
    wire [63:0] _22082;
    wire [63:0] _22083;
    wire [62:0] _22084;
    wire [63:0] _22086;
    wire _22087;
    wire _22088;
    wire _22076;
    wire [63:0] _22073;
    wire [63:0] _22074;
    wire [62:0] _22075;
    wire [63:0] _22077;
    wire _22078;
    wire _22079;
    wire _22067;
    wire [63:0] _22064;
    wire [63:0] _22065;
    wire [62:0] _22066;
    wire [63:0] _22068;
    wire _22069;
    wire _22070;
    wire _22058;
    wire [63:0] _22055;
    wire [63:0] _22056;
    wire [62:0] _22057;
    wire [63:0] _22059;
    wire _22060;
    wire _22061;
    wire _22049;
    wire [63:0] _22046;
    wire [63:0] _22047;
    wire [62:0] _22048;
    wire [63:0] _22050;
    wire _22051;
    wire _22052;
    wire _22040;
    wire [63:0] _22037;
    wire [63:0] _22038;
    wire [62:0] _22039;
    wire [63:0] _22041;
    wire _22042;
    wire _22043;
    wire _22031;
    wire [63:0] _22028;
    wire [63:0] _22029;
    wire [62:0] _22030;
    wire [63:0] _22032;
    wire _22033;
    wire _22034;
    wire _22022;
    wire [63:0] _22019;
    wire [63:0] _22020;
    wire [62:0] _22021;
    wire [63:0] _22023;
    wire _22024;
    wire _22025;
    wire _22013;
    wire [63:0] _22010;
    wire [63:0] _22011;
    wire [62:0] _22012;
    wire [63:0] _22014;
    wire _22015;
    wire _22016;
    wire _22004;
    wire [63:0] _22001;
    wire [63:0] _22002;
    wire [62:0] _22003;
    wire [63:0] _22005;
    wire _22006;
    wire _22007;
    wire _21995;
    wire [63:0] _21992;
    wire [63:0] _21993;
    wire [62:0] _21994;
    wire [63:0] _21996;
    wire _21997;
    wire _21998;
    wire _21986;
    wire [63:0] _21983;
    wire [63:0] _21984;
    wire [62:0] _21985;
    wire [63:0] _21987;
    wire _21988;
    wire _21989;
    wire _21977;
    wire [63:0] _21974;
    wire [63:0] _21975;
    wire [62:0] _21976;
    wire [63:0] _21978;
    wire _21979;
    wire _21980;
    wire _21968;
    wire [63:0] _21965;
    wire [63:0] _21966;
    wire [62:0] _21967;
    wire [63:0] _21969;
    wire _21970;
    wire _21971;
    wire _21959;
    wire [63:0] _21956;
    wire [63:0] _21957;
    wire [62:0] _21958;
    wire [63:0] _21960;
    wire _21961;
    wire _21962;
    wire _21950;
    wire [63:0] _21947;
    wire [63:0] _21948;
    wire [62:0] _21949;
    wire [63:0] _21951;
    wire _21952;
    wire _21953;
    wire _21941;
    wire [63:0] _21938;
    wire [63:0] _21939;
    wire [62:0] _21940;
    wire [63:0] _21942;
    wire _21943;
    wire _21944;
    wire _21932;
    wire [63:0] _21929;
    wire [63:0] _21930;
    wire [62:0] _21931;
    wire [63:0] _21933;
    wire _21934;
    wire _21935;
    wire _21923;
    wire [63:0] _21920;
    wire [63:0] _21921;
    wire [62:0] _21922;
    wire [63:0] _21924;
    wire _21925;
    wire _21926;
    wire _21914;
    wire [63:0] _21911;
    wire [63:0] _21912;
    wire [62:0] _21913;
    wire [63:0] _21915;
    wire _21916;
    wire _21917;
    wire _21905;
    wire [63:0] _21902;
    wire [63:0] _21903;
    wire [62:0] _21904;
    wire [63:0] _21906;
    wire _21907;
    wire _21908;
    wire _21896;
    wire [63:0] _21893;
    wire [63:0] _21894;
    wire [62:0] _21895;
    wire [63:0] _21897;
    wire _21898;
    wire _21899;
    wire _21887;
    wire [63:0] _21884;
    wire [63:0] _21885;
    wire [62:0] _21886;
    wire [63:0] _21888;
    wire _21889;
    wire _21890;
    wire _21878;
    wire [63:0] _21875;
    wire [63:0] _21876;
    wire [62:0] _21877;
    wire [63:0] _21879;
    wire _21880;
    wire _21881;
    wire _21869;
    wire [63:0] _21866;
    wire [63:0] _21867;
    wire [62:0] _21868;
    wire [63:0] _21870;
    wire _21871;
    wire _21872;
    wire _21860;
    wire [63:0] _21857;
    wire [63:0] _21858;
    wire [62:0] _21859;
    wire [63:0] _21861;
    wire _21862;
    wire _21863;
    wire _21851;
    wire [63:0] _21848;
    wire [63:0] _21849;
    wire [62:0] _21850;
    wire [63:0] _21852;
    wire _21853;
    wire _21854;
    wire _21842;
    wire [63:0] _21839;
    wire [63:0] _21840;
    wire [62:0] _21841;
    wire [63:0] _21843;
    wire _21844;
    wire _21845;
    wire _21833;
    wire [63:0] _21830;
    wire [63:0] _21831;
    wire [62:0] _21832;
    wire [63:0] _21834;
    wire _21835;
    wire _21836;
    wire _21824;
    wire [63:0] _21821;
    wire [63:0] _21822;
    wire [62:0] _21823;
    wire [63:0] _21825;
    wire _21826;
    wire _21827;
    wire _21815;
    wire [63:0] _21812;
    wire [63:0] _21813;
    wire [62:0] _21814;
    wire [63:0] _21816;
    wire _21817;
    wire _21818;
    wire _21806;
    wire [63:0] _21803;
    wire [63:0] _21804;
    wire [62:0] _21805;
    wire [63:0] _21807;
    wire _21808;
    wire _21809;
    wire _21797;
    wire [63:0] _21794;
    wire [63:0] _21795;
    wire [62:0] _21796;
    wire [63:0] _21798;
    wire _21799;
    wire _21800;
    wire _21788;
    wire [63:0] _21785;
    wire [63:0] _21786;
    wire [62:0] _21787;
    wire [63:0] _21789;
    wire _21790;
    wire _21791;
    wire _21779;
    wire [63:0] _21776;
    wire [63:0] _21777;
    wire [62:0] _21778;
    wire [63:0] _21780;
    wire _21781;
    wire _21782;
    wire _21770;
    wire [63:0] _21767;
    wire [63:0] _21768;
    wire [62:0] _21769;
    wire [63:0] _21771;
    wire _21772;
    wire _21773;
    wire _21761;
    wire [63:0] _21758;
    wire [63:0] _21759;
    wire [62:0] _21760;
    wire [63:0] _21762;
    wire _21763;
    wire _21764;
    wire _21752;
    wire [63:0] _21749;
    wire [63:0] _21750;
    wire [62:0] _21751;
    wire [63:0] _21753;
    wire _21754;
    wire _21755;
    wire _21743;
    wire [63:0] _21740;
    wire [63:0] _21741;
    wire [62:0] _21742;
    wire [63:0] _21744;
    wire _21745;
    wire _21746;
    wire _21734;
    wire [63:0] _21731;
    wire [63:0] _21732;
    wire [62:0] _21733;
    wire [63:0] _21735;
    wire _21736;
    wire _21737;
    wire _21725;
    wire [63:0] _21722;
    wire [63:0] _21723;
    wire [62:0] _21724;
    wire [63:0] _21726;
    wire _21727;
    wire _21728;
    wire _21716;
    wire [63:0] _21713;
    wire [63:0] _21714;
    wire [62:0] _21715;
    wire [63:0] _21717;
    wire _21718;
    wire _21719;
    wire _21707;
    wire [63:0] _21704;
    wire [63:0] _21705;
    wire [62:0] _21706;
    wire [63:0] _21708;
    wire _21709;
    wire _21710;
    wire _21698;
    wire [63:0] _21695;
    wire [63:0] _21696;
    wire [62:0] _21697;
    wire [63:0] _21699;
    wire _21700;
    wire _21701;
    wire _21689;
    wire [63:0] _21686;
    wire [63:0] _21687;
    wire [62:0] _21688;
    wire [63:0] _21690;
    wire _21691;
    wire _21692;
    wire _21680;
    wire [63:0] _21677;
    wire [63:0] _21678;
    wire [62:0] _21679;
    wire [63:0] _21681;
    wire _21682;
    wire _21683;
    wire _21671;
    wire [63:0] _21668;
    wire [63:0] _21669;
    wire [62:0] _21670;
    wire [63:0] _21672;
    wire _21673;
    wire _21674;
    wire _21662;
    wire [63:0] _21659;
    wire [63:0] _21660;
    wire [62:0] _21661;
    wire [63:0] _21663;
    wire _21664;
    wire _21665;
    wire _21653;
    wire [63:0] _21650;
    wire [63:0] _21651;
    wire [62:0] _21652;
    wire [63:0] _21654;
    wire _21655;
    wire _21656;
    wire _21644;
    wire [63:0] _21641;
    wire [63:0] _21642;
    wire [62:0] _21643;
    wire [63:0] _21645;
    wire _21646;
    wire _21647;
    wire _21635;
    wire [63:0] _21632;
    wire [63:0] _21633;
    wire [62:0] _21634;
    wire [63:0] _21636;
    wire _21637;
    wire _21638;
    wire _21626;
    wire [63:0] _21623;
    wire [63:0] _21624;
    wire [62:0] _21625;
    wire [63:0] _21627;
    wire _21628;
    wire _21629;
    wire _21617;
    wire [63:0] _21614;
    wire [63:0] _21615;
    wire [62:0] _21616;
    wire [63:0] _21618;
    wire _21619;
    wire _21620;
    wire [63:0] _21607;
    wire _21608;
    wire [63:0] _21609;
    wire _21610;
    wire _21611;
    wire [63:0] _21612;
    wire [62:0] _21613;
    wire [63:0] _21621;
    wire [62:0] _21622;
    wire [63:0] _21630;
    wire [62:0] _21631;
    wire [63:0] _21639;
    wire [62:0] _21640;
    wire [63:0] _21648;
    wire [62:0] _21649;
    wire [63:0] _21657;
    wire [62:0] _21658;
    wire [63:0] _21666;
    wire [62:0] _21667;
    wire [63:0] _21675;
    wire [62:0] _21676;
    wire [63:0] _21684;
    wire [62:0] _21685;
    wire [63:0] _21693;
    wire [62:0] _21694;
    wire [63:0] _21702;
    wire [62:0] _21703;
    wire [63:0] _21711;
    wire [62:0] _21712;
    wire [63:0] _21720;
    wire [62:0] _21721;
    wire [63:0] _21729;
    wire [62:0] _21730;
    wire [63:0] _21738;
    wire [62:0] _21739;
    wire [63:0] _21747;
    wire [62:0] _21748;
    wire [63:0] _21756;
    wire [62:0] _21757;
    wire [63:0] _21765;
    wire [62:0] _21766;
    wire [63:0] _21774;
    wire [62:0] _21775;
    wire [63:0] _21783;
    wire [62:0] _21784;
    wire [63:0] _21792;
    wire [62:0] _21793;
    wire [63:0] _21801;
    wire [62:0] _21802;
    wire [63:0] _21810;
    wire [62:0] _21811;
    wire [63:0] _21819;
    wire [62:0] _21820;
    wire [63:0] _21828;
    wire [62:0] _21829;
    wire [63:0] _21837;
    wire [62:0] _21838;
    wire [63:0] _21846;
    wire [62:0] _21847;
    wire [63:0] _21855;
    wire [62:0] _21856;
    wire [63:0] _21864;
    wire [62:0] _21865;
    wire [63:0] _21873;
    wire [62:0] _21874;
    wire [63:0] _21882;
    wire [62:0] _21883;
    wire [63:0] _21891;
    wire [62:0] _21892;
    wire [63:0] _21900;
    wire [62:0] _21901;
    wire [63:0] _21909;
    wire [62:0] _21910;
    wire [63:0] _21918;
    wire [62:0] _21919;
    wire [63:0] _21927;
    wire [62:0] _21928;
    wire [63:0] _21936;
    wire [62:0] _21937;
    wire [63:0] _21945;
    wire [62:0] _21946;
    wire [63:0] _21954;
    wire [62:0] _21955;
    wire [63:0] _21963;
    wire [62:0] _21964;
    wire [63:0] _21972;
    wire [62:0] _21973;
    wire [63:0] _21981;
    wire [62:0] _21982;
    wire [63:0] _21990;
    wire [62:0] _21991;
    wire [63:0] _21999;
    wire [62:0] _22000;
    wire [63:0] _22008;
    wire [62:0] _22009;
    wire [63:0] _22017;
    wire [62:0] _22018;
    wire [63:0] _22026;
    wire [62:0] _22027;
    wire [63:0] _22035;
    wire [62:0] _22036;
    wire [63:0] _22044;
    wire [62:0] _22045;
    wire [63:0] _22053;
    wire [62:0] _22054;
    wire [63:0] _22062;
    wire [62:0] _22063;
    wire [63:0] _22071;
    wire [62:0] _22072;
    wire [63:0] _22080;
    wire [62:0] _22081;
    wire [63:0] _22089;
    wire [62:0] _22090;
    wire [63:0] _22098;
    wire [62:0] _22099;
    wire [63:0] _22107;
    wire [62:0] _22108;
    wire [63:0] _22116;
    wire [62:0] _22117;
    wire [63:0] _22125;
    wire [62:0] _22126;
    wire [63:0] _22134;
    wire [62:0] _22135;
    wire [63:0] _22143;
    wire [62:0] _22144;
    wire [63:0] _22152;
    wire [62:0] _22153;
    wire [63:0] _22161;
    wire [62:0] _22162;
    wire [63:0] _22170;
    wire [62:0] _22171;
    wire [63:0] _22179;
    wire [63:0] _22181;
    wire [127:0] _22182;
    wire [63:0] _22183;
    wire [63:0] _22765;
    wire [63:0] _21604;
    wire _21593;
    wire [63:0] _21590;
    wire [63:0] _21591;
    wire [62:0] _21592;
    wire [63:0] _21594;
    wire _21595;
    wire _21596;
    wire _21584;
    wire [63:0] _21581;
    wire [63:0] _21582;
    wire [62:0] _21583;
    wire [63:0] _21585;
    wire _21586;
    wire _21587;
    wire _21575;
    wire [63:0] _21572;
    wire [63:0] _21573;
    wire [62:0] _21574;
    wire [63:0] _21576;
    wire _21577;
    wire _21578;
    wire _21566;
    wire [63:0] _21563;
    wire [63:0] _21564;
    wire [62:0] _21565;
    wire [63:0] _21567;
    wire _21568;
    wire _21569;
    wire _21557;
    wire [63:0] _21554;
    wire [63:0] _21555;
    wire [62:0] _21556;
    wire [63:0] _21558;
    wire _21559;
    wire _21560;
    wire _21548;
    wire [63:0] _21545;
    wire [63:0] _21546;
    wire [62:0] _21547;
    wire [63:0] _21549;
    wire _21550;
    wire _21551;
    wire _21539;
    wire [63:0] _21536;
    wire [63:0] _21537;
    wire [62:0] _21538;
    wire [63:0] _21540;
    wire _21541;
    wire _21542;
    wire _21530;
    wire [63:0] _21527;
    wire [63:0] _21528;
    wire [62:0] _21529;
    wire [63:0] _21531;
    wire _21532;
    wire _21533;
    wire _21521;
    wire [63:0] _21518;
    wire [63:0] _21519;
    wire [62:0] _21520;
    wire [63:0] _21522;
    wire _21523;
    wire _21524;
    wire _21512;
    wire [63:0] _21509;
    wire [63:0] _21510;
    wire [62:0] _21511;
    wire [63:0] _21513;
    wire _21514;
    wire _21515;
    wire _21503;
    wire [63:0] _21500;
    wire [63:0] _21501;
    wire [62:0] _21502;
    wire [63:0] _21504;
    wire _21505;
    wire _21506;
    wire _21494;
    wire [63:0] _21491;
    wire [63:0] _21492;
    wire [62:0] _21493;
    wire [63:0] _21495;
    wire _21496;
    wire _21497;
    wire _21485;
    wire [63:0] _21482;
    wire [63:0] _21483;
    wire [62:0] _21484;
    wire [63:0] _21486;
    wire _21487;
    wire _21488;
    wire _21476;
    wire [63:0] _21473;
    wire [63:0] _21474;
    wire [62:0] _21475;
    wire [63:0] _21477;
    wire _21478;
    wire _21479;
    wire _21467;
    wire [63:0] _21464;
    wire [63:0] _21465;
    wire [62:0] _21466;
    wire [63:0] _21468;
    wire _21469;
    wire _21470;
    wire _21458;
    wire [63:0] _21455;
    wire [63:0] _21456;
    wire [62:0] _21457;
    wire [63:0] _21459;
    wire _21460;
    wire _21461;
    wire _21449;
    wire [63:0] _21446;
    wire [63:0] _21447;
    wire [62:0] _21448;
    wire [63:0] _21450;
    wire _21451;
    wire _21452;
    wire _21440;
    wire [63:0] _21437;
    wire [63:0] _21438;
    wire [62:0] _21439;
    wire [63:0] _21441;
    wire _21442;
    wire _21443;
    wire _21431;
    wire [63:0] _21428;
    wire [63:0] _21429;
    wire [62:0] _21430;
    wire [63:0] _21432;
    wire _21433;
    wire _21434;
    wire _21422;
    wire [63:0] _21419;
    wire [63:0] _21420;
    wire [62:0] _21421;
    wire [63:0] _21423;
    wire _21424;
    wire _21425;
    wire _21413;
    wire [63:0] _21410;
    wire [63:0] _21411;
    wire [62:0] _21412;
    wire [63:0] _21414;
    wire _21415;
    wire _21416;
    wire _21404;
    wire [63:0] _21401;
    wire [63:0] _21402;
    wire [62:0] _21403;
    wire [63:0] _21405;
    wire _21406;
    wire _21407;
    wire _21395;
    wire [63:0] _21392;
    wire [63:0] _21393;
    wire [62:0] _21394;
    wire [63:0] _21396;
    wire _21397;
    wire _21398;
    wire _21386;
    wire [63:0] _21383;
    wire [63:0] _21384;
    wire [62:0] _21385;
    wire [63:0] _21387;
    wire _21388;
    wire _21389;
    wire _21377;
    wire [63:0] _21374;
    wire [63:0] _21375;
    wire [62:0] _21376;
    wire [63:0] _21378;
    wire _21379;
    wire _21380;
    wire _21368;
    wire [63:0] _21365;
    wire [63:0] _21366;
    wire [62:0] _21367;
    wire [63:0] _21369;
    wire _21370;
    wire _21371;
    wire _21359;
    wire [63:0] _21356;
    wire [63:0] _21357;
    wire [62:0] _21358;
    wire [63:0] _21360;
    wire _21361;
    wire _21362;
    wire _21350;
    wire [63:0] _21347;
    wire [63:0] _21348;
    wire [62:0] _21349;
    wire [63:0] _21351;
    wire _21352;
    wire _21353;
    wire _21341;
    wire [63:0] _21338;
    wire [63:0] _21339;
    wire [62:0] _21340;
    wire [63:0] _21342;
    wire _21343;
    wire _21344;
    wire _21332;
    wire [63:0] _21329;
    wire [63:0] _21330;
    wire [62:0] _21331;
    wire [63:0] _21333;
    wire _21334;
    wire _21335;
    wire _21323;
    wire [63:0] _21320;
    wire [63:0] _21321;
    wire [62:0] _21322;
    wire [63:0] _21324;
    wire _21325;
    wire _21326;
    wire _21314;
    wire [63:0] _21311;
    wire [63:0] _21312;
    wire [62:0] _21313;
    wire [63:0] _21315;
    wire _21316;
    wire _21317;
    wire _21305;
    wire [63:0] _21302;
    wire [63:0] _21303;
    wire [62:0] _21304;
    wire [63:0] _21306;
    wire _21307;
    wire _21308;
    wire _21296;
    wire [63:0] _21293;
    wire [63:0] _21294;
    wire [62:0] _21295;
    wire [63:0] _21297;
    wire _21298;
    wire _21299;
    wire _21287;
    wire [63:0] _21284;
    wire [63:0] _21285;
    wire [62:0] _21286;
    wire [63:0] _21288;
    wire _21289;
    wire _21290;
    wire _21278;
    wire [63:0] _21275;
    wire [63:0] _21276;
    wire [62:0] _21277;
    wire [63:0] _21279;
    wire _21280;
    wire _21281;
    wire _21269;
    wire [63:0] _21266;
    wire [63:0] _21267;
    wire [62:0] _21268;
    wire [63:0] _21270;
    wire _21271;
    wire _21272;
    wire _21260;
    wire [63:0] _21257;
    wire [63:0] _21258;
    wire [62:0] _21259;
    wire [63:0] _21261;
    wire _21262;
    wire _21263;
    wire _21251;
    wire [63:0] _21248;
    wire [63:0] _21249;
    wire [62:0] _21250;
    wire [63:0] _21252;
    wire _21253;
    wire _21254;
    wire _21242;
    wire [63:0] _21239;
    wire [63:0] _21240;
    wire [62:0] _21241;
    wire [63:0] _21243;
    wire _21244;
    wire _21245;
    wire _21233;
    wire [63:0] _21230;
    wire [63:0] _21231;
    wire [62:0] _21232;
    wire [63:0] _21234;
    wire _21235;
    wire _21236;
    wire _21224;
    wire [63:0] _21221;
    wire [63:0] _21222;
    wire [62:0] _21223;
    wire [63:0] _21225;
    wire _21226;
    wire _21227;
    wire _21215;
    wire [63:0] _21212;
    wire [63:0] _21213;
    wire [62:0] _21214;
    wire [63:0] _21216;
    wire _21217;
    wire _21218;
    wire _21206;
    wire [63:0] _21203;
    wire [63:0] _21204;
    wire [62:0] _21205;
    wire [63:0] _21207;
    wire _21208;
    wire _21209;
    wire _21197;
    wire [63:0] _21194;
    wire [63:0] _21195;
    wire [62:0] _21196;
    wire [63:0] _21198;
    wire _21199;
    wire _21200;
    wire _21188;
    wire [63:0] _21185;
    wire [63:0] _21186;
    wire [62:0] _21187;
    wire [63:0] _21189;
    wire _21190;
    wire _21191;
    wire _21179;
    wire [63:0] _21176;
    wire [63:0] _21177;
    wire [62:0] _21178;
    wire [63:0] _21180;
    wire _21181;
    wire _21182;
    wire _21170;
    wire [63:0] _21167;
    wire [63:0] _21168;
    wire [62:0] _21169;
    wire [63:0] _21171;
    wire _21172;
    wire _21173;
    wire _21161;
    wire [63:0] _21158;
    wire [63:0] _21159;
    wire [62:0] _21160;
    wire [63:0] _21162;
    wire _21163;
    wire _21164;
    wire _21152;
    wire [63:0] _21149;
    wire [63:0] _21150;
    wire [62:0] _21151;
    wire [63:0] _21153;
    wire _21154;
    wire _21155;
    wire _21143;
    wire [63:0] _21140;
    wire [63:0] _21141;
    wire [62:0] _21142;
    wire [63:0] _21144;
    wire _21145;
    wire _21146;
    wire _21134;
    wire [63:0] _21131;
    wire [63:0] _21132;
    wire [62:0] _21133;
    wire [63:0] _21135;
    wire _21136;
    wire _21137;
    wire _21125;
    wire [63:0] _21122;
    wire [63:0] _21123;
    wire [62:0] _21124;
    wire [63:0] _21126;
    wire _21127;
    wire _21128;
    wire _21116;
    wire [63:0] _21113;
    wire [63:0] _21114;
    wire [62:0] _21115;
    wire [63:0] _21117;
    wire _21118;
    wire _21119;
    wire _21107;
    wire [63:0] _21104;
    wire [63:0] _21105;
    wire [62:0] _21106;
    wire [63:0] _21108;
    wire _21109;
    wire _21110;
    wire _21098;
    wire [63:0] _21095;
    wire [63:0] _21096;
    wire [62:0] _21097;
    wire [63:0] _21099;
    wire _21100;
    wire _21101;
    wire _21089;
    wire [63:0] _21086;
    wire [63:0] _21087;
    wire [62:0] _21088;
    wire [63:0] _21090;
    wire _21091;
    wire _21092;
    wire _21080;
    wire [63:0] _21077;
    wire [63:0] _21078;
    wire [62:0] _21079;
    wire [63:0] _21081;
    wire _21082;
    wire _21083;
    wire _21071;
    wire [63:0] _21068;
    wire [63:0] _21069;
    wire [62:0] _21070;
    wire [63:0] _21072;
    wire _21073;
    wire _21074;
    wire _21062;
    wire [63:0] _21059;
    wire [63:0] _21060;
    wire [62:0] _21061;
    wire [63:0] _21063;
    wire _21064;
    wire _21065;
    wire _21053;
    wire [63:0] _21050;
    wire [63:0] _21051;
    wire [62:0] _21052;
    wire [63:0] _21054;
    wire _21055;
    wire _21056;
    wire _21044;
    wire [63:0] _21041;
    wire [63:0] _21042;
    wire [62:0] _21043;
    wire [63:0] _21045;
    wire _21046;
    wire _21047;
    wire _21035;
    wire [63:0] _21032;
    wire [63:0] _21033;
    wire [62:0] _21034;
    wire [63:0] _21036;
    wire _21037;
    wire _21038;
    wire [63:0] _21027;
    wire [63:0] _21023;
    wire [63:0] _21024;
    wire _21025;
    wire [63:0] _21026;
    wire _21028;
    wire _21029;
    wire [63:0] _21030;
    wire [62:0] _21031;
    wire [63:0] _21039;
    wire [62:0] _21040;
    wire [63:0] _21048;
    wire [62:0] _21049;
    wire [63:0] _21057;
    wire [62:0] _21058;
    wire [63:0] _21066;
    wire [62:0] _21067;
    wire [63:0] _21075;
    wire [62:0] _21076;
    wire [63:0] _21084;
    wire [62:0] _21085;
    wire [63:0] _21093;
    wire [62:0] _21094;
    wire [63:0] _21102;
    wire [62:0] _21103;
    wire [63:0] _21111;
    wire [62:0] _21112;
    wire [63:0] _21120;
    wire [62:0] _21121;
    wire [63:0] _21129;
    wire [62:0] _21130;
    wire [63:0] _21138;
    wire [62:0] _21139;
    wire [63:0] _21147;
    wire [62:0] _21148;
    wire [63:0] _21156;
    wire [62:0] _21157;
    wire [63:0] _21165;
    wire [62:0] _21166;
    wire [63:0] _21174;
    wire [62:0] _21175;
    wire [63:0] _21183;
    wire [62:0] _21184;
    wire [63:0] _21192;
    wire [62:0] _21193;
    wire [63:0] _21201;
    wire [62:0] _21202;
    wire [63:0] _21210;
    wire [62:0] _21211;
    wire [63:0] _21219;
    wire [62:0] _21220;
    wire [63:0] _21228;
    wire [62:0] _21229;
    wire [63:0] _21237;
    wire [62:0] _21238;
    wire [63:0] _21246;
    wire [62:0] _21247;
    wire [63:0] _21255;
    wire [62:0] _21256;
    wire [63:0] _21264;
    wire [62:0] _21265;
    wire [63:0] _21273;
    wire [62:0] _21274;
    wire [63:0] _21282;
    wire [62:0] _21283;
    wire [63:0] _21291;
    wire [62:0] _21292;
    wire [63:0] _21300;
    wire [62:0] _21301;
    wire [63:0] _21309;
    wire [62:0] _21310;
    wire [63:0] _21318;
    wire [62:0] _21319;
    wire [63:0] _21327;
    wire [62:0] _21328;
    wire [63:0] _21336;
    wire [62:0] _21337;
    wire [63:0] _21345;
    wire [62:0] _21346;
    wire [63:0] _21354;
    wire [62:0] _21355;
    wire [63:0] _21363;
    wire [62:0] _21364;
    wire [63:0] _21372;
    wire [62:0] _21373;
    wire [63:0] _21381;
    wire [62:0] _21382;
    wire [63:0] _21390;
    wire [62:0] _21391;
    wire [63:0] _21399;
    wire [62:0] _21400;
    wire [63:0] _21408;
    wire [62:0] _21409;
    wire [63:0] _21417;
    wire [62:0] _21418;
    wire [63:0] _21426;
    wire [62:0] _21427;
    wire [63:0] _21435;
    wire [62:0] _21436;
    wire [63:0] _21444;
    wire [62:0] _21445;
    wire [63:0] _21453;
    wire [62:0] _21454;
    wire [63:0] _21462;
    wire [62:0] _21463;
    wire [63:0] _21471;
    wire [62:0] _21472;
    wire [63:0] _21480;
    wire [62:0] _21481;
    wire [63:0] _21489;
    wire [62:0] _21490;
    wire [63:0] _21498;
    wire [62:0] _21499;
    wire [63:0] _21507;
    wire [62:0] _21508;
    wire [63:0] _21516;
    wire [62:0] _21517;
    wire [63:0] _21525;
    wire [62:0] _21526;
    wire [63:0] _21534;
    wire [62:0] _21535;
    wire [63:0] _21543;
    wire [62:0] _21544;
    wire [63:0] _21552;
    wire [62:0] _21553;
    wire [63:0] _21561;
    wire [62:0] _21562;
    wire [63:0] _21570;
    wire [62:0] _21571;
    wire [63:0] _21579;
    wire [62:0] _21580;
    wire [63:0] _21588;
    wire [62:0] _21589;
    wire [63:0] _21597;
    wire [127:0] _21598;
    wire [63:0] _21599;
    wire _21600;
    wire [63:0] _21601;
    wire [63:0] _21017;
    wire _21018;
    wire [63:0] _21019;
    wire _21602;
    wire _21603;
    wire [63:0] _22766;
    wire _21008;
    wire [63:0] _21005;
    wire [63:0] _21006;
    wire [62:0] _21007;
    wire [63:0] _21009;
    wire _21010;
    wire _21011;
    wire _20999;
    wire [63:0] _20996;
    wire [63:0] _20997;
    wire [62:0] _20998;
    wire [63:0] _21000;
    wire _21001;
    wire _21002;
    wire _20990;
    wire [63:0] _20987;
    wire [63:0] _20988;
    wire [62:0] _20989;
    wire [63:0] _20991;
    wire _20992;
    wire _20993;
    wire _20981;
    wire [63:0] _20978;
    wire [63:0] _20979;
    wire [62:0] _20980;
    wire [63:0] _20982;
    wire _20983;
    wire _20984;
    wire _20972;
    wire [63:0] _20969;
    wire [63:0] _20970;
    wire [62:0] _20971;
    wire [63:0] _20973;
    wire _20974;
    wire _20975;
    wire _20963;
    wire [63:0] _20960;
    wire [63:0] _20961;
    wire [62:0] _20962;
    wire [63:0] _20964;
    wire _20965;
    wire _20966;
    wire _20954;
    wire [63:0] _20951;
    wire [63:0] _20952;
    wire [62:0] _20953;
    wire [63:0] _20955;
    wire _20956;
    wire _20957;
    wire _20945;
    wire [63:0] _20942;
    wire [63:0] _20943;
    wire [62:0] _20944;
    wire [63:0] _20946;
    wire _20947;
    wire _20948;
    wire _20936;
    wire [63:0] _20933;
    wire [63:0] _20934;
    wire [62:0] _20935;
    wire [63:0] _20937;
    wire _20938;
    wire _20939;
    wire _20927;
    wire [63:0] _20924;
    wire [63:0] _20925;
    wire [62:0] _20926;
    wire [63:0] _20928;
    wire _20929;
    wire _20930;
    wire _20918;
    wire [63:0] _20915;
    wire [63:0] _20916;
    wire [62:0] _20917;
    wire [63:0] _20919;
    wire _20920;
    wire _20921;
    wire _20909;
    wire [63:0] _20906;
    wire [63:0] _20907;
    wire [62:0] _20908;
    wire [63:0] _20910;
    wire _20911;
    wire _20912;
    wire _20900;
    wire [63:0] _20897;
    wire [63:0] _20898;
    wire [62:0] _20899;
    wire [63:0] _20901;
    wire _20902;
    wire _20903;
    wire _20891;
    wire [63:0] _20888;
    wire [63:0] _20889;
    wire [62:0] _20890;
    wire [63:0] _20892;
    wire _20893;
    wire _20894;
    wire _20882;
    wire [63:0] _20879;
    wire [63:0] _20880;
    wire [62:0] _20881;
    wire [63:0] _20883;
    wire _20884;
    wire _20885;
    wire _20873;
    wire [63:0] _20870;
    wire [63:0] _20871;
    wire [62:0] _20872;
    wire [63:0] _20874;
    wire _20875;
    wire _20876;
    wire _20864;
    wire [63:0] _20861;
    wire [63:0] _20862;
    wire [62:0] _20863;
    wire [63:0] _20865;
    wire _20866;
    wire _20867;
    wire _20855;
    wire [63:0] _20852;
    wire [63:0] _20853;
    wire [62:0] _20854;
    wire [63:0] _20856;
    wire _20857;
    wire _20858;
    wire _20846;
    wire [63:0] _20843;
    wire [63:0] _20844;
    wire [62:0] _20845;
    wire [63:0] _20847;
    wire _20848;
    wire _20849;
    wire _20837;
    wire [63:0] _20834;
    wire [63:0] _20835;
    wire [62:0] _20836;
    wire [63:0] _20838;
    wire _20839;
    wire _20840;
    wire _20828;
    wire [63:0] _20825;
    wire [63:0] _20826;
    wire [62:0] _20827;
    wire [63:0] _20829;
    wire _20830;
    wire _20831;
    wire _20819;
    wire [63:0] _20816;
    wire [63:0] _20817;
    wire [62:0] _20818;
    wire [63:0] _20820;
    wire _20821;
    wire _20822;
    wire _20810;
    wire [63:0] _20807;
    wire [63:0] _20808;
    wire [62:0] _20809;
    wire [63:0] _20811;
    wire _20812;
    wire _20813;
    wire _20801;
    wire [63:0] _20798;
    wire [63:0] _20799;
    wire [62:0] _20800;
    wire [63:0] _20802;
    wire _20803;
    wire _20804;
    wire _20792;
    wire [63:0] _20789;
    wire [63:0] _20790;
    wire [62:0] _20791;
    wire [63:0] _20793;
    wire _20794;
    wire _20795;
    wire _20783;
    wire [63:0] _20780;
    wire [63:0] _20781;
    wire [62:0] _20782;
    wire [63:0] _20784;
    wire _20785;
    wire _20786;
    wire _20774;
    wire [63:0] _20771;
    wire [63:0] _20772;
    wire [62:0] _20773;
    wire [63:0] _20775;
    wire _20776;
    wire _20777;
    wire _20765;
    wire [63:0] _20762;
    wire [63:0] _20763;
    wire [62:0] _20764;
    wire [63:0] _20766;
    wire _20767;
    wire _20768;
    wire _20756;
    wire [63:0] _20753;
    wire [63:0] _20754;
    wire [62:0] _20755;
    wire [63:0] _20757;
    wire _20758;
    wire _20759;
    wire _20747;
    wire [63:0] _20744;
    wire [63:0] _20745;
    wire [62:0] _20746;
    wire [63:0] _20748;
    wire _20749;
    wire _20750;
    wire _20738;
    wire [63:0] _20735;
    wire [63:0] _20736;
    wire [62:0] _20737;
    wire [63:0] _20739;
    wire _20740;
    wire _20741;
    wire _20729;
    wire [63:0] _20726;
    wire [63:0] _20727;
    wire [62:0] _20728;
    wire [63:0] _20730;
    wire _20731;
    wire _20732;
    wire _20720;
    wire [63:0] _20717;
    wire [63:0] _20718;
    wire [62:0] _20719;
    wire [63:0] _20721;
    wire _20722;
    wire _20723;
    wire _20711;
    wire [63:0] _20708;
    wire [63:0] _20709;
    wire [62:0] _20710;
    wire [63:0] _20712;
    wire _20713;
    wire _20714;
    wire _20702;
    wire [63:0] _20699;
    wire [63:0] _20700;
    wire [62:0] _20701;
    wire [63:0] _20703;
    wire _20704;
    wire _20705;
    wire _20693;
    wire [63:0] _20690;
    wire [63:0] _20691;
    wire [62:0] _20692;
    wire [63:0] _20694;
    wire _20695;
    wire _20696;
    wire _20684;
    wire [63:0] _20681;
    wire [63:0] _20682;
    wire [62:0] _20683;
    wire [63:0] _20685;
    wire _20686;
    wire _20687;
    wire _20675;
    wire [63:0] _20672;
    wire [63:0] _20673;
    wire [62:0] _20674;
    wire [63:0] _20676;
    wire _20677;
    wire _20678;
    wire _20666;
    wire [63:0] _20663;
    wire [63:0] _20664;
    wire [62:0] _20665;
    wire [63:0] _20667;
    wire _20668;
    wire _20669;
    wire _20657;
    wire [63:0] _20654;
    wire [63:0] _20655;
    wire [62:0] _20656;
    wire [63:0] _20658;
    wire _20659;
    wire _20660;
    wire _20648;
    wire [63:0] _20645;
    wire [63:0] _20646;
    wire [62:0] _20647;
    wire [63:0] _20649;
    wire _20650;
    wire _20651;
    wire _20639;
    wire [63:0] _20636;
    wire [63:0] _20637;
    wire [62:0] _20638;
    wire [63:0] _20640;
    wire _20641;
    wire _20642;
    wire _20630;
    wire [63:0] _20627;
    wire [63:0] _20628;
    wire [62:0] _20629;
    wire [63:0] _20631;
    wire _20632;
    wire _20633;
    wire _20621;
    wire [63:0] _20618;
    wire [63:0] _20619;
    wire [62:0] _20620;
    wire [63:0] _20622;
    wire _20623;
    wire _20624;
    wire _20612;
    wire [63:0] _20609;
    wire [63:0] _20610;
    wire [62:0] _20611;
    wire [63:0] _20613;
    wire _20614;
    wire _20615;
    wire _20603;
    wire [63:0] _20600;
    wire [63:0] _20601;
    wire [62:0] _20602;
    wire [63:0] _20604;
    wire _20605;
    wire _20606;
    wire _20594;
    wire [63:0] _20591;
    wire [63:0] _20592;
    wire [62:0] _20593;
    wire [63:0] _20595;
    wire _20596;
    wire _20597;
    wire _20585;
    wire [63:0] _20582;
    wire [63:0] _20583;
    wire [62:0] _20584;
    wire [63:0] _20586;
    wire _20587;
    wire _20588;
    wire _20576;
    wire [63:0] _20573;
    wire [63:0] _20574;
    wire [62:0] _20575;
    wire [63:0] _20577;
    wire _20578;
    wire _20579;
    wire _20567;
    wire [63:0] _20564;
    wire [63:0] _20565;
    wire [62:0] _20566;
    wire [63:0] _20568;
    wire _20569;
    wire _20570;
    wire _20558;
    wire [63:0] _20555;
    wire [63:0] _20556;
    wire [62:0] _20557;
    wire [63:0] _20559;
    wire _20560;
    wire _20561;
    wire _20549;
    wire [63:0] _20546;
    wire [63:0] _20547;
    wire [62:0] _20548;
    wire [63:0] _20550;
    wire _20551;
    wire _20552;
    wire _20540;
    wire [63:0] _20537;
    wire [63:0] _20538;
    wire [62:0] _20539;
    wire [63:0] _20541;
    wire _20542;
    wire _20543;
    wire _20531;
    wire [63:0] _20528;
    wire [63:0] _20529;
    wire [62:0] _20530;
    wire [63:0] _20532;
    wire _20533;
    wire _20534;
    wire _20522;
    wire [63:0] _20519;
    wire [63:0] _20520;
    wire [62:0] _20521;
    wire [63:0] _20523;
    wire _20524;
    wire _20525;
    wire _20513;
    wire [63:0] _20510;
    wire [63:0] _20511;
    wire [62:0] _20512;
    wire [63:0] _20514;
    wire _20515;
    wire _20516;
    wire _20504;
    wire [63:0] _20501;
    wire [63:0] _20502;
    wire [62:0] _20503;
    wire [63:0] _20505;
    wire _20506;
    wire _20507;
    wire _20495;
    wire [63:0] _20492;
    wire [63:0] _20493;
    wire [62:0] _20494;
    wire [63:0] _20496;
    wire _20497;
    wire _20498;
    wire _20486;
    wire [63:0] _20483;
    wire [63:0] _20484;
    wire [62:0] _20485;
    wire [63:0] _20487;
    wire _20488;
    wire _20489;
    wire _20477;
    wire [63:0] _20474;
    wire [63:0] _20475;
    wire [62:0] _20476;
    wire [63:0] _20478;
    wire _20479;
    wire _20480;
    wire _20468;
    wire [63:0] _20465;
    wire [63:0] _20466;
    wire [62:0] _20467;
    wire [63:0] _20469;
    wire _20470;
    wire _20471;
    wire _20459;
    wire [63:0] _20456;
    wire [63:0] _20457;
    wire [62:0] _20458;
    wire [63:0] _20460;
    wire _20461;
    wire _20462;
    wire _20450;
    wire [63:0] _20447;
    wire [63:0] _20448;
    wire [62:0] _20449;
    wire [63:0] _20451;
    wire _20452;
    wire _20453;
    wire [63:0] _20437;
    wire [127:0] _20438;
    wire [63:0] _20439;
    wire _20440;
    wire [63:0] _20441;
    wire _20443;
    wire _20444;
    wire [63:0] _20445;
    wire [62:0] _20446;
    wire [63:0] _20454;
    wire [62:0] _20455;
    wire [63:0] _20463;
    wire [62:0] _20464;
    wire [63:0] _20472;
    wire [62:0] _20473;
    wire [63:0] _20481;
    wire [62:0] _20482;
    wire [63:0] _20490;
    wire [62:0] _20491;
    wire [63:0] _20499;
    wire [62:0] _20500;
    wire [63:0] _20508;
    wire [62:0] _20509;
    wire [63:0] _20517;
    wire [62:0] _20518;
    wire [63:0] _20526;
    wire [62:0] _20527;
    wire [63:0] _20535;
    wire [62:0] _20536;
    wire [63:0] _20544;
    wire [62:0] _20545;
    wire [63:0] _20553;
    wire [62:0] _20554;
    wire [63:0] _20562;
    wire [62:0] _20563;
    wire [63:0] _20571;
    wire [62:0] _20572;
    wire [63:0] _20580;
    wire [62:0] _20581;
    wire [63:0] _20589;
    wire [62:0] _20590;
    wire [63:0] _20598;
    wire [62:0] _20599;
    wire [63:0] _20607;
    wire [62:0] _20608;
    wire [63:0] _20616;
    wire [62:0] _20617;
    wire [63:0] _20625;
    wire [62:0] _20626;
    wire [63:0] _20634;
    wire [62:0] _20635;
    wire [63:0] _20643;
    wire [62:0] _20644;
    wire [63:0] _20652;
    wire [62:0] _20653;
    wire [63:0] _20661;
    wire [62:0] _20662;
    wire [63:0] _20670;
    wire [62:0] _20671;
    wire [63:0] _20679;
    wire [62:0] _20680;
    wire [63:0] _20688;
    wire [62:0] _20689;
    wire [63:0] _20697;
    wire [62:0] _20698;
    wire [63:0] _20706;
    wire [62:0] _20707;
    wire [63:0] _20715;
    wire [62:0] _20716;
    wire [63:0] _20724;
    wire [62:0] _20725;
    wire [63:0] _20733;
    wire [62:0] _20734;
    wire [63:0] _20742;
    wire [62:0] _20743;
    wire [63:0] _20751;
    wire [62:0] _20752;
    wire [63:0] _20760;
    wire [62:0] _20761;
    wire [63:0] _20769;
    wire [62:0] _20770;
    wire [63:0] _20778;
    wire [62:0] _20779;
    wire [63:0] _20787;
    wire [62:0] _20788;
    wire [63:0] _20796;
    wire [62:0] _20797;
    wire [63:0] _20805;
    wire [62:0] _20806;
    wire [63:0] _20814;
    wire [62:0] _20815;
    wire [63:0] _20823;
    wire [62:0] _20824;
    wire [63:0] _20832;
    wire [62:0] _20833;
    wire [63:0] _20841;
    wire [62:0] _20842;
    wire [63:0] _20850;
    wire [62:0] _20851;
    wire [63:0] _20859;
    wire [62:0] _20860;
    wire [63:0] _20868;
    wire [62:0] _20869;
    wire [63:0] _20877;
    wire [62:0] _20878;
    wire [63:0] _20886;
    wire [62:0] _20887;
    wire [63:0] _20895;
    wire [62:0] _20896;
    wire [63:0] _20904;
    wire [62:0] _20905;
    wire [63:0] _20913;
    wire [62:0] _20914;
    wire [63:0] _20922;
    wire [62:0] _20923;
    wire [63:0] _20931;
    wire [62:0] _20932;
    wire [63:0] _20940;
    wire [62:0] _20941;
    wire [63:0] _20949;
    wire [62:0] _20950;
    wire [63:0] _20958;
    wire [62:0] _20959;
    wire [63:0] _20967;
    wire [62:0] _20968;
    wire [63:0] _20976;
    wire [62:0] _20977;
    wire [63:0] _20985;
    wire [62:0] _20986;
    wire [63:0] _20994;
    wire [62:0] _20995;
    wire [63:0] _21003;
    wire [62:0] _21004;
    wire [63:0] _21012;
    wire [127:0] _21013;
    wire [63:0] _21014;
    wire _20425;
    wire [63:0] _20422;
    wire [63:0] _20423;
    wire [62:0] _20424;
    wire [63:0] _20426;
    wire _20427;
    wire _20428;
    wire _20416;
    wire [63:0] _20413;
    wire [63:0] _20414;
    wire [62:0] _20415;
    wire [63:0] _20417;
    wire _20418;
    wire _20419;
    wire _20407;
    wire [63:0] _20404;
    wire [63:0] _20405;
    wire [62:0] _20406;
    wire [63:0] _20408;
    wire _20409;
    wire _20410;
    wire _20398;
    wire [63:0] _20395;
    wire [63:0] _20396;
    wire [62:0] _20397;
    wire [63:0] _20399;
    wire _20400;
    wire _20401;
    wire _20389;
    wire [63:0] _20386;
    wire [63:0] _20387;
    wire [62:0] _20388;
    wire [63:0] _20390;
    wire _20391;
    wire _20392;
    wire _20380;
    wire [63:0] _20377;
    wire [63:0] _20378;
    wire [62:0] _20379;
    wire [63:0] _20381;
    wire _20382;
    wire _20383;
    wire _20371;
    wire [63:0] _20368;
    wire [63:0] _20369;
    wire [62:0] _20370;
    wire [63:0] _20372;
    wire _20373;
    wire _20374;
    wire _20362;
    wire [63:0] _20359;
    wire [63:0] _20360;
    wire [62:0] _20361;
    wire [63:0] _20363;
    wire _20364;
    wire _20365;
    wire _20353;
    wire [63:0] _20350;
    wire [63:0] _20351;
    wire [62:0] _20352;
    wire [63:0] _20354;
    wire _20355;
    wire _20356;
    wire _20344;
    wire [63:0] _20341;
    wire [63:0] _20342;
    wire [62:0] _20343;
    wire [63:0] _20345;
    wire _20346;
    wire _20347;
    wire _20335;
    wire [63:0] _20332;
    wire [63:0] _20333;
    wire [62:0] _20334;
    wire [63:0] _20336;
    wire _20337;
    wire _20338;
    wire _20326;
    wire [63:0] _20323;
    wire [63:0] _20324;
    wire [62:0] _20325;
    wire [63:0] _20327;
    wire _20328;
    wire _20329;
    wire _20317;
    wire [63:0] _20314;
    wire [63:0] _20315;
    wire [62:0] _20316;
    wire [63:0] _20318;
    wire _20319;
    wire _20320;
    wire _20308;
    wire [63:0] _20305;
    wire [63:0] _20306;
    wire [62:0] _20307;
    wire [63:0] _20309;
    wire _20310;
    wire _20311;
    wire _20299;
    wire [63:0] _20296;
    wire [63:0] _20297;
    wire [62:0] _20298;
    wire [63:0] _20300;
    wire _20301;
    wire _20302;
    wire _20290;
    wire [63:0] _20287;
    wire [63:0] _20288;
    wire [62:0] _20289;
    wire [63:0] _20291;
    wire _20292;
    wire _20293;
    wire _20281;
    wire [63:0] _20278;
    wire [63:0] _20279;
    wire [62:0] _20280;
    wire [63:0] _20282;
    wire _20283;
    wire _20284;
    wire _20272;
    wire [63:0] _20269;
    wire [63:0] _20270;
    wire [62:0] _20271;
    wire [63:0] _20273;
    wire _20274;
    wire _20275;
    wire _20263;
    wire [63:0] _20260;
    wire [63:0] _20261;
    wire [62:0] _20262;
    wire [63:0] _20264;
    wire _20265;
    wire _20266;
    wire _20254;
    wire [63:0] _20251;
    wire [63:0] _20252;
    wire [62:0] _20253;
    wire [63:0] _20255;
    wire _20256;
    wire _20257;
    wire _20245;
    wire [63:0] _20242;
    wire [63:0] _20243;
    wire [62:0] _20244;
    wire [63:0] _20246;
    wire _20247;
    wire _20248;
    wire _20236;
    wire [63:0] _20233;
    wire [63:0] _20234;
    wire [62:0] _20235;
    wire [63:0] _20237;
    wire _20238;
    wire _20239;
    wire _20227;
    wire [63:0] _20224;
    wire [63:0] _20225;
    wire [62:0] _20226;
    wire [63:0] _20228;
    wire _20229;
    wire _20230;
    wire _20218;
    wire [63:0] _20215;
    wire [63:0] _20216;
    wire [62:0] _20217;
    wire [63:0] _20219;
    wire _20220;
    wire _20221;
    wire _20209;
    wire [63:0] _20206;
    wire [63:0] _20207;
    wire [62:0] _20208;
    wire [63:0] _20210;
    wire _20211;
    wire _20212;
    wire _20200;
    wire [63:0] _20197;
    wire [63:0] _20198;
    wire [62:0] _20199;
    wire [63:0] _20201;
    wire _20202;
    wire _20203;
    wire _20191;
    wire [63:0] _20188;
    wire [63:0] _20189;
    wire [62:0] _20190;
    wire [63:0] _20192;
    wire _20193;
    wire _20194;
    wire _20182;
    wire [63:0] _20179;
    wire [63:0] _20180;
    wire [62:0] _20181;
    wire [63:0] _20183;
    wire _20184;
    wire _20185;
    wire _20173;
    wire [63:0] _20170;
    wire [63:0] _20171;
    wire [62:0] _20172;
    wire [63:0] _20174;
    wire _20175;
    wire _20176;
    wire _20164;
    wire [63:0] _20161;
    wire [63:0] _20162;
    wire [62:0] _20163;
    wire [63:0] _20165;
    wire _20166;
    wire _20167;
    wire _20155;
    wire [63:0] _20152;
    wire [63:0] _20153;
    wire [62:0] _20154;
    wire [63:0] _20156;
    wire _20157;
    wire _20158;
    wire _20146;
    wire [63:0] _20143;
    wire [63:0] _20144;
    wire [62:0] _20145;
    wire [63:0] _20147;
    wire _20148;
    wire _20149;
    wire _20137;
    wire [63:0] _20134;
    wire [63:0] _20135;
    wire [62:0] _20136;
    wire [63:0] _20138;
    wire _20139;
    wire _20140;
    wire _20128;
    wire [63:0] _20125;
    wire [63:0] _20126;
    wire [62:0] _20127;
    wire [63:0] _20129;
    wire _20130;
    wire _20131;
    wire _20119;
    wire [63:0] _20116;
    wire [63:0] _20117;
    wire [62:0] _20118;
    wire [63:0] _20120;
    wire _20121;
    wire _20122;
    wire _20110;
    wire [63:0] _20107;
    wire [63:0] _20108;
    wire [62:0] _20109;
    wire [63:0] _20111;
    wire _20112;
    wire _20113;
    wire _20101;
    wire [63:0] _20098;
    wire [63:0] _20099;
    wire [62:0] _20100;
    wire [63:0] _20102;
    wire _20103;
    wire _20104;
    wire _20092;
    wire [63:0] _20089;
    wire [63:0] _20090;
    wire [62:0] _20091;
    wire [63:0] _20093;
    wire _20094;
    wire _20095;
    wire _20083;
    wire [63:0] _20080;
    wire [63:0] _20081;
    wire [62:0] _20082;
    wire [63:0] _20084;
    wire _20085;
    wire _20086;
    wire _20074;
    wire [63:0] _20071;
    wire [63:0] _20072;
    wire [62:0] _20073;
    wire [63:0] _20075;
    wire _20076;
    wire _20077;
    wire _20065;
    wire [63:0] _20062;
    wire [63:0] _20063;
    wire [62:0] _20064;
    wire [63:0] _20066;
    wire _20067;
    wire _20068;
    wire _20056;
    wire [63:0] _20053;
    wire [63:0] _20054;
    wire [62:0] _20055;
    wire [63:0] _20057;
    wire _20058;
    wire _20059;
    wire _20047;
    wire [63:0] _20044;
    wire [63:0] _20045;
    wire [62:0] _20046;
    wire [63:0] _20048;
    wire _20049;
    wire _20050;
    wire _20038;
    wire [63:0] _20035;
    wire [63:0] _20036;
    wire [62:0] _20037;
    wire [63:0] _20039;
    wire _20040;
    wire _20041;
    wire _20029;
    wire [63:0] _20026;
    wire [63:0] _20027;
    wire [62:0] _20028;
    wire [63:0] _20030;
    wire _20031;
    wire _20032;
    wire _20020;
    wire [63:0] _20017;
    wire [63:0] _20018;
    wire [62:0] _20019;
    wire [63:0] _20021;
    wire _20022;
    wire _20023;
    wire _20011;
    wire [63:0] _20008;
    wire [63:0] _20009;
    wire [62:0] _20010;
    wire [63:0] _20012;
    wire _20013;
    wire _20014;
    wire _20002;
    wire [63:0] _19999;
    wire [63:0] _20000;
    wire [62:0] _20001;
    wire [63:0] _20003;
    wire _20004;
    wire _20005;
    wire _19993;
    wire [63:0] _19990;
    wire [63:0] _19991;
    wire [62:0] _19992;
    wire [63:0] _19994;
    wire _19995;
    wire _19996;
    wire _19984;
    wire [63:0] _19981;
    wire [63:0] _19982;
    wire [62:0] _19983;
    wire [63:0] _19985;
    wire _19986;
    wire _19987;
    wire _19975;
    wire [63:0] _19972;
    wire [63:0] _19973;
    wire [62:0] _19974;
    wire [63:0] _19976;
    wire _19977;
    wire _19978;
    wire _19966;
    wire [63:0] _19963;
    wire [63:0] _19964;
    wire [62:0] _19965;
    wire [63:0] _19967;
    wire _19968;
    wire _19969;
    wire _19957;
    wire [63:0] _19954;
    wire [63:0] _19955;
    wire [62:0] _19956;
    wire [63:0] _19958;
    wire _19959;
    wire _19960;
    wire _19948;
    wire [63:0] _19945;
    wire [63:0] _19946;
    wire [62:0] _19947;
    wire [63:0] _19949;
    wire _19950;
    wire _19951;
    wire _19939;
    wire [63:0] _19936;
    wire [63:0] _19937;
    wire [62:0] _19938;
    wire [63:0] _19940;
    wire _19941;
    wire _19942;
    wire _19930;
    wire [63:0] _19927;
    wire [63:0] _19928;
    wire [62:0] _19929;
    wire [63:0] _19931;
    wire _19932;
    wire _19933;
    wire _19921;
    wire [63:0] _19918;
    wire [63:0] _19919;
    wire [62:0] _19920;
    wire [63:0] _19922;
    wire _19923;
    wire _19924;
    wire _19912;
    wire [63:0] _19909;
    wire [63:0] _19910;
    wire [62:0] _19911;
    wire [63:0] _19913;
    wire _19914;
    wire _19915;
    wire _19903;
    wire [63:0] _19900;
    wire [63:0] _19901;
    wire [62:0] _19902;
    wire [63:0] _19904;
    wire _19905;
    wire _19906;
    wire _19894;
    wire [63:0] _19891;
    wire [63:0] _19892;
    wire [62:0] _19893;
    wire [63:0] _19895;
    wire _19896;
    wire _19897;
    wire _19885;
    wire [63:0] _19882;
    wire [63:0] _19883;
    wire [62:0] _19884;
    wire [63:0] _19886;
    wire _19887;
    wire _19888;
    wire _19876;
    wire [63:0] _19873;
    wire [63:0] _19874;
    wire [62:0] _19875;
    wire [63:0] _19877;
    wire _19878;
    wire _19879;
    wire _19867;
    wire [63:0] _19864;
    wire [63:0] _19865;
    wire [62:0] _19866;
    wire [63:0] _19868;
    wire _19869;
    wire _19870;
    wire [63:0] _19857;
    wire _19858;
    wire [63:0] _19859;
    wire _19860;
    wire _19861;
    wire [63:0] _19862;
    wire [62:0] _19863;
    wire [63:0] _19871;
    wire [62:0] _19872;
    wire [63:0] _19880;
    wire [62:0] _19881;
    wire [63:0] _19889;
    wire [62:0] _19890;
    wire [63:0] _19898;
    wire [62:0] _19899;
    wire [63:0] _19907;
    wire [62:0] _19908;
    wire [63:0] _19916;
    wire [62:0] _19917;
    wire [63:0] _19925;
    wire [62:0] _19926;
    wire [63:0] _19934;
    wire [62:0] _19935;
    wire [63:0] _19943;
    wire [62:0] _19944;
    wire [63:0] _19952;
    wire [62:0] _19953;
    wire [63:0] _19961;
    wire [62:0] _19962;
    wire [63:0] _19970;
    wire [62:0] _19971;
    wire [63:0] _19979;
    wire [62:0] _19980;
    wire [63:0] _19988;
    wire [62:0] _19989;
    wire [63:0] _19997;
    wire [62:0] _19998;
    wire [63:0] _20006;
    wire [62:0] _20007;
    wire [63:0] _20015;
    wire [62:0] _20016;
    wire [63:0] _20024;
    wire [62:0] _20025;
    wire [63:0] _20033;
    wire [62:0] _20034;
    wire [63:0] _20042;
    wire [62:0] _20043;
    wire [63:0] _20051;
    wire [62:0] _20052;
    wire [63:0] _20060;
    wire [62:0] _20061;
    wire [63:0] _20069;
    wire [62:0] _20070;
    wire [63:0] _20078;
    wire [62:0] _20079;
    wire [63:0] _20087;
    wire [62:0] _20088;
    wire [63:0] _20096;
    wire [62:0] _20097;
    wire [63:0] _20105;
    wire [62:0] _20106;
    wire [63:0] _20114;
    wire [62:0] _20115;
    wire [63:0] _20123;
    wire [62:0] _20124;
    wire [63:0] _20132;
    wire [62:0] _20133;
    wire [63:0] _20141;
    wire [62:0] _20142;
    wire [63:0] _20150;
    wire [62:0] _20151;
    wire [63:0] _20159;
    wire [62:0] _20160;
    wire [63:0] _20168;
    wire [62:0] _20169;
    wire [63:0] _20177;
    wire [62:0] _20178;
    wire [63:0] _20186;
    wire [62:0] _20187;
    wire [63:0] _20195;
    wire [62:0] _20196;
    wire [63:0] _20204;
    wire [62:0] _20205;
    wire [63:0] _20213;
    wire [62:0] _20214;
    wire [63:0] _20222;
    wire [62:0] _20223;
    wire [63:0] _20231;
    wire [62:0] _20232;
    wire [63:0] _20240;
    wire [62:0] _20241;
    wire [63:0] _20249;
    wire [62:0] _20250;
    wire [63:0] _20258;
    wire [62:0] _20259;
    wire [63:0] _20267;
    wire [62:0] _20268;
    wire [63:0] _20276;
    wire [62:0] _20277;
    wire [63:0] _20285;
    wire [62:0] _20286;
    wire [63:0] _20294;
    wire [62:0] _20295;
    wire [63:0] _20303;
    wire [62:0] _20304;
    wire [63:0] _20312;
    wire [62:0] _20313;
    wire [63:0] _20321;
    wire [62:0] _20322;
    wire [63:0] _20330;
    wire [62:0] _20331;
    wire [63:0] _20339;
    wire [62:0] _20340;
    wire [63:0] _20348;
    wire [62:0] _20349;
    wire [63:0] _20357;
    wire [62:0] _20358;
    wire [63:0] _20366;
    wire [62:0] _20367;
    wire [63:0] _20375;
    wire [62:0] _20376;
    wire [63:0] _20384;
    wire [62:0] _20385;
    wire [63:0] _20393;
    wire [62:0] _20394;
    wire [63:0] _20402;
    wire [62:0] _20403;
    wire [63:0] _20411;
    wire [62:0] _20412;
    wire [63:0] _20420;
    wire [62:0] _20421;
    wire [63:0] _20429;
    wire [63:0] _20431;
    wire [127:0] _20432;
    wire [63:0] _20433;
    wire [63:0] _21015;
    wire _19843;
    wire [63:0] _19840;
    wire [63:0] _19841;
    wire [62:0] _19842;
    wire [63:0] _19844;
    wire _19845;
    wire _19846;
    wire _19834;
    wire [63:0] _19831;
    wire [63:0] _19832;
    wire [62:0] _19833;
    wire [63:0] _19835;
    wire _19836;
    wire _19837;
    wire _19825;
    wire [63:0] _19822;
    wire [63:0] _19823;
    wire [62:0] _19824;
    wire [63:0] _19826;
    wire _19827;
    wire _19828;
    wire _19816;
    wire [63:0] _19813;
    wire [63:0] _19814;
    wire [62:0] _19815;
    wire [63:0] _19817;
    wire _19818;
    wire _19819;
    wire _19807;
    wire [63:0] _19804;
    wire [63:0] _19805;
    wire [62:0] _19806;
    wire [63:0] _19808;
    wire _19809;
    wire _19810;
    wire _19798;
    wire [63:0] _19795;
    wire [63:0] _19796;
    wire [62:0] _19797;
    wire [63:0] _19799;
    wire _19800;
    wire _19801;
    wire _19789;
    wire [63:0] _19786;
    wire [63:0] _19787;
    wire [62:0] _19788;
    wire [63:0] _19790;
    wire _19791;
    wire _19792;
    wire _19780;
    wire [63:0] _19777;
    wire [63:0] _19778;
    wire [62:0] _19779;
    wire [63:0] _19781;
    wire _19782;
    wire _19783;
    wire _19771;
    wire [63:0] _19768;
    wire [63:0] _19769;
    wire [62:0] _19770;
    wire [63:0] _19772;
    wire _19773;
    wire _19774;
    wire _19762;
    wire [63:0] _19759;
    wire [63:0] _19760;
    wire [62:0] _19761;
    wire [63:0] _19763;
    wire _19764;
    wire _19765;
    wire _19753;
    wire [63:0] _19750;
    wire [63:0] _19751;
    wire [62:0] _19752;
    wire [63:0] _19754;
    wire _19755;
    wire _19756;
    wire _19744;
    wire [63:0] _19741;
    wire [63:0] _19742;
    wire [62:0] _19743;
    wire [63:0] _19745;
    wire _19746;
    wire _19747;
    wire _19735;
    wire [63:0] _19732;
    wire [63:0] _19733;
    wire [62:0] _19734;
    wire [63:0] _19736;
    wire _19737;
    wire _19738;
    wire _19726;
    wire [63:0] _19723;
    wire [63:0] _19724;
    wire [62:0] _19725;
    wire [63:0] _19727;
    wire _19728;
    wire _19729;
    wire _19717;
    wire [63:0] _19714;
    wire [63:0] _19715;
    wire [62:0] _19716;
    wire [63:0] _19718;
    wire _19719;
    wire _19720;
    wire _19708;
    wire [63:0] _19705;
    wire [63:0] _19706;
    wire [62:0] _19707;
    wire [63:0] _19709;
    wire _19710;
    wire _19711;
    wire _19699;
    wire [63:0] _19696;
    wire [63:0] _19697;
    wire [62:0] _19698;
    wire [63:0] _19700;
    wire _19701;
    wire _19702;
    wire _19690;
    wire [63:0] _19687;
    wire [63:0] _19688;
    wire [62:0] _19689;
    wire [63:0] _19691;
    wire _19692;
    wire _19693;
    wire _19681;
    wire [63:0] _19678;
    wire [63:0] _19679;
    wire [62:0] _19680;
    wire [63:0] _19682;
    wire _19683;
    wire _19684;
    wire _19672;
    wire [63:0] _19669;
    wire [63:0] _19670;
    wire [62:0] _19671;
    wire [63:0] _19673;
    wire _19674;
    wire _19675;
    wire _19663;
    wire [63:0] _19660;
    wire [63:0] _19661;
    wire [62:0] _19662;
    wire [63:0] _19664;
    wire _19665;
    wire _19666;
    wire _19654;
    wire [63:0] _19651;
    wire [63:0] _19652;
    wire [62:0] _19653;
    wire [63:0] _19655;
    wire _19656;
    wire _19657;
    wire _19645;
    wire [63:0] _19642;
    wire [63:0] _19643;
    wire [62:0] _19644;
    wire [63:0] _19646;
    wire _19647;
    wire _19648;
    wire _19636;
    wire [63:0] _19633;
    wire [63:0] _19634;
    wire [62:0] _19635;
    wire [63:0] _19637;
    wire _19638;
    wire _19639;
    wire _19627;
    wire [63:0] _19624;
    wire [63:0] _19625;
    wire [62:0] _19626;
    wire [63:0] _19628;
    wire _19629;
    wire _19630;
    wire _19618;
    wire [63:0] _19615;
    wire [63:0] _19616;
    wire [62:0] _19617;
    wire [63:0] _19619;
    wire _19620;
    wire _19621;
    wire _19609;
    wire [63:0] _19606;
    wire [63:0] _19607;
    wire [62:0] _19608;
    wire [63:0] _19610;
    wire _19611;
    wire _19612;
    wire _19600;
    wire [63:0] _19597;
    wire [63:0] _19598;
    wire [62:0] _19599;
    wire [63:0] _19601;
    wire _19602;
    wire _19603;
    wire _19591;
    wire [63:0] _19588;
    wire [63:0] _19589;
    wire [62:0] _19590;
    wire [63:0] _19592;
    wire _19593;
    wire _19594;
    wire _19582;
    wire [63:0] _19579;
    wire [63:0] _19580;
    wire [62:0] _19581;
    wire [63:0] _19583;
    wire _19584;
    wire _19585;
    wire _19573;
    wire [63:0] _19570;
    wire [63:0] _19571;
    wire [62:0] _19572;
    wire [63:0] _19574;
    wire _19575;
    wire _19576;
    wire _19564;
    wire [63:0] _19561;
    wire [63:0] _19562;
    wire [62:0] _19563;
    wire [63:0] _19565;
    wire _19566;
    wire _19567;
    wire _19555;
    wire [63:0] _19552;
    wire [63:0] _19553;
    wire [62:0] _19554;
    wire [63:0] _19556;
    wire _19557;
    wire _19558;
    wire _19546;
    wire [63:0] _19543;
    wire [63:0] _19544;
    wire [62:0] _19545;
    wire [63:0] _19547;
    wire _19548;
    wire _19549;
    wire _19537;
    wire [63:0] _19534;
    wire [63:0] _19535;
    wire [62:0] _19536;
    wire [63:0] _19538;
    wire _19539;
    wire _19540;
    wire _19528;
    wire [63:0] _19525;
    wire [63:0] _19526;
    wire [62:0] _19527;
    wire [63:0] _19529;
    wire _19530;
    wire _19531;
    wire _19519;
    wire [63:0] _19516;
    wire [63:0] _19517;
    wire [62:0] _19518;
    wire [63:0] _19520;
    wire _19521;
    wire _19522;
    wire _19510;
    wire [63:0] _19507;
    wire [63:0] _19508;
    wire [62:0] _19509;
    wire [63:0] _19511;
    wire _19512;
    wire _19513;
    wire _19501;
    wire [63:0] _19498;
    wire [63:0] _19499;
    wire [62:0] _19500;
    wire [63:0] _19502;
    wire _19503;
    wire _19504;
    wire _19492;
    wire [63:0] _19489;
    wire [63:0] _19490;
    wire [62:0] _19491;
    wire [63:0] _19493;
    wire _19494;
    wire _19495;
    wire _19483;
    wire [63:0] _19480;
    wire [63:0] _19481;
    wire [62:0] _19482;
    wire [63:0] _19484;
    wire _19485;
    wire _19486;
    wire _19474;
    wire [63:0] _19471;
    wire [63:0] _19472;
    wire [62:0] _19473;
    wire [63:0] _19475;
    wire _19476;
    wire _19477;
    wire _19465;
    wire [63:0] _19462;
    wire [63:0] _19463;
    wire [62:0] _19464;
    wire [63:0] _19466;
    wire _19467;
    wire _19468;
    wire _19456;
    wire [63:0] _19453;
    wire [63:0] _19454;
    wire [62:0] _19455;
    wire [63:0] _19457;
    wire _19458;
    wire _19459;
    wire _19447;
    wire [63:0] _19444;
    wire [63:0] _19445;
    wire [62:0] _19446;
    wire [63:0] _19448;
    wire _19449;
    wire _19450;
    wire _19438;
    wire [63:0] _19435;
    wire [63:0] _19436;
    wire [62:0] _19437;
    wire [63:0] _19439;
    wire _19440;
    wire _19441;
    wire _19429;
    wire [63:0] _19426;
    wire [63:0] _19427;
    wire [62:0] _19428;
    wire [63:0] _19430;
    wire _19431;
    wire _19432;
    wire _19420;
    wire [63:0] _19417;
    wire [63:0] _19418;
    wire [62:0] _19419;
    wire [63:0] _19421;
    wire _19422;
    wire _19423;
    wire _19411;
    wire [63:0] _19408;
    wire [63:0] _19409;
    wire [62:0] _19410;
    wire [63:0] _19412;
    wire _19413;
    wire _19414;
    wire _19402;
    wire [63:0] _19399;
    wire [63:0] _19400;
    wire [62:0] _19401;
    wire [63:0] _19403;
    wire _19404;
    wire _19405;
    wire _19393;
    wire [63:0] _19390;
    wire [63:0] _19391;
    wire [62:0] _19392;
    wire [63:0] _19394;
    wire _19395;
    wire _19396;
    wire _19384;
    wire [63:0] _19381;
    wire [63:0] _19382;
    wire [62:0] _19383;
    wire [63:0] _19385;
    wire _19386;
    wire _19387;
    wire _19375;
    wire [63:0] _19372;
    wire [63:0] _19373;
    wire [62:0] _19374;
    wire [63:0] _19376;
    wire _19377;
    wire _19378;
    wire _19366;
    wire [63:0] _19363;
    wire [63:0] _19364;
    wire [62:0] _19365;
    wire [63:0] _19367;
    wire _19368;
    wire _19369;
    wire _19357;
    wire [63:0] _19354;
    wire [63:0] _19355;
    wire [62:0] _19356;
    wire [63:0] _19358;
    wire _19359;
    wire _19360;
    wire _19348;
    wire [63:0] _19345;
    wire [63:0] _19346;
    wire [62:0] _19347;
    wire [63:0] _19349;
    wire _19350;
    wire _19351;
    wire _19339;
    wire [63:0] _19336;
    wire [63:0] _19337;
    wire [62:0] _19338;
    wire [63:0] _19340;
    wire _19341;
    wire _19342;
    wire _19330;
    wire [63:0] _19327;
    wire [63:0] _19328;
    wire [62:0] _19329;
    wire [63:0] _19331;
    wire _19332;
    wire _19333;
    wire _19321;
    wire [63:0] _19318;
    wire [63:0] _19319;
    wire [62:0] _19320;
    wire [63:0] _19322;
    wire _19323;
    wire _19324;
    wire _19312;
    wire [63:0] _19309;
    wire [63:0] _19310;
    wire [62:0] _19311;
    wire [63:0] _19313;
    wire _19314;
    wire _19315;
    wire _19303;
    wire [63:0] _19300;
    wire [63:0] _19301;
    wire [62:0] _19302;
    wire [63:0] _19304;
    wire _19305;
    wire _19306;
    wire _19294;
    wire [63:0] _19291;
    wire [63:0] _19292;
    wire [62:0] _19293;
    wire [63:0] _19295;
    wire _19296;
    wire _19297;
    wire _19285;
    wire [63:0] _19282;
    wire [63:0] _19283;
    wire [62:0] _19284;
    wire [63:0] _19286;
    wire _19287;
    wire _19288;
    wire [63:0] _19277;
    wire [63:0] _19273;
    wire [63:0] _19274;
    wire _19275;
    wire [63:0] _19276;
    wire _19278;
    wire _19279;
    wire [63:0] _19280;
    wire [62:0] _19281;
    wire [63:0] _19289;
    wire [62:0] _19290;
    wire [63:0] _19298;
    wire [62:0] _19299;
    wire [63:0] _19307;
    wire [62:0] _19308;
    wire [63:0] _19316;
    wire [62:0] _19317;
    wire [63:0] _19325;
    wire [62:0] _19326;
    wire [63:0] _19334;
    wire [62:0] _19335;
    wire [63:0] _19343;
    wire [62:0] _19344;
    wire [63:0] _19352;
    wire [62:0] _19353;
    wire [63:0] _19361;
    wire [62:0] _19362;
    wire [63:0] _19370;
    wire [62:0] _19371;
    wire [63:0] _19379;
    wire [62:0] _19380;
    wire [63:0] _19388;
    wire [62:0] _19389;
    wire [63:0] _19397;
    wire [62:0] _19398;
    wire [63:0] _19406;
    wire [62:0] _19407;
    wire [63:0] _19415;
    wire [62:0] _19416;
    wire [63:0] _19424;
    wire [62:0] _19425;
    wire [63:0] _19433;
    wire [62:0] _19434;
    wire [63:0] _19442;
    wire [62:0] _19443;
    wire [63:0] _19451;
    wire [62:0] _19452;
    wire [63:0] _19460;
    wire [62:0] _19461;
    wire [63:0] _19469;
    wire [62:0] _19470;
    wire [63:0] _19478;
    wire [62:0] _19479;
    wire [63:0] _19487;
    wire [62:0] _19488;
    wire [63:0] _19496;
    wire [62:0] _19497;
    wire [63:0] _19505;
    wire [62:0] _19506;
    wire [63:0] _19514;
    wire [62:0] _19515;
    wire [63:0] _19523;
    wire [62:0] _19524;
    wire [63:0] _19532;
    wire [62:0] _19533;
    wire [63:0] _19541;
    wire [62:0] _19542;
    wire [63:0] _19550;
    wire [62:0] _19551;
    wire [63:0] _19559;
    wire [62:0] _19560;
    wire [63:0] _19568;
    wire [62:0] _19569;
    wire [63:0] _19577;
    wire [62:0] _19578;
    wire [63:0] _19586;
    wire [62:0] _19587;
    wire [63:0] _19595;
    wire [62:0] _19596;
    wire [63:0] _19604;
    wire [62:0] _19605;
    wire [63:0] _19613;
    wire [62:0] _19614;
    wire [63:0] _19622;
    wire [62:0] _19623;
    wire [63:0] _19631;
    wire [62:0] _19632;
    wire [63:0] _19640;
    wire [62:0] _19641;
    wire [63:0] _19649;
    wire [62:0] _19650;
    wire [63:0] _19658;
    wire [62:0] _19659;
    wire [63:0] _19667;
    wire [62:0] _19668;
    wire [63:0] _19676;
    wire [62:0] _19677;
    wire [63:0] _19685;
    wire [62:0] _19686;
    wire [63:0] _19694;
    wire [62:0] _19695;
    wire [63:0] _19703;
    wire [62:0] _19704;
    wire [63:0] _19712;
    wire [62:0] _19713;
    wire [63:0] _19721;
    wire [62:0] _19722;
    wire [63:0] _19730;
    wire [62:0] _19731;
    wire [63:0] _19739;
    wire [62:0] _19740;
    wire [63:0] _19748;
    wire [62:0] _19749;
    wire [63:0] _19757;
    wire [62:0] _19758;
    wire [63:0] _19766;
    wire [62:0] _19767;
    wire [63:0] _19775;
    wire [62:0] _19776;
    wire [63:0] _19784;
    wire [62:0] _19785;
    wire [63:0] _19793;
    wire [62:0] _19794;
    wire [63:0] _19802;
    wire [62:0] _19803;
    wire [63:0] _19811;
    wire [62:0] _19812;
    wire [63:0] _19820;
    wire [62:0] _19821;
    wire [63:0] _19829;
    wire [62:0] _19830;
    wire [63:0] _19838;
    wire [62:0] _19839;
    wire [63:0] _19847;
    wire [127:0] _19848;
    wire [63:0] _19849;
    wire _19850;
    wire [63:0] _19851;
    wire [63:0] _19267;
    wire _19268;
    wire [63:0] _19269;
    wire _19852;
    wire _19853;
    wire [63:0] _21016;
    wire [63:0] _22767;
    wire _19256;
    wire [63:0] _19253;
    wire [63:0] _19254;
    wire [62:0] _19255;
    wire [63:0] _19257;
    wire _19258;
    wire _19259;
    wire _19247;
    wire [63:0] _19244;
    wire [63:0] _19245;
    wire [62:0] _19246;
    wire [63:0] _19248;
    wire _19249;
    wire _19250;
    wire _19238;
    wire [63:0] _19235;
    wire [63:0] _19236;
    wire [62:0] _19237;
    wire [63:0] _19239;
    wire _19240;
    wire _19241;
    wire _19229;
    wire [63:0] _19226;
    wire [63:0] _19227;
    wire [62:0] _19228;
    wire [63:0] _19230;
    wire _19231;
    wire _19232;
    wire _19220;
    wire [63:0] _19217;
    wire [63:0] _19218;
    wire [62:0] _19219;
    wire [63:0] _19221;
    wire _19222;
    wire _19223;
    wire _19211;
    wire [63:0] _19208;
    wire [63:0] _19209;
    wire [62:0] _19210;
    wire [63:0] _19212;
    wire _19213;
    wire _19214;
    wire _19202;
    wire [63:0] _19199;
    wire [63:0] _19200;
    wire [62:0] _19201;
    wire [63:0] _19203;
    wire _19204;
    wire _19205;
    wire _19193;
    wire [63:0] _19190;
    wire [63:0] _19191;
    wire [62:0] _19192;
    wire [63:0] _19194;
    wire _19195;
    wire _19196;
    wire _19184;
    wire [63:0] _19181;
    wire [63:0] _19182;
    wire [62:0] _19183;
    wire [63:0] _19185;
    wire _19186;
    wire _19187;
    wire _19175;
    wire [63:0] _19172;
    wire [63:0] _19173;
    wire [62:0] _19174;
    wire [63:0] _19176;
    wire _19177;
    wire _19178;
    wire _19166;
    wire [63:0] _19163;
    wire [63:0] _19164;
    wire [62:0] _19165;
    wire [63:0] _19167;
    wire _19168;
    wire _19169;
    wire _19157;
    wire [63:0] _19154;
    wire [63:0] _19155;
    wire [62:0] _19156;
    wire [63:0] _19158;
    wire _19159;
    wire _19160;
    wire _19148;
    wire [63:0] _19145;
    wire [63:0] _19146;
    wire [62:0] _19147;
    wire [63:0] _19149;
    wire _19150;
    wire _19151;
    wire _19139;
    wire [63:0] _19136;
    wire [63:0] _19137;
    wire [62:0] _19138;
    wire [63:0] _19140;
    wire _19141;
    wire _19142;
    wire _19130;
    wire [63:0] _19127;
    wire [63:0] _19128;
    wire [62:0] _19129;
    wire [63:0] _19131;
    wire _19132;
    wire _19133;
    wire _19121;
    wire [63:0] _19118;
    wire [63:0] _19119;
    wire [62:0] _19120;
    wire [63:0] _19122;
    wire _19123;
    wire _19124;
    wire _19112;
    wire [63:0] _19109;
    wire [63:0] _19110;
    wire [62:0] _19111;
    wire [63:0] _19113;
    wire _19114;
    wire _19115;
    wire _19103;
    wire [63:0] _19100;
    wire [63:0] _19101;
    wire [62:0] _19102;
    wire [63:0] _19104;
    wire _19105;
    wire _19106;
    wire _19094;
    wire [63:0] _19091;
    wire [63:0] _19092;
    wire [62:0] _19093;
    wire [63:0] _19095;
    wire _19096;
    wire _19097;
    wire _19085;
    wire [63:0] _19082;
    wire [63:0] _19083;
    wire [62:0] _19084;
    wire [63:0] _19086;
    wire _19087;
    wire _19088;
    wire _19076;
    wire [63:0] _19073;
    wire [63:0] _19074;
    wire [62:0] _19075;
    wire [63:0] _19077;
    wire _19078;
    wire _19079;
    wire _19067;
    wire [63:0] _19064;
    wire [63:0] _19065;
    wire [62:0] _19066;
    wire [63:0] _19068;
    wire _19069;
    wire _19070;
    wire _19058;
    wire [63:0] _19055;
    wire [63:0] _19056;
    wire [62:0] _19057;
    wire [63:0] _19059;
    wire _19060;
    wire _19061;
    wire _19049;
    wire [63:0] _19046;
    wire [63:0] _19047;
    wire [62:0] _19048;
    wire [63:0] _19050;
    wire _19051;
    wire _19052;
    wire _19040;
    wire [63:0] _19037;
    wire [63:0] _19038;
    wire [62:0] _19039;
    wire [63:0] _19041;
    wire _19042;
    wire _19043;
    wire _19031;
    wire [63:0] _19028;
    wire [63:0] _19029;
    wire [62:0] _19030;
    wire [63:0] _19032;
    wire _19033;
    wire _19034;
    wire _19022;
    wire [63:0] _19019;
    wire [63:0] _19020;
    wire [62:0] _19021;
    wire [63:0] _19023;
    wire _19024;
    wire _19025;
    wire _19013;
    wire [63:0] _19010;
    wire [63:0] _19011;
    wire [62:0] _19012;
    wire [63:0] _19014;
    wire _19015;
    wire _19016;
    wire _19004;
    wire [63:0] _19001;
    wire [63:0] _19002;
    wire [62:0] _19003;
    wire [63:0] _19005;
    wire _19006;
    wire _19007;
    wire _18995;
    wire [63:0] _18992;
    wire [63:0] _18993;
    wire [62:0] _18994;
    wire [63:0] _18996;
    wire _18997;
    wire _18998;
    wire _18986;
    wire [63:0] _18983;
    wire [63:0] _18984;
    wire [62:0] _18985;
    wire [63:0] _18987;
    wire _18988;
    wire _18989;
    wire _18977;
    wire [63:0] _18974;
    wire [63:0] _18975;
    wire [62:0] _18976;
    wire [63:0] _18978;
    wire _18979;
    wire _18980;
    wire _18968;
    wire [63:0] _18965;
    wire [63:0] _18966;
    wire [62:0] _18967;
    wire [63:0] _18969;
    wire _18970;
    wire _18971;
    wire _18959;
    wire [63:0] _18956;
    wire [63:0] _18957;
    wire [62:0] _18958;
    wire [63:0] _18960;
    wire _18961;
    wire _18962;
    wire _18950;
    wire [63:0] _18947;
    wire [63:0] _18948;
    wire [62:0] _18949;
    wire [63:0] _18951;
    wire _18952;
    wire _18953;
    wire _18941;
    wire [63:0] _18938;
    wire [63:0] _18939;
    wire [62:0] _18940;
    wire [63:0] _18942;
    wire _18943;
    wire _18944;
    wire _18932;
    wire [63:0] _18929;
    wire [63:0] _18930;
    wire [62:0] _18931;
    wire [63:0] _18933;
    wire _18934;
    wire _18935;
    wire _18923;
    wire [63:0] _18920;
    wire [63:0] _18921;
    wire [62:0] _18922;
    wire [63:0] _18924;
    wire _18925;
    wire _18926;
    wire _18914;
    wire [63:0] _18911;
    wire [63:0] _18912;
    wire [62:0] _18913;
    wire [63:0] _18915;
    wire _18916;
    wire _18917;
    wire _18905;
    wire [63:0] _18902;
    wire [63:0] _18903;
    wire [62:0] _18904;
    wire [63:0] _18906;
    wire _18907;
    wire _18908;
    wire _18896;
    wire [63:0] _18893;
    wire [63:0] _18894;
    wire [62:0] _18895;
    wire [63:0] _18897;
    wire _18898;
    wire _18899;
    wire _18887;
    wire [63:0] _18884;
    wire [63:0] _18885;
    wire [62:0] _18886;
    wire [63:0] _18888;
    wire _18889;
    wire _18890;
    wire _18878;
    wire [63:0] _18875;
    wire [63:0] _18876;
    wire [62:0] _18877;
    wire [63:0] _18879;
    wire _18880;
    wire _18881;
    wire _18869;
    wire [63:0] _18866;
    wire [63:0] _18867;
    wire [62:0] _18868;
    wire [63:0] _18870;
    wire _18871;
    wire _18872;
    wire _18860;
    wire [63:0] _18857;
    wire [63:0] _18858;
    wire [62:0] _18859;
    wire [63:0] _18861;
    wire _18862;
    wire _18863;
    wire _18851;
    wire [63:0] _18848;
    wire [63:0] _18849;
    wire [62:0] _18850;
    wire [63:0] _18852;
    wire _18853;
    wire _18854;
    wire _18842;
    wire [63:0] _18839;
    wire [63:0] _18840;
    wire [62:0] _18841;
    wire [63:0] _18843;
    wire _18844;
    wire _18845;
    wire _18833;
    wire [63:0] _18830;
    wire [63:0] _18831;
    wire [62:0] _18832;
    wire [63:0] _18834;
    wire _18835;
    wire _18836;
    wire _18824;
    wire [63:0] _18821;
    wire [63:0] _18822;
    wire [62:0] _18823;
    wire [63:0] _18825;
    wire _18826;
    wire _18827;
    wire _18815;
    wire [63:0] _18812;
    wire [63:0] _18813;
    wire [62:0] _18814;
    wire [63:0] _18816;
    wire _18817;
    wire _18818;
    wire _18806;
    wire [63:0] _18803;
    wire [63:0] _18804;
    wire [62:0] _18805;
    wire [63:0] _18807;
    wire _18808;
    wire _18809;
    wire _18797;
    wire [63:0] _18794;
    wire [63:0] _18795;
    wire [62:0] _18796;
    wire [63:0] _18798;
    wire _18799;
    wire _18800;
    wire _18788;
    wire [63:0] _18785;
    wire [63:0] _18786;
    wire [62:0] _18787;
    wire [63:0] _18789;
    wire _18790;
    wire _18791;
    wire _18779;
    wire [63:0] _18776;
    wire [63:0] _18777;
    wire [62:0] _18778;
    wire [63:0] _18780;
    wire _18781;
    wire _18782;
    wire _18770;
    wire [63:0] _18767;
    wire [63:0] _18768;
    wire [62:0] _18769;
    wire [63:0] _18771;
    wire _18772;
    wire _18773;
    wire _18761;
    wire [63:0] _18758;
    wire [63:0] _18759;
    wire [62:0] _18760;
    wire [63:0] _18762;
    wire _18763;
    wire _18764;
    wire _18752;
    wire [63:0] _18749;
    wire [63:0] _18750;
    wire [62:0] _18751;
    wire [63:0] _18753;
    wire _18754;
    wire _18755;
    wire _18743;
    wire [63:0] _18740;
    wire [63:0] _18741;
    wire [62:0] _18742;
    wire [63:0] _18744;
    wire _18745;
    wire _18746;
    wire _18734;
    wire [63:0] _18731;
    wire [63:0] _18732;
    wire [62:0] _18733;
    wire [63:0] _18735;
    wire _18736;
    wire _18737;
    wire _18725;
    wire [63:0] _18722;
    wire [63:0] _18723;
    wire [62:0] _18724;
    wire [63:0] _18726;
    wire _18727;
    wire _18728;
    wire _18716;
    wire [63:0] _18713;
    wire [63:0] _18714;
    wire [62:0] _18715;
    wire [63:0] _18717;
    wire _18718;
    wire _18719;
    wire _18707;
    wire [63:0] _18704;
    wire [63:0] _18705;
    wire [62:0] _18706;
    wire [63:0] _18708;
    wire _18709;
    wire _18710;
    wire _18698;
    wire [63:0] _18695;
    wire [63:0] _18696;
    wire [62:0] _18697;
    wire [63:0] _18699;
    wire _18700;
    wire _18701;
    wire [63:0] _18685;
    wire [127:0] _18686;
    wire [63:0] _18687;
    wire _18688;
    wire [63:0] _18689;
    wire _18691;
    wire _18692;
    wire [63:0] _18693;
    wire [62:0] _18694;
    wire [63:0] _18702;
    wire [62:0] _18703;
    wire [63:0] _18711;
    wire [62:0] _18712;
    wire [63:0] _18720;
    wire [62:0] _18721;
    wire [63:0] _18729;
    wire [62:0] _18730;
    wire [63:0] _18738;
    wire [62:0] _18739;
    wire [63:0] _18747;
    wire [62:0] _18748;
    wire [63:0] _18756;
    wire [62:0] _18757;
    wire [63:0] _18765;
    wire [62:0] _18766;
    wire [63:0] _18774;
    wire [62:0] _18775;
    wire [63:0] _18783;
    wire [62:0] _18784;
    wire [63:0] _18792;
    wire [62:0] _18793;
    wire [63:0] _18801;
    wire [62:0] _18802;
    wire [63:0] _18810;
    wire [62:0] _18811;
    wire [63:0] _18819;
    wire [62:0] _18820;
    wire [63:0] _18828;
    wire [62:0] _18829;
    wire [63:0] _18837;
    wire [62:0] _18838;
    wire [63:0] _18846;
    wire [62:0] _18847;
    wire [63:0] _18855;
    wire [62:0] _18856;
    wire [63:0] _18864;
    wire [62:0] _18865;
    wire [63:0] _18873;
    wire [62:0] _18874;
    wire [63:0] _18882;
    wire [62:0] _18883;
    wire [63:0] _18891;
    wire [62:0] _18892;
    wire [63:0] _18900;
    wire [62:0] _18901;
    wire [63:0] _18909;
    wire [62:0] _18910;
    wire [63:0] _18918;
    wire [62:0] _18919;
    wire [63:0] _18927;
    wire [62:0] _18928;
    wire [63:0] _18936;
    wire [62:0] _18937;
    wire [63:0] _18945;
    wire [62:0] _18946;
    wire [63:0] _18954;
    wire [62:0] _18955;
    wire [63:0] _18963;
    wire [62:0] _18964;
    wire [63:0] _18972;
    wire [62:0] _18973;
    wire [63:0] _18981;
    wire [62:0] _18982;
    wire [63:0] _18990;
    wire [62:0] _18991;
    wire [63:0] _18999;
    wire [62:0] _19000;
    wire [63:0] _19008;
    wire [62:0] _19009;
    wire [63:0] _19017;
    wire [62:0] _19018;
    wire [63:0] _19026;
    wire [62:0] _19027;
    wire [63:0] _19035;
    wire [62:0] _19036;
    wire [63:0] _19044;
    wire [62:0] _19045;
    wire [63:0] _19053;
    wire [62:0] _19054;
    wire [63:0] _19062;
    wire [62:0] _19063;
    wire [63:0] _19071;
    wire [62:0] _19072;
    wire [63:0] _19080;
    wire [62:0] _19081;
    wire [63:0] _19089;
    wire [62:0] _19090;
    wire [63:0] _19098;
    wire [62:0] _19099;
    wire [63:0] _19107;
    wire [62:0] _19108;
    wire [63:0] _19116;
    wire [62:0] _19117;
    wire [63:0] _19125;
    wire [62:0] _19126;
    wire [63:0] _19134;
    wire [62:0] _19135;
    wire [63:0] _19143;
    wire [62:0] _19144;
    wire [63:0] _19152;
    wire [62:0] _19153;
    wire [63:0] _19161;
    wire [62:0] _19162;
    wire [63:0] _19170;
    wire [62:0] _19171;
    wire [63:0] _19179;
    wire [62:0] _19180;
    wire [63:0] _19188;
    wire [62:0] _19189;
    wire [63:0] _19197;
    wire [62:0] _19198;
    wire [63:0] _19206;
    wire [62:0] _19207;
    wire [63:0] _19215;
    wire [62:0] _19216;
    wire [63:0] _19224;
    wire [62:0] _19225;
    wire [63:0] _19233;
    wire [62:0] _19234;
    wire [63:0] _19242;
    wire [62:0] _19243;
    wire [63:0] _19251;
    wire [62:0] _19252;
    wire [63:0] _19260;
    wire [127:0] _19261;
    wire [63:0] _19262;
    wire _18673;
    wire [63:0] _18670;
    wire [63:0] _18671;
    wire [62:0] _18672;
    wire [63:0] _18674;
    wire _18675;
    wire _18676;
    wire _18664;
    wire [63:0] _18661;
    wire [63:0] _18662;
    wire [62:0] _18663;
    wire [63:0] _18665;
    wire _18666;
    wire _18667;
    wire _18655;
    wire [63:0] _18652;
    wire [63:0] _18653;
    wire [62:0] _18654;
    wire [63:0] _18656;
    wire _18657;
    wire _18658;
    wire _18646;
    wire [63:0] _18643;
    wire [63:0] _18644;
    wire [62:0] _18645;
    wire [63:0] _18647;
    wire _18648;
    wire _18649;
    wire _18637;
    wire [63:0] _18634;
    wire [63:0] _18635;
    wire [62:0] _18636;
    wire [63:0] _18638;
    wire _18639;
    wire _18640;
    wire _18628;
    wire [63:0] _18625;
    wire [63:0] _18626;
    wire [62:0] _18627;
    wire [63:0] _18629;
    wire _18630;
    wire _18631;
    wire _18619;
    wire [63:0] _18616;
    wire [63:0] _18617;
    wire [62:0] _18618;
    wire [63:0] _18620;
    wire _18621;
    wire _18622;
    wire _18610;
    wire [63:0] _18607;
    wire [63:0] _18608;
    wire [62:0] _18609;
    wire [63:0] _18611;
    wire _18612;
    wire _18613;
    wire _18601;
    wire [63:0] _18598;
    wire [63:0] _18599;
    wire [62:0] _18600;
    wire [63:0] _18602;
    wire _18603;
    wire _18604;
    wire _18592;
    wire [63:0] _18589;
    wire [63:0] _18590;
    wire [62:0] _18591;
    wire [63:0] _18593;
    wire _18594;
    wire _18595;
    wire _18583;
    wire [63:0] _18580;
    wire [63:0] _18581;
    wire [62:0] _18582;
    wire [63:0] _18584;
    wire _18585;
    wire _18586;
    wire _18574;
    wire [63:0] _18571;
    wire [63:0] _18572;
    wire [62:0] _18573;
    wire [63:0] _18575;
    wire _18576;
    wire _18577;
    wire _18565;
    wire [63:0] _18562;
    wire [63:0] _18563;
    wire [62:0] _18564;
    wire [63:0] _18566;
    wire _18567;
    wire _18568;
    wire _18556;
    wire [63:0] _18553;
    wire [63:0] _18554;
    wire [62:0] _18555;
    wire [63:0] _18557;
    wire _18558;
    wire _18559;
    wire _18547;
    wire [63:0] _18544;
    wire [63:0] _18545;
    wire [62:0] _18546;
    wire [63:0] _18548;
    wire _18549;
    wire _18550;
    wire _18538;
    wire [63:0] _18535;
    wire [63:0] _18536;
    wire [62:0] _18537;
    wire [63:0] _18539;
    wire _18540;
    wire _18541;
    wire _18529;
    wire [63:0] _18526;
    wire [63:0] _18527;
    wire [62:0] _18528;
    wire [63:0] _18530;
    wire _18531;
    wire _18532;
    wire _18520;
    wire [63:0] _18517;
    wire [63:0] _18518;
    wire [62:0] _18519;
    wire [63:0] _18521;
    wire _18522;
    wire _18523;
    wire _18511;
    wire [63:0] _18508;
    wire [63:0] _18509;
    wire [62:0] _18510;
    wire [63:0] _18512;
    wire _18513;
    wire _18514;
    wire _18502;
    wire [63:0] _18499;
    wire [63:0] _18500;
    wire [62:0] _18501;
    wire [63:0] _18503;
    wire _18504;
    wire _18505;
    wire _18493;
    wire [63:0] _18490;
    wire [63:0] _18491;
    wire [62:0] _18492;
    wire [63:0] _18494;
    wire _18495;
    wire _18496;
    wire _18484;
    wire [63:0] _18481;
    wire [63:0] _18482;
    wire [62:0] _18483;
    wire [63:0] _18485;
    wire _18486;
    wire _18487;
    wire _18475;
    wire [63:0] _18472;
    wire [63:0] _18473;
    wire [62:0] _18474;
    wire [63:0] _18476;
    wire _18477;
    wire _18478;
    wire _18466;
    wire [63:0] _18463;
    wire [63:0] _18464;
    wire [62:0] _18465;
    wire [63:0] _18467;
    wire _18468;
    wire _18469;
    wire _18457;
    wire [63:0] _18454;
    wire [63:0] _18455;
    wire [62:0] _18456;
    wire [63:0] _18458;
    wire _18459;
    wire _18460;
    wire _18448;
    wire [63:0] _18445;
    wire [63:0] _18446;
    wire [62:0] _18447;
    wire [63:0] _18449;
    wire _18450;
    wire _18451;
    wire _18439;
    wire [63:0] _18436;
    wire [63:0] _18437;
    wire [62:0] _18438;
    wire [63:0] _18440;
    wire _18441;
    wire _18442;
    wire _18430;
    wire [63:0] _18427;
    wire [63:0] _18428;
    wire [62:0] _18429;
    wire [63:0] _18431;
    wire _18432;
    wire _18433;
    wire _18421;
    wire [63:0] _18418;
    wire [63:0] _18419;
    wire [62:0] _18420;
    wire [63:0] _18422;
    wire _18423;
    wire _18424;
    wire _18412;
    wire [63:0] _18409;
    wire [63:0] _18410;
    wire [62:0] _18411;
    wire [63:0] _18413;
    wire _18414;
    wire _18415;
    wire _18403;
    wire [63:0] _18400;
    wire [63:0] _18401;
    wire [62:0] _18402;
    wire [63:0] _18404;
    wire _18405;
    wire _18406;
    wire _18394;
    wire [63:0] _18391;
    wire [63:0] _18392;
    wire [62:0] _18393;
    wire [63:0] _18395;
    wire _18396;
    wire _18397;
    wire _18385;
    wire [63:0] _18382;
    wire [63:0] _18383;
    wire [62:0] _18384;
    wire [63:0] _18386;
    wire _18387;
    wire _18388;
    wire _18376;
    wire [63:0] _18373;
    wire [63:0] _18374;
    wire [62:0] _18375;
    wire [63:0] _18377;
    wire _18378;
    wire _18379;
    wire _18367;
    wire [63:0] _18364;
    wire [63:0] _18365;
    wire [62:0] _18366;
    wire [63:0] _18368;
    wire _18369;
    wire _18370;
    wire _18358;
    wire [63:0] _18355;
    wire [63:0] _18356;
    wire [62:0] _18357;
    wire [63:0] _18359;
    wire _18360;
    wire _18361;
    wire _18349;
    wire [63:0] _18346;
    wire [63:0] _18347;
    wire [62:0] _18348;
    wire [63:0] _18350;
    wire _18351;
    wire _18352;
    wire _18340;
    wire [63:0] _18337;
    wire [63:0] _18338;
    wire [62:0] _18339;
    wire [63:0] _18341;
    wire _18342;
    wire _18343;
    wire _18331;
    wire [63:0] _18328;
    wire [63:0] _18329;
    wire [62:0] _18330;
    wire [63:0] _18332;
    wire _18333;
    wire _18334;
    wire _18322;
    wire [63:0] _18319;
    wire [63:0] _18320;
    wire [62:0] _18321;
    wire [63:0] _18323;
    wire _18324;
    wire _18325;
    wire _18313;
    wire [63:0] _18310;
    wire [63:0] _18311;
    wire [62:0] _18312;
    wire [63:0] _18314;
    wire _18315;
    wire _18316;
    wire _18304;
    wire [63:0] _18301;
    wire [63:0] _18302;
    wire [62:0] _18303;
    wire [63:0] _18305;
    wire _18306;
    wire _18307;
    wire _18295;
    wire [63:0] _18292;
    wire [63:0] _18293;
    wire [62:0] _18294;
    wire [63:0] _18296;
    wire _18297;
    wire _18298;
    wire _18286;
    wire [63:0] _18283;
    wire [63:0] _18284;
    wire [62:0] _18285;
    wire [63:0] _18287;
    wire _18288;
    wire _18289;
    wire _18277;
    wire [63:0] _18274;
    wire [63:0] _18275;
    wire [62:0] _18276;
    wire [63:0] _18278;
    wire _18279;
    wire _18280;
    wire _18268;
    wire [63:0] _18265;
    wire [63:0] _18266;
    wire [62:0] _18267;
    wire [63:0] _18269;
    wire _18270;
    wire _18271;
    wire _18259;
    wire [63:0] _18256;
    wire [63:0] _18257;
    wire [62:0] _18258;
    wire [63:0] _18260;
    wire _18261;
    wire _18262;
    wire _18250;
    wire [63:0] _18247;
    wire [63:0] _18248;
    wire [62:0] _18249;
    wire [63:0] _18251;
    wire _18252;
    wire _18253;
    wire _18241;
    wire [63:0] _18238;
    wire [63:0] _18239;
    wire [62:0] _18240;
    wire [63:0] _18242;
    wire _18243;
    wire _18244;
    wire _18232;
    wire [63:0] _18229;
    wire [63:0] _18230;
    wire [62:0] _18231;
    wire [63:0] _18233;
    wire _18234;
    wire _18235;
    wire _18223;
    wire [63:0] _18220;
    wire [63:0] _18221;
    wire [62:0] _18222;
    wire [63:0] _18224;
    wire _18225;
    wire _18226;
    wire _18214;
    wire [63:0] _18211;
    wire [63:0] _18212;
    wire [62:0] _18213;
    wire [63:0] _18215;
    wire _18216;
    wire _18217;
    wire _18205;
    wire [63:0] _18202;
    wire [63:0] _18203;
    wire [62:0] _18204;
    wire [63:0] _18206;
    wire _18207;
    wire _18208;
    wire _18196;
    wire [63:0] _18193;
    wire [63:0] _18194;
    wire [62:0] _18195;
    wire [63:0] _18197;
    wire _18198;
    wire _18199;
    wire _18187;
    wire [63:0] _18184;
    wire [63:0] _18185;
    wire [62:0] _18186;
    wire [63:0] _18188;
    wire _18189;
    wire _18190;
    wire _18178;
    wire [63:0] _18175;
    wire [63:0] _18176;
    wire [62:0] _18177;
    wire [63:0] _18179;
    wire _18180;
    wire _18181;
    wire _18169;
    wire [63:0] _18166;
    wire [63:0] _18167;
    wire [62:0] _18168;
    wire [63:0] _18170;
    wire _18171;
    wire _18172;
    wire _18160;
    wire [63:0] _18157;
    wire [63:0] _18158;
    wire [62:0] _18159;
    wire [63:0] _18161;
    wire _18162;
    wire _18163;
    wire _18151;
    wire [63:0] _18148;
    wire [63:0] _18149;
    wire [62:0] _18150;
    wire [63:0] _18152;
    wire _18153;
    wire _18154;
    wire _18142;
    wire [63:0] _18139;
    wire [63:0] _18140;
    wire [62:0] _18141;
    wire [63:0] _18143;
    wire _18144;
    wire _18145;
    wire _18133;
    wire [63:0] _18130;
    wire [63:0] _18131;
    wire [62:0] _18132;
    wire [63:0] _18134;
    wire _18135;
    wire _18136;
    wire _18124;
    wire [63:0] _18121;
    wire [63:0] _18122;
    wire [62:0] _18123;
    wire [63:0] _18125;
    wire _18126;
    wire _18127;
    wire _18115;
    wire [63:0] _18112;
    wire [63:0] _18113;
    wire [62:0] _18114;
    wire [63:0] _18116;
    wire _18117;
    wire _18118;
    wire [63:0] _18105;
    wire _18106;
    wire [63:0] _18107;
    wire _18108;
    wire _18109;
    wire [63:0] _18110;
    wire [62:0] _18111;
    wire [63:0] _18119;
    wire [62:0] _18120;
    wire [63:0] _18128;
    wire [62:0] _18129;
    wire [63:0] _18137;
    wire [62:0] _18138;
    wire [63:0] _18146;
    wire [62:0] _18147;
    wire [63:0] _18155;
    wire [62:0] _18156;
    wire [63:0] _18164;
    wire [62:0] _18165;
    wire [63:0] _18173;
    wire [62:0] _18174;
    wire [63:0] _18182;
    wire [62:0] _18183;
    wire [63:0] _18191;
    wire [62:0] _18192;
    wire [63:0] _18200;
    wire [62:0] _18201;
    wire [63:0] _18209;
    wire [62:0] _18210;
    wire [63:0] _18218;
    wire [62:0] _18219;
    wire [63:0] _18227;
    wire [62:0] _18228;
    wire [63:0] _18236;
    wire [62:0] _18237;
    wire [63:0] _18245;
    wire [62:0] _18246;
    wire [63:0] _18254;
    wire [62:0] _18255;
    wire [63:0] _18263;
    wire [62:0] _18264;
    wire [63:0] _18272;
    wire [62:0] _18273;
    wire [63:0] _18281;
    wire [62:0] _18282;
    wire [63:0] _18290;
    wire [62:0] _18291;
    wire [63:0] _18299;
    wire [62:0] _18300;
    wire [63:0] _18308;
    wire [62:0] _18309;
    wire [63:0] _18317;
    wire [62:0] _18318;
    wire [63:0] _18326;
    wire [62:0] _18327;
    wire [63:0] _18335;
    wire [62:0] _18336;
    wire [63:0] _18344;
    wire [62:0] _18345;
    wire [63:0] _18353;
    wire [62:0] _18354;
    wire [63:0] _18362;
    wire [62:0] _18363;
    wire [63:0] _18371;
    wire [62:0] _18372;
    wire [63:0] _18380;
    wire [62:0] _18381;
    wire [63:0] _18389;
    wire [62:0] _18390;
    wire [63:0] _18398;
    wire [62:0] _18399;
    wire [63:0] _18407;
    wire [62:0] _18408;
    wire [63:0] _18416;
    wire [62:0] _18417;
    wire [63:0] _18425;
    wire [62:0] _18426;
    wire [63:0] _18434;
    wire [62:0] _18435;
    wire [63:0] _18443;
    wire [62:0] _18444;
    wire [63:0] _18452;
    wire [62:0] _18453;
    wire [63:0] _18461;
    wire [62:0] _18462;
    wire [63:0] _18470;
    wire [62:0] _18471;
    wire [63:0] _18479;
    wire [62:0] _18480;
    wire [63:0] _18488;
    wire [62:0] _18489;
    wire [63:0] _18497;
    wire [62:0] _18498;
    wire [63:0] _18506;
    wire [62:0] _18507;
    wire [63:0] _18515;
    wire [62:0] _18516;
    wire [63:0] _18524;
    wire [62:0] _18525;
    wire [63:0] _18533;
    wire [62:0] _18534;
    wire [63:0] _18542;
    wire [62:0] _18543;
    wire [63:0] _18551;
    wire [62:0] _18552;
    wire [63:0] _18560;
    wire [62:0] _18561;
    wire [63:0] _18569;
    wire [62:0] _18570;
    wire [63:0] _18578;
    wire [62:0] _18579;
    wire [63:0] _18587;
    wire [62:0] _18588;
    wire [63:0] _18596;
    wire [62:0] _18597;
    wire [63:0] _18605;
    wire [62:0] _18606;
    wire [63:0] _18614;
    wire [62:0] _18615;
    wire [63:0] _18623;
    wire [62:0] _18624;
    wire [63:0] _18632;
    wire [62:0] _18633;
    wire [63:0] _18641;
    wire [62:0] _18642;
    wire [63:0] _18650;
    wire [62:0] _18651;
    wire [63:0] _18659;
    wire [62:0] _18660;
    wire [63:0] _18668;
    wire [62:0] _18669;
    wire [63:0] _18677;
    wire [63:0] _18679;
    wire [127:0] _18680;
    wire [63:0] _18681;
    wire [63:0] _19263;
    wire _18091;
    wire [63:0] _18088;
    wire [63:0] _18089;
    wire [62:0] _18090;
    wire [63:0] _18092;
    wire _18093;
    wire _18094;
    wire _18082;
    wire [63:0] _18079;
    wire [63:0] _18080;
    wire [62:0] _18081;
    wire [63:0] _18083;
    wire _18084;
    wire _18085;
    wire _18073;
    wire [63:0] _18070;
    wire [63:0] _18071;
    wire [62:0] _18072;
    wire [63:0] _18074;
    wire _18075;
    wire _18076;
    wire _18064;
    wire [63:0] _18061;
    wire [63:0] _18062;
    wire [62:0] _18063;
    wire [63:0] _18065;
    wire _18066;
    wire _18067;
    wire _18055;
    wire [63:0] _18052;
    wire [63:0] _18053;
    wire [62:0] _18054;
    wire [63:0] _18056;
    wire _18057;
    wire _18058;
    wire _18046;
    wire [63:0] _18043;
    wire [63:0] _18044;
    wire [62:0] _18045;
    wire [63:0] _18047;
    wire _18048;
    wire _18049;
    wire _18037;
    wire [63:0] _18034;
    wire [63:0] _18035;
    wire [62:0] _18036;
    wire [63:0] _18038;
    wire _18039;
    wire _18040;
    wire _18028;
    wire [63:0] _18025;
    wire [63:0] _18026;
    wire [62:0] _18027;
    wire [63:0] _18029;
    wire _18030;
    wire _18031;
    wire _18019;
    wire [63:0] _18016;
    wire [63:0] _18017;
    wire [62:0] _18018;
    wire [63:0] _18020;
    wire _18021;
    wire _18022;
    wire _18010;
    wire [63:0] _18007;
    wire [63:0] _18008;
    wire [62:0] _18009;
    wire [63:0] _18011;
    wire _18012;
    wire _18013;
    wire _18001;
    wire [63:0] _17998;
    wire [63:0] _17999;
    wire [62:0] _18000;
    wire [63:0] _18002;
    wire _18003;
    wire _18004;
    wire _17992;
    wire [63:0] _17989;
    wire [63:0] _17990;
    wire [62:0] _17991;
    wire [63:0] _17993;
    wire _17994;
    wire _17995;
    wire _17983;
    wire [63:0] _17980;
    wire [63:0] _17981;
    wire [62:0] _17982;
    wire [63:0] _17984;
    wire _17985;
    wire _17986;
    wire _17974;
    wire [63:0] _17971;
    wire [63:0] _17972;
    wire [62:0] _17973;
    wire [63:0] _17975;
    wire _17976;
    wire _17977;
    wire _17965;
    wire [63:0] _17962;
    wire [63:0] _17963;
    wire [62:0] _17964;
    wire [63:0] _17966;
    wire _17967;
    wire _17968;
    wire _17956;
    wire [63:0] _17953;
    wire [63:0] _17954;
    wire [62:0] _17955;
    wire [63:0] _17957;
    wire _17958;
    wire _17959;
    wire _17947;
    wire [63:0] _17944;
    wire [63:0] _17945;
    wire [62:0] _17946;
    wire [63:0] _17948;
    wire _17949;
    wire _17950;
    wire _17938;
    wire [63:0] _17935;
    wire [63:0] _17936;
    wire [62:0] _17937;
    wire [63:0] _17939;
    wire _17940;
    wire _17941;
    wire _17929;
    wire [63:0] _17926;
    wire [63:0] _17927;
    wire [62:0] _17928;
    wire [63:0] _17930;
    wire _17931;
    wire _17932;
    wire _17920;
    wire [63:0] _17917;
    wire [63:0] _17918;
    wire [62:0] _17919;
    wire [63:0] _17921;
    wire _17922;
    wire _17923;
    wire _17911;
    wire [63:0] _17908;
    wire [63:0] _17909;
    wire [62:0] _17910;
    wire [63:0] _17912;
    wire _17913;
    wire _17914;
    wire _17902;
    wire [63:0] _17899;
    wire [63:0] _17900;
    wire [62:0] _17901;
    wire [63:0] _17903;
    wire _17904;
    wire _17905;
    wire _17893;
    wire [63:0] _17890;
    wire [63:0] _17891;
    wire [62:0] _17892;
    wire [63:0] _17894;
    wire _17895;
    wire _17896;
    wire _17884;
    wire [63:0] _17881;
    wire [63:0] _17882;
    wire [62:0] _17883;
    wire [63:0] _17885;
    wire _17886;
    wire _17887;
    wire _17875;
    wire [63:0] _17872;
    wire [63:0] _17873;
    wire [62:0] _17874;
    wire [63:0] _17876;
    wire _17877;
    wire _17878;
    wire _17866;
    wire [63:0] _17863;
    wire [63:0] _17864;
    wire [62:0] _17865;
    wire [63:0] _17867;
    wire _17868;
    wire _17869;
    wire _17857;
    wire [63:0] _17854;
    wire [63:0] _17855;
    wire [62:0] _17856;
    wire [63:0] _17858;
    wire _17859;
    wire _17860;
    wire _17848;
    wire [63:0] _17845;
    wire [63:0] _17846;
    wire [62:0] _17847;
    wire [63:0] _17849;
    wire _17850;
    wire _17851;
    wire _17839;
    wire [63:0] _17836;
    wire [63:0] _17837;
    wire [62:0] _17838;
    wire [63:0] _17840;
    wire _17841;
    wire _17842;
    wire _17830;
    wire [63:0] _17827;
    wire [63:0] _17828;
    wire [62:0] _17829;
    wire [63:0] _17831;
    wire _17832;
    wire _17833;
    wire _17821;
    wire [63:0] _17818;
    wire [63:0] _17819;
    wire [62:0] _17820;
    wire [63:0] _17822;
    wire _17823;
    wire _17824;
    wire _17812;
    wire [63:0] _17809;
    wire [63:0] _17810;
    wire [62:0] _17811;
    wire [63:0] _17813;
    wire _17814;
    wire _17815;
    wire _17803;
    wire [63:0] _17800;
    wire [63:0] _17801;
    wire [62:0] _17802;
    wire [63:0] _17804;
    wire _17805;
    wire _17806;
    wire _17794;
    wire [63:0] _17791;
    wire [63:0] _17792;
    wire [62:0] _17793;
    wire [63:0] _17795;
    wire _17796;
    wire _17797;
    wire _17785;
    wire [63:0] _17782;
    wire [63:0] _17783;
    wire [62:0] _17784;
    wire [63:0] _17786;
    wire _17787;
    wire _17788;
    wire _17776;
    wire [63:0] _17773;
    wire [63:0] _17774;
    wire [62:0] _17775;
    wire [63:0] _17777;
    wire _17778;
    wire _17779;
    wire _17767;
    wire [63:0] _17764;
    wire [63:0] _17765;
    wire [62:0] _17766;
    wire [63:0] _17768;
    wire _17769;
    wire _17770;
    wire _17758;
    wire [63:0] _17755;
    wire [63:0] _17756;
    wire [62:0] _17757;
    wire [63:0] _17759;
    wire _17760;
    wire _17761;
    wire _17749;
    wire [63:0] _17746;
    wire [63:0] _17747;
    wire [62:0] _17748;
    wire [63:0] _17750;
    wire _17751;
    wire _17752;
    wire _17740;
    wire [63:0] _17737;
    wire [63:0] _17738;
    wire [62:0] _17739;
    wire [63:0] _17741;
    wire _17742;
    wire _17743;
    wire _17731;
    wire [63:0] _17728;
    wire [63:0] _17729;
    wire [62:0] _17730;
    wire [63:0] _17732;
    wire _17733;
    wire _17734;
    wire _17722;
    wire [63:0] _17719;
    wire [63:0] _17720;
    wire [62:0] _17721;
    wire [63:0] _17723;
    wire _17724;
    wire _17725;
    wire _17713;
    wire [63:0] _17710;
    wire [63:0] _17711;
    wire [62:0] _17712;
    wire [63:0] _17714;
    wire _17715;
    wire _17716;
    wire _17704;
    wire [63:0] _17701;
    wire [63:0] _17702;
    wire [62:0] _17703;
    wire [63:0] _17705;
    wire _17706;
    wire _17707;
    wire _17695;
    wire [63:0] _17692;
    wire [63:0] _17693;
    wire [62:0] _17694;
    wire [63:0] _17696;
    wire _17697;
    wire _17698;
    wire _17686;
    wire [63:0] _17683;
    wire [63:0] _17684;
    wire [62:0] _17685;
    wire [63:0] _17687;
    wire _17688;
    wire _17689;
    wire _17677;
    wire [63:0] _17674;
    wire [63:0] _17675;
    wire [62:0] _17676;
    wire [63:0] _17678;
    wire _17679;
    wire _17680;
    wire _17668;
    wire [63:0] _17665;
    wire [63:0] _17666;
    wire [62:0] _17667;
    wire [63:0] _17669;
    wire _17670;
    wire _17671;
    wire _17659;
    wire [63:0] _17656;
    wire [63:0] _17657;
    wire [62:0] _17658;
    wire [63:0] _17660;
    wire _17661;
    wire _17662;
    wire _17650;
    wire [63:0] _17647;
    wire [63:0] _17648;
    wire [62:0] _17649;
    wire [63:0] _17651;
    wire _17652;
    wire _17653;
    wire _17641;
    wire [63:0] _17638;
    wire [63:0] _17639;
    wire [62:0] _17640;
    wire [63:0] _17642;
    wire _17643;
    wire _17644;
    wire _17632;
    wire [63:0] _17629;
    wire [63:0] _17630;
    wire [62:0] _17631;
    wire [63:0] _17633;
    wire _17634;
    wire _17635;
    wire _17623;
    wire [63:0] _17620;
    wire [63:0] _17621;
    wire [62:0] _17622;
    wire [63:0] _17624;
    wire _17625;
    wire _17626;
    wire _17614;
    wire [63:0] _17611;
    wire [63:0] _17612;
    wire [62:0] _17613;
    wire [63:0] _17615;
    wire _17616;
    wire _17617;
    wire _17605;
    wire [63:0] _17602;
    wire [63:0] _17603;
    wire [62:0] _17604;
    wire [63:0] _17606;
    wire _17607;
    wire _17608;
    wire _17596;
    wire [63:0] _17593;
    wire [63:0] _17594;
    wire [62:0] _17595;
    wire [63:0] _17597;
    wire _17598;
    wire _17599;
    wire _17587;
    wire [63:0] _17584;
    wire [63:0] _17585;
    wire [62:0] _17586;
    wire [63:0] _17588;
    wire _17589;
    wire _17590;
    wire _17578;
    wire [63:0] _17575;
    wire [63:0] _17576;
    wire [62:0] _17577;
    wire [63:0] _17579;
    wire _17580;
    wire _17581;
    wire _17569;
    wire [63:0] _17566;
    wire [63:0] _17567;
    wire [62:0] _17568;
    wire [63:0] _17570;
    wire _17571;
    wire _17572;
    wire _17560;
    wire [63:0] _17557;
    wire [63:0] _17558;
    wire [62:0] _17559;
    wire [63:0] _17561;
    wire _17562;
    wire _17563;
    wire _17551;
    wire [63:0] _17548;
    wire [63:0] _17549;
    wire [62:0] _17550;
    wire [63:0] _17552;
    wire _17553;
    wire _17554;
    wire _17542;
    wire [63:0] _17539;
    wire [63:0] _17540;
    wire [62:0] _17541;
    wire [63:0] _17543;
    wire _17544;
    wire _17545;
    wire _17533;
    wire [63:0] _17530;
    wire [63:0] _17531;
    wire [62:0] _17532;
    wire [63:0] _17534;
    wire _17535;
    wire _17536;
    wire [63:0] _17525;
    wire [63:0] _17521;
    wire [63:0] _17522;
    wire _17523;
    wire [63:0] _17524;
    wire _17526;
    wire _17527;
    wire [63:0] _17528;
    wire [62:0] _17529;
    wire [63:0] _17537;
    wire [62:0] _17538;
    wire [63:0] _17546;
    wire [62:0] _17547;
    wire [63:0] _17555;
    wire [62:0] _17556;
    wire [63:0] _17564;
    wire [62:0] _17565;
    wire [63:0] _17573;
    wire [62:0] _17574;
    wire [63:0] _17582;
    wire [62:0] _17583;
    wire [63:0] _17591;
    wire [62:0] _17592;
    wire [63:0] _17600;
    wire [62:0] _17601;
    wire [63:0] _17609;
    wire [62:0] _17610;
    wire [63:0] _17618;
    wire [62:0] _17619;
    wire [63:0] _17627;
    wire [62:0] _17628;
    wire [63:0] _17636;
    wire [62:0] _17637;
    wire [63:0] _17645;
    wire [62:0] _17646;
    wire [63:0] _17654;
    wire [62:0] _17655;
    wire [63:0] _17663;
    wire [62:0] _17664;
    wire [63:0] _17672;
    wire [62:0] _17673;
    wire [63:0] _17681;
    wire [62:0] _17682;
    wire [63:0] _17690;
    wire [62:0] _17691;
    wire [63:0] _17699;
    wire [62:0] _17700;
    wire [63:0] _17708;
    wire [62:0] _17709;
    wire [63:0] _17717;
    wire [62:0] _17718;
    wire [63:0] _17726;
    wire [62:0] _17727;
    wire [63:0] _17735;
    wire [62:0] _17736;
    wire [63:0] _17744;
    wire [62:0] _17745;
    wire [63:0] _17753;
    wire [62:0] _17754;
    wire [63:0] _17762;
    wire [62:0] _17763;
    wire [63:0] _17771;
    wire [62:0] _17772;
    wire [63:0] _17780;
    wire [62:0] _17781;
    wire [63:0] _17789;
    wire [62:0] _17790;
    wire [63:0] _17798;
    wire [62:0] _17799;
    wire [63:0] _17807;
    wire [62:0] _17808;
    wire [63:0] _17816;
    wire [62:0] _17817;
    wire [63:0] _17825;
    wire [62:0] _17826;
    wire [63:0] _17834;
    wire [62:0] _17835;
    wire [63:0] _17843;
    wire [62:0] _17844;
    wire [63:0] _17852;
    wire [62:0] _17853;
    wire [63:0] _17861;
    wire [62:0] _17862;
    wire [63:0] _17870;
    wire [62:0] _17871;
    wire [63:0] _17879;
    wire [62:0] _17880;
    wire [63:0] _17888;
    wire [62:0] _17889;
    wire [63:0] _17897;
    wire [62:0] _17898;
    wire [63:0] _17906;
    wire [62:0] _17907;
    wire [63:0] _17915;
    wire [62:0] _17916;
    wire [63:0] _17924;
    wire [62:0] _17925;
    wire [63:0] _17933;
    wire [62:0] _17934;
    wire [63:0] _17942;
    wire [62:0] _17943;
    wire [63:0] _17951;
    wire [62:0] _17952;
    wire [63:0] _17960;
    wire [62:0] _17961;
    wire [63:0] _17969;
    wire [62:0] _17970;
    wire [63:0] _17978;
    wire [62:0] _17979;
    wire [63:0] _17987;
    wire [62:0] _17988;
    wire [63:0] _17996;
    wire [62:0] _17997;
    wire [63:0] _18005;
    wire [62:0] _18006;
    wire [63:0] _18014;
    wire [62:0] _18015;
    wire [63:0] _18023;
    wire [62:0] _18024;
    wire [63:0] _18032;
    wire [62:0] _18033;
    wire [63:0] _18041;
    wire [62:0] _18042;
    wire [63:0] _18050;
    wire [62:0] _18051;
    wire [63:0] _18059;
    wire [62:0] _18060;
    wire [63:0] _18068;
    wire [62:0] _18069;
    wire [63:0] _18077;
    wire [62:0] _18078;
    wire [63:0] _18086;
    wire [62:0] _18087;
    wire [63:0] _18095;
    wire [127:0] _18096;
    wire [63:0] _18097;
    wire [63:0] _17518;
    wire _18098;
    wire [63:0] _18099;
    wire _17516;
    wire [63:0] _17517;
    wire _18100;
    wire _18101;
    wire [63:0] _19264;
    wire _17505;
    wire [63:0] _17502;
    wire [63:0] _17503;
    wire [62:0] _17504;
    wire [63:0] _17506;
    wire _17507;
    wire _17508;
    wire _17496;
    wire [63:0] _17493;
    wire [63:0] _17494;
    wire [62:0] _17495;
    wire [63:0] _17497;
    wire _17498;
    wire _17499;
    wire _17487;
    wire [63:0] _17484;
    wire [63:0] _17485;
    wire [62:0] _17486;
    wire [63:0] _17488;
    wire _17489;
    wire _17490;
    wire _17478;
    wire [63:0] _17475;
    wire [63:0] _17476;
    wire [62:0] _17477;
    wire [63:0] _17479;
    wire _17480;
    wire _17481;
    wire _17469;
    wire [63:0] _17466;
    wire [63:0] _17467;
    wire [62:0] _17468;
    wire [63:0] _17470;
    wire _17471;
    wire _17472;
    wire _17460;
    wire [63:0] _17457;
    wire [63:0] _17458;
    wire [62:0] _17459;
    wire [63:0] _17461;
    wire _17462;
    wire _17463;
    wire _17451;
    wire [63:0] _17448;
    wire [63:0] _17449;
    wire [62:0] _17450;
    wire [63:0] _17452;
    wire _17453;
    wire _17454;
    wire _17442;
    wire [63:0] _17439;
    wire [63:0] _17440;
    wire [62:0] _17441;
    wire [63:0] _17443;
    wire _17444;
    wire _17445;
    wire _17433;
    wire [63:0] _17430;
    wire [63:0] _17431;
    wire [62:0] _17432;
    wire [63:0] _17434;
    wire _17435;
    wire _17436;
    wire _17424;
    wire [63:0] _17421;
    wire [63:0] _17422;
    wire [62:0] _17423;
    wire [63:0] _17425;
    wire _17426;
    wire _17427;
    wire _17415;
    wire [63:0] _17412;
    wire [63:0] _17413;
    wire [62:0] _17414;
    wire [63:0] _17416;
    wire _17417;
    wire _17418;
    wire _17406;
    wire [63:0] _17403;
    wire [63:0] _17404;
    wire [62:0] _17405;
    wire [63:0] _17407;
    wire _17408;
    wire _17409;
    wire _17397;
    wire [63:0] _17394;
    wire [63:0] _17395;
    wire [62:0] _17396;
    wire [63:0] _17398;
    wire _17399;
    wire _17400;
    wire _17388;
    wire [63:0] _17385;
    wire [63:0] _17386;
    wire [62:0] _17387;
    wire [63:0] _17389;
    wire _17390;
    wire _17391;
    wire _17379;
    wire [63:0] _17376;
    wire [63:0] _17377;
    wire [62:0] _17378;
    wire [63:0] _17380;
    wire _17381;
    wire _17382;
    wire _17370;
    wire [63:0] _17367;
    wire [63:0] _17368;
    wire [62:0] _17369;
    wire [63:0] _17371;
    wire _17372;
    wire _17373;
    wire _17361;
    wire [63:0] _17358;
    wire [63:0] _17359;
    wire [62:0] _17360;
    wire [63:0] _17362;
    wire _17363;
    wire _17364;
    wire _17352;
    wire [63:0] _17349;
    wire [63:0] _17350;
    wire [62:0] _17351;
    wire [63:0] _17353;
    wire _17354;
    wire _17355;
    wire _17343;
    wire [63:0] _17340;
    wire [63:0] _17341;
    wire [62:0] _17342;
    wire [63:0] _17344;
    wire _17345;
    wire _17346;
    wire _17334;
    wire [63:0] _17331;
    wire [63:0] _17332;
    wire [62:0] _17333;
    wire [63:0] _17335;
    wire _17336;
    wire _17337;
    wire _17325;
    wire [63:0] _17322;
    wire [63:0] _17323;
    wire [62:0] _17324;
    wire [63:0] _17326;
    wire _17327;
    wire _17328;
    wire _17316;
    wire [63:0] _17313;
    wire [63:0] _17314;
    wire [62:0] _17315;
    wire [63:0] _17317;
    wire _17318;
    wire _17319;
    wire _17307;
    wire [63:0] _17304;
    wire [63:0] _17305;
    wire [62:0] _17306;
    wire [63:0] _17308;
    wire _17309;
    wire _17310;
    wire _17298;
    wire [63:0] _17295;
    wire [63:0] _17296;
    wire [62:0] _17297;
    wire [63:0] _17299;
    wire _17300;
    wire _17301;
    wire _17289;
    wire [63:0] _17286;
    wire [63:0] _17287;
    wire [62:0] _17288;
    wire [63:0] _17290;
    wire _17291;
    wire _17292;
    wire _17280;
    wire [63:0] _17277;
    wire [63:0] _17278;
    wire [62:0] _17279;
    wire [63:0] _17281;
    wire _17282;
    wire _17283;
    wire _17271;
    wire [63:0] _17268;
    wire [63:0] _17269;
    wire [62:0] _17270;
    wire [63:0] _17272;
    wire _17273;
    wire _17274;
    wire _17262;
    wire [63:0] _17259;
    wire [63:0] _17260;
    wire [62:0] _17261;
    wire [63:0] _17263;
    wire _17264;
    wire _17265;
    wire _17253;
    wire [63:0] _17250;
    wire [63:0] _17251;
    wire [62:0] _17252;
    wire [63:0] _17254;
    wire _17255;
    wire _17256;
    wire _17244;
    wire [63:0] _17241;
    wire [63:0] _17242;
    wire [62:0] _17243;
    wire [63:0] _17245;
    wire _17246;
    wire _17247;
    wire _17235;
    wire [63:0] _17232;
    wire [63:0] _17233;
    wire [62:0] _17234;
    wire [63:0] _17236;
    wire _17237;
    wire _17238;
    wire _17226;
    wire [63:0] _17223;
    wire [63:0] _17224;
    wire [62:0] _17225;
    wire [63:0] _17227;
    wire _17228;
    wire _17229;
    wire _17217;
    wire [63:0] _17214;
    wire [63:0] _17215;
    wire [62:0] _17216;
    wire [63:0] _17218;
    wire _17219;
    wire _17220;
    wire _17208;
    wire [63:0] _17205;
    wire [63:0] _17206;
    wire [62:0] _17207;
    wire [63:0] _17209;
    wire _17210;
    wire _17211;
    wire _17199;
    wire [63:0] _17196;
    wire [63:0] _17197;
    wire [62:0] _17198;
    wire [63:0] _17200;
    wire _17201;
    wire _17202;
    wire _17190;
    wire [63:0] _17187;
    wire [63:0] _17188;
    wire [62:0] _17189;
    wire [63:0] _17191;
    wire _17192;
    wire _17193;
    wire _17181;
    wire [63:0] _17178;
    wire [63:0] _17179;
    wire [62:0] _17180;
    wire [63:0] _17182;
    wire _17183;
    wire _17184;
    wire _17172;
    wire [63:0] _17169;
    wire [63:0] _17170;
    wire [62:0] _17171;
    wire [63:0] _17173;
    wire _17174;
    wire _17175;
    wire _17163;
    wire [63:0] _17160;
    wire [63:0] _17161;
    wire [62:0] _17162;
    wire [63:0] _17164;
    wire _17165;
    wire _17166;
    wire _17154;
    wire [63:0] _17151;
    wire [63:0] _17152;
    wire [62:0] _17153;
    wire [63:0] _17155;
    wire _17156;
    wire _17157;
    wire _17145;
    wire [63:0] _17142;
    wire [63:0] _17143;
    wire [62:0] _17144;
    wire [63:0] _17146;
    wire _17147;
    wire _17148;
    wire _17136;
    wire [63:0] _17133;
    wire [63:0] _17134;
    wire [62:0] _17135;
    wire [63:0] _17137;
    wire _17138;
    wire _17139;
    wire _17127;
    wire [63:0] _17124;
    wire [63:0] _17125;
    wire [62:0] _17126;
    wire [63:0] _17128;
    wire _17129;
    wire _17130;
    wire _17118;
    wire [63:0] _17115;
    wire [63:0] _17116;
    wire [62:0] _17117;
    wire [63:0] _17119;
    wire _17120;
    wire _17121;
    wire _17109;
    wire [63:0] _17106;
    wire [63:0] _17107;
    wire [62:0] _17108;
    wire [63:0] _17110;
    wire _17111;
    wire _17112;
    wire _17100;
    wire [63:0] _17097;
    wire [63:0] _17098;
    wire [62:0] _17099;
    wire [63:0] _17101;
    wire _17102;
    wire _17103;
    wire _17091;
    wire [63:0] _17088;
    wire [63:0] _17089;
    wire [62:0] _17090;
    wire [63:0] _17092;
    wire _17093;
    wire _17094;
    wire _17082;
    wire [63:0] _17079;
    wire [63:0] _17080;
    wire [62:0] _17081;
    wire [63:0] _17083;
    wire _17084;
    wire _17085;
    wire _17073;
    wire [63:0] _17070;
    wire [63:0] _17071;
    wire [62:0] _17072;
    wire [63:0] _17074;
    wire _17075;
    wire _17076;
    wire _17064;
    wire [63:0] _17061;
    wire [63:0] _17062;
    wire [62:0] _17063;
    wire [63:0] _17065;
    wire _17066;
    wire _17067;
    wire _17055;
    wire [63:0] _17052;
    wire [63:0] _17053;
    wire [62:0] _17054;
    wire [63:0] _17056;
    wire _17057;
    wire _17058;
    wire _17046;
    wire [63:0] _17043;
    wire [63:0] _17044;
    wire [62:0] _17045;
    wire [63:0] _17047;
    wire _17048;
    wire _17049;
    wire _17037;
    wire [63:0] _17034;
    wire [63:0] _17035;
    wire [62:0] _17036;
    wire [63:0] _17038;
    wire _17039;
    wire _17040;
    wire _17028;
    wire [63:0] _17025;
    wire [63:0] _17026;
    wire [62:0] _17027;
    wire [63:0] _17029;
    wire _17030;
    wire _17031;
    wire _17019;
    wire [63:0] _17016;
    wire [63:0] _17017;
    wire [62:0] _17018;
    wire [63:0] _17020;
    wire _17021;
    wire _17022;
    wire _17010;
    wire [63:0] _17007;
    wire [63:0] _17008;
    wire [62:0] _17009;
    wire [63:0] _17011;
    wire _17012;
    wire _17013;
    wire _17001;
    wire [63:0] _16998;
    wire [63:0] _16999;
    wire [62:0] _17000;
    wire [63:0] _17002;
    wire _17003;
    wire _17004;
    wire _16992;
    wire [63:0] _16989;
    wire [63:0] _16990;
    wire [62:0] _16991;
    wire [63:0] _16993;
    wire _16994;
    wire _16995;
    wire _16983;
    wire [63:0] _16980;
    wire [63:0] _16981;
    wire [62:0] _16982;
    wire [63:0] _16984;
    wire _16985;
    wire _16986;
    wire _16974;
    wire [63:0] _16971;
    wire [63:0] _16972;
    wire [62:0] _16973;
    wire [63:0] _16975;
    wire _16976;
    wire _16977;
    wire _16965;
    wire [63:0] _16962;
    wire [63:0] _16963;
    wire [62:0] _16964;
    wire [63:0] _16966;
    wire _16967;
    wire _16968;
    wire _16956;
    wire [63:0] _16953;
    wire [63:0] _16954;
    wire [62:0] _16955;
    wire [63:0] _16957;
    wire _16958;
    wire _16959;
    wire _16947;
    wire [63:0] _16944;
    wire [63:0] _16945;
    wire [62:0] _16946;
    wire [63:0] _16948;
    wire _16949;
    wire _16950;
    wire [63:0] _16934;
    wire [127:0] _16935;
    wire [63:0] _16936;
    wire _16937;
    wire [63:0] _16938;
    wire _16940;
    wire _16941;
    wire [63:0] _16942;
    wire [62:0] _16943;
    wire [63:0] _16951;
    wire [62:0] _16952;
    wire [63:0] _16960;
    wire [62:0] _16961;
    wire [63:0] _16969;
    wire [62:0] _16970;
    wire [63:0] _16978;
    wire [62:0] _16979;
    wire [63:0] _16987;
    wire [62:0] _16988;
    wire [63:0] _16996;
    wire [62:0] _16997;
    wire [63:0] _17005;
    wire [62:0] _17006;
    wire [63:0] _17014;
    wire [62:0] _17015;
    wire [63:0] _17023;
    wire [62:0] _17024;
    wire [63:0] _17032;
    wire [62:0] _17033;
    wire [63:0] _17041;
    wire [62:0] _17042;
    wire [63:0] _17050;
    wire [62:0] _17051;
    wire [63:0] _17059;
    wire [62:0] _17060;
    wire [63:0] _17068;
    wire [62:0] _17069;
    wire [63:0] _17077;
    wire [62:0] _17078;
    wire [63:0] _17086;
    wire [62:0] _17087;
    wire [63:0] _17095;
    wire [62:0] _17096;
    wire [63:0] _17104;
    wire [62:0] _17105;
    wire [63:0] _17113;
    wire [62:0] _17114;
    wire [63:0] _17122;
    wire [62:0] _17123;
    wire [63:0] _17131;
    wire [62:0] _17132;
    wire [63:0] _17140;
    wire [62:0] _17141;
    wire [63:0] _17149;
    wire [62:0] _17150;
    wire [63:0] _17158;
    wire [62:0] _17159;
    wire [63:0] _17167;
    wire [62:0] _17168;
    wire [63:0] _17176;
    wire [62:0] _17177;
    wire [63:0] _17185;
    wire [62:0] _17186;
    wire [63:0] _17194;
    wire [62:0] _17195;
    wire [63:0] _17203;
    wire [62:0] _17204;
    wire [63:0] _17212;
    wire [62:0] _17213;
    wire [63:0] _17221;
    wire [62:0] _17222;
    wire [63:0] _17230;
    wire [62:0] _17231;
    wire [63:0] _17239;
    wire [62:0] _17240;
    wire [63:0] _17248;
    wire [62:0] _17249;
    wire [63:0] _17257;
    wire [62:0] _17258;
    wire [63:0] _17266;
    wire [62:0] _17267;
    wire [63:0] _17275;
    wire [62:0] _17276;
    wire [63:0] _17284;
    wire [62:0] _17285;
    wire [63:0] _17293;
    wire [62:0] _17294;
    wire [63:0] _17302;
    wire [62:0] _17303;
    wire [63:0] _17311;
    wire [62:0] _17312;
    wire [63:0] _17320;
    wire [62:0] _17321;
    wire [63:0] _17329;
    wire [62:0] _17330;
    wire [63:0] _17338;
    wire [62:0] _17339;
    wire [63:0] _17347;
    wire [62:0] _17348;
    wire [63:0] _17356;
    wire [62:0] _17357;
    wire [63:0] _17365;
    wire [62:0] _17366;
    wire [63:0] _17374;
    wire [62:0] _17375;
    wire [63:0] _17383;
    wire [62:0] _17384;
    wire [63:0] _17392;
    wire [62:0] _17393;
    wire [63:0] _17401;
    wire [62:0] _17402;
    wire [63:0] _17410;
    wire [62:0] _17411;
    wire [63:0] _17419;
    wire [62:0] _17420;
    wire [63:0] _17428;
    wire [62:0] _17429;
    wire [63:0] _17437;
    wire [62:0] _17438;
    wire [63:0] _17446;
    wire [62:0] _17447;
    wire [63:0] _17455;
    wire [62:0] _17456;
    wire [63:0] _17464;
    wire [62:0] _17465;
    wire [63:0] _17473;
    wire [62:0] _17474;
    wire [63:0] _17482;
    wire [62:0] _17483;
    wire [63:0] _17491;
    wire [62:0] _17492;
    wire [63:0] _17500;
    wire [62:0] _17501;
    wire [63:0] _17509;
    wire [127:0] _17510;
    wire [63:0] _17511;
    wire _16922;
    wire [63:0] _16919;
    wire [63:0] _16920;
    wire [62:0] _16921;
    wire [63:0] _16923;
    wire _16924;
    wire _16925;
    wire _16913;
    wire [63:0] _16910;
    wire [63:0] _16911;
    wire [62:0] _16912;
    wire [63:0] _16914;
    wire _16915;
    wire _16916;
    wire _16904;
    wire [63:0] _16901;
    wire [63:0] _16902;
    wire [62:0] _16903;
    wire [63:0] _16905;
    wire _16906;
    wire _16907;
    wire _16895;
    wire [63:0] _16892;
    wire [63:0] _16893;
    wire [62:0] _16894;
    wire [63:0] _16896;
    wire _16897;
    wire _16898;
    wire _16886;
    wire [63:0] _16883;
    wire [63:0] _16884;
    wire [62:0] _16885;
    wire [63:0] _16887;
    wire _16888;
    wire _16889;
    wire _16877;
    wire [63:0] _16874;
    wire [63:0] _16875;
    wire [62:0] _16876;
    wire [63:0] _16878;
    wire _16879;
    wire _16880;
    wire _16868;
    wire [63:0] _16865;
    wire [63:0] _16866;
    wire [62:0] _16867;
    wire [63:0] _16869;
    wire _16870;
    wire _16871;
    wire _16859;
    wire [63:0] _16856;
    wire [63:0] _16857;
    wire [62:0] _16858;
    wire [63:0] _16860;
    wire _16861;
    wire _16862;
    wire _16850;
    wire [63:0] _16847;
    wire [63:0] _16848;
    wire [62:0] _16849;
    wire [63:0] _16851;
    wire _16852;
    wire _16853;
    wire _16841;
    wire [63:0] _16838;
    wire [63:0] _16839;
    wire [62:0] _16840;
    wire [63:0] _16842;
    wire _16843;
    wire _16844;
    wire _16832;
    wire [63:0] _16829;
    wire [63:0] _16830;
    wire [62:0] _16831;
    wire [63:0] _16833;
    wire _16834;
    wire _16835;
    wire _16823;
    wire [63:0] _16820;
    wire [63:0] _16821;
    wire [62:0] _16822;
    wire [63:0] _16824;
    wire _16825;
    wire _16826;
    wire _16814;
    wire [63:0] _16811;
    wire [63:0] _16812;
    wire [62:0] _16813;
    wire [63:0] _16815;
    wire _16816;
    wire _16817;
    wire _16805;
    wire [63:0] _16802;
    wire [63:0] _16803;
    wire [62:0] _16804;
    wire [63:0] _16806;
    wire _16807;
    wire _16808;
    wire _16796;
    wire [63:0] _16793;
    wire [63:0] _16794;
    wire [62:0] _16795;
    wire [63:0] _16797;
    wire _16798;
    wire _16799;
    wire _16787;
    wire [63:0] _16784;
    wire [63:0] _16785;
    wire [62:0] _16786;
    wire [63:0] _16788;
    wire _16789;
    wire _16790;
    wire _16778;
    wire [63:0] _16775;
    wire [63:0] _16776;
    wire [62:0] _16777;
    wire [63:0] _16779;
    wire _16780;
    wire _16781;
    wire _16769;
    wire [63:0] _16766;
    wire [63:0] _16767;
    wire [62:0] _16768;
    wire [63:0] _16770;
    wire _16771;
    wire _16772;
    wire _16760;
    wire [63:0] _16757;
    wire [63:0] _16758;
    wire [62:0] _16759;
    wire [63:0] _16761;
    wire _16762;
    wire _16763;
    wire _16751;
    wire [63:0] _16748;
    wire [63:0] _16749;
    wire [62:0] _16750;
    wire [63:0] _16752;
    wire _16753;
    wire _16754;
    wire _16742;
    wire [63:0] _16739;
    wire [63:0] _16740;
    wire [62:0] _16741;
    wire [63:0] _16743;
    wire _16744;
    wire _16745;
    wire _16733;
    wire [63:0] _16730;
    wire [63:0] _16731;
    wire [62:0] _16732;
    wire [63:0] _16734;
    wire _16735;
    wire _16736;
    wire _16724;
    wire [63:0] _16721;
    wire [63:0] _16722;
    wire [62:0] _16723;
    wire [63:0] _16725;
    wire _16726;
    wire _16727;
    wire _16715;
    wire [63:0] _16712;
    wire [63:0] _16713;
    wire [62:0] _16714;
    wire [63:0] _16716;
    wire _16717;
    wire _16718;
    wire _16706;
    wire [63:0] _16703;
    wire [63:0] _16704;
    wire [62:0] _16705;
    wire [63:0] _16707;
    wire _16708;
    wire _16709;
    wire _16697;
    wire [63:0] _16694;
    wire [63:0] _16695;
    wire [62:0] _16696;
    wire [63:0] _16698;
    wire _16699;
    wire _16700;
    wire _16688;
    wire [63:0] _16685;
    wire [63:0] _16686;
    wire [62:0] _16687;
    wire [63:0] _16689;
    wire _16690;
    wire _16691;
    wire _16679;
    wire [63:0] _16676;
    wire [63:0] _16677;
    wire [62:0] _16678;
    wire [63:0] _16680;
    wire _16681;
    wire _16682;
    wire _16670;
    wire [63:0] _16667;
    wire [63:0] _16668;
    wire [62:0] _16669;
    wire [63:0] _16671;
    wire _16672;
    wire _16673;
    wire _16661;
    wire [63:0] _16658;
    wire [63:0] _16659;
    wire [62:0] _16660;
    wire [63:0] _16662;
    wire _16663;
    wire _16664;
    wire _16652;
    wire [63:0] _16649;
    wire [63:0] _16650;
    wire [62:0] _16651;
    wire [63:0] _16653;
    wire _16654;
    wire _16655;
    wire _16643;
    wire [63:0] _16640;
    wire [63:0] _16641;
    wire [62:0] _16642;
    wire [63:0] _16644;
    wire _16645;
    wire _16646;
    wire _16634;
    wire [63:0] _16631;
    wire [63:0] _16632;
    wire [62:0] _16633;
    wire [63:0] _16635;
    wire _16636;
    wire _16637;
    wire _16625;
    wire [63:0] _16622;
    wire [63:0] _16623;
    wire [62:0] _16624;
    wire [63:0] _16626;
    wire _16627;
    wire _16628;
    wire _16616;
    wire [63:0] _16613;
    wire [63:0] _16614;
    wire [62:0] _16615;
    wire [63:0] _16617;
    wire _16618;
    wire _16619;
    wire _16607;
    wire [63:0] _16604;
    wire [63:0] _16605;
    wire [62:0] _16606;
    wire [63:0] _16608;
    wire _16609;
    wire _16610;
    wire _16598;
    wire [63:0] _16595;
    wire [63:0] _16596;
    wire [62:0] _16597;
    wire [63:0] _16599;
    wire _16600;
    wire _16601;
    wire _16589;
    wire [63:0] _16586;
    wire [63:0] _16587;
    wire [62:0] _16588;
    wire [63:0] _16590;
    wire _16591;
    wire _16592;
    wire _16580;
    wire [63:0] _16577;
    wire [63:0] _16578;
    wire [62:0] _16579;
    wire [63:0] _16581;
    wire _16582;
    wire _16583;
    wire _16571;
    wire [63:0] _16568;
    wire [63:0] _16569;
    wire [62:0] _16570;
    wire [63:0] _16572;
    wire _16573;
    wire _16574;
    wire _16562;
    wire [63:0] _16559;
    wire [63:0] _16560;
    wire [62:0] _16561;
    wire [63:0] _16563;
    wire _16564;
    wire _16565;
    wire _16553;
    wire [63:0] _16550;
    wire [63:0] _16551;
    wire [62:0] _16552;
    wire [63:0] _16554;
    wire _16555;
    wire _16556;
    wire _16544;
    wire [63:0] _16541;
    wire [63:0] _16542;
    wire [62:0] _16543;
    wire [63:0] _16545;
    wire _16546;
    wire _16547;
    wire _16535;
    wire [63:0] _16532;
    wire [63:0] _16533;
    wire [62:0] _16534;
    wire [63:0] _16536;
    wire _16537;
    wire _16538;
    wire _16526;
    wire [63:0] _16523;
    wire [63:0] _16524;
    wire [62:0] _16525;
    wire [63:0] _16527;
    wire _16528;
    wire _16529;
    wire _16517;
    wire [63:0] _16514;
    wire [63:0] _16515;
    wire [62:0] _16516;
    wire [63:0] _16518;
    wire _16519;
    wire _16520;
    wire _16508;
    wire [63:0] _16505;
    wire [63:0] _16506;
    wire [62:0] _16507;
    wire [63:0] _16509;
    wire _16510;
    wire _16511;
    wire _16499;
    wire [63:0] _16496;
    wire [63:0] _16497;
    wire [62:0] _16498;
    wire [63:0] _16500;
    wire _16501;
    wire _16502;
    wire _16490;
    wire [63:0] _16487;
    wire [63:0] _16488;
    wire [62:0] _16489;
    wire [63:0] _16491;
    wire _16492;
    wire _16493;
    wire _16481;
    wire [63:0] _16478;
    wire [63:0] _16479;
    wire [62:0] _16480;
    wire [63:0] _16482;
    wire _16483;
    wire _16484;
    wire _16472;
    wire [63:0] _16469;
    wire [63:0] _16470;
    wire [62:0] _16471;
    wire [63:0] _16473;
    wire _16474;
    wire _16475;
    wire _16463;
    wire [63:0] _16460;
    wire [63:0] _16461;
    wire [62:0] _16462;
    wire [63:0] _16464;
    wire _16465;
    wire _16466;
    wire _16454;
    wire [63:0] _16451;
    wire [63:0] _16452;
    wire [62:0] _16453;
    wire [63:0] _16455;
    wire _16456;
    wire _16457;
    wire _16445;
    wire [63:0] _16442;
    wire [63:0] _16443;
    wire [62:0] _16444;
    wire [63:0] _16446;
    wire _16447;
    wire _16448;
    wire _16436;
    wire [63:0] _16433;
    wire [63:0] _16434;
    wire [62:0] _16435;
    wire [63:0] _16437;
    wire _16438;
    wire _16439;
    wire _16427;
    wire [63:0] _16424;
    wire [63:0] _16425;
    wire [62:0] _16426;
    wire [63:0] _16428;
    wire _16429;
    wire _16430;
    wire _16418;
    wire [63:0] _16415;
    wire [63:0] _16416;
    wire [62:0] _16417;
    wire [63:0] _16419;
    wire _16420;
    wire _16421;
    wire _16409;
    wire [63:0] _16406;
    wire [63:0] _16407;
    wire [62:0] _16408;
    wire [63:0] _16410;
    wire _16411;
    wire _16412;
    wire _16400;
    wire [63:0] _16397;
    wire [63:0] _16398;
    wire [62:0] _16399;
    wire [63:0] _16401;
    wire _16402;
    wire _16403;
    wire _16391;
    wire [63:0] _16388;
    wire [63:0] _16389;
    wire [62:0] _16390;
    wire [63:0] _16392;
    wire _16393;
    wire _16394;
    wire _16382;
    wire [63:0] _16379;
    wire [63:0] _16380;
    wire [62:0] _16381;
    wire [63:0] _16383;
    wire _16384;
    wire _16385;
    wire _16373;
    wire [63:0] _16370;
    wire [63:0] _16371;
    wire [62:0] _16372;
    wire [63:0] _16374;
    wire _16375;
    wire _16376;
    wire _16364;
    wire [63:0] _16361;
    wire [63:0] _16362;
    wire [62:0] _16363;
    wire [63:0] _16365;
    wire _16366;
    wire _16367;
    wire [63:0] _16354;
    wire _16355;
    wire [63:0] _16356;
    wire _16357;
    wire _16358;
    wire [63:0] _16359;
    wire [62:0] _16360;
    wire [63:0] _16368;
    wire [62:0] _16369;
    wire [63:0] _16377;
    wire [62:0] _16378;
    wire [63:0] _16386;
    wire [62:0] _16387;
    wire [63:0] _16395;
    wire [62:0] _16396;
    wire [63:0] _16404;
    wire [62:0] _16405;
    wire [63:0] _16413;
    wire [62:0] _16414;
    wire [63:0] _16422;
    wire [62:0] _16423;
    wire [63:0] _16431;
    wire [62:0] _16432;
    wire [63:0] _16440;
    wire [62:0] _16441;
    wire [63:0] _16449;
    wire [62:0] _16450;
    wire [63:0] _16458;
    wire [62:0] _16459;
    wire [63:0] _16467;
    wire [62:0] _16468;
    wire [63:0] _16476;
    wire [62:0] _16477;
    wire [63:0] _16485;
    wire [62:0] _16486;
    wire [63:0] _16494;
    wire [62:0] _16495;
    wire [63:0] _16503;
    wire [62:0] _16504;
    wire [63:0] _16512;
    wire [62:0] _16513;
    wire [63:0] _16521;
    wire [62:0] _16522;
    wire [63:0] _16530;
    wire [62:0] _16531;
    wire [63:0] _16539;
    wire [62:0] _16540;
    wire [63:0] _16548;
    wire [62:0] _16549;
    wire [63:0] _16557;
    wire [62:0] _16558;
    wire [63:0] _16566;
    wire [62:0] _16567;
    wire [63:0] _16575;
    wire [62:0] _16576;
    wire [63:0] _16584;
    wire [62:0] _16585;
    wire [63:0] _16593;
    wire [62:0] _16594;
    wire [63:0] _16602;
    wire [62:0] _16603;
    wire [63:0] _16611;
    wire [62:0] _16612;
    wire [63:0] _16620;
    wire [62:0] _16621;
    wire [63:0] _16629;
    wire [62:0] _16630;
    wire [63:0] _16638;
    wire [62:0] _16639;
    wire [63:0] _16647;
    wire [62:0] _16648;
    wire [63:0] _16656;
    wire [62:0] _16657;
    wire [63:0] _16665;
    wire [62:0] _16666;
    wire [63:0] _16674;
    wire [62:0] _16675;
    wire [63:0] _16683;
    wire [62:0] _16684;
    wire [63:0] _16692;
    wire [62:0] _16693;
    wire [63:0] _16701;
    wire [62:0] _16702;
    wire [63:0] _16710;
    wire [62:0] _16711;
    wire [63:0] _16719;
    wire [62:0] _16720;
    wire [63:0] _16728;
    wire [62:0] _16729;
    wire [63:0] _16737;
    wire [62:0] _16738;
    wire [63:0] _16746;
    wire [62:0] _16747;
    wire [63:0] _16755;
    wire [62:0] _16756;
    wire [63:0] _16764;
    wire [62:0] _16765;
    wire [63:0] _16773;
    wire [62:0] _16774;
    wire [63:0] _16782;
    wire [62:0] _16783;
    wire [63:0] _16791;
    wire [62:0] _16792;
    wire [63:0] _16800;
    wire [62:0] _16801;
    wire [63:0] _16809;
    wire [62:0] _16810;
    wire [63:0] _16818;
    wire [62:0] _16819;
    wire [63:0] _16827;
    wire [62:0] _16828;
    wire [63:0] _16836;
    wire [62:0] _16837;
    wire [63:0] _16845;
    wire [62:0] _16846;
    wire [63:0] _16854;
    wire [62:0] _16855;
    wire [63:0] _16863;
    wire [62:0] _16864;
    wire [63:0] _16872;
    wire [62:0] _16873;
    wire [63:0] _16881;
    wire [62:0] _16882;
    wire [63:0] _16890;
    wire [62:0] _16891;
    wire [63:0] _16899;
    wire [62:0] _16900;
    wire [63:0] _16908;
    wire [62:0] _16909;
    wire [63:0] _16917;
    wire [62:0] _16918;
    wire [63:0] _16926;
    wire [63:0] _16928;
    wire [127:0] _16929;
    wire [63:0] _16930;
    wire [63:0] _17512;
    wire _16340;
    wire [63:0] _16337;
    wire [63:0] _16338;
    wire [62:0] _16339;
    wire [63:0] _16341;
    wire _16342;
    wire _16343;
    wire _16331;
    wire [63:0] _16328;
    wire [63:0] _16329;
    wire [62:0] _16330;
    wire [63:0] _16332;
    wire _16333;
    wire _16334;
    wire _16322;
    wire [63:0] _16319;
    wire [63:0] _16320;
    wire [62:0] _16321;
    wire [63:0] _16323;
    wire _16324;
    wire _16325;
    wire _16313;
    wire [63:0] _16310;
    wire [63:0] _16311;
    wire [62:0] _16312;
    wire [63:0] _16314;
    wire _16315;
    wire _16316;
    wire _16304;
    wire [63:0] _16301;
    wire [63:0] _16302;
    wire [62:0] _16303;
    wire [63:0] _16305;
    wire _16306;
    wire _16307;
    wire _16295;
    wire [63:0] _16292;
    wire [63:0] _16293;
    wire [62:0] _16294;
    wire [63:0] _16296;
    wire _16297;
    wire _16298;
    wire _16286;
    wire [63:0] _16283;
    wire [63:0] _16284;
    wire [62:0] _16285;
    wire [63:0] _16287;
    wire _16288;
    wire _16289;
    wire _16277;
    wire [63:0] _16274;
    wire [63:0] _16275;
    wire [62:0] _16276;
    wire [63:0] _16278;
    wire _16279;
    wire _16280;
    wire _16268;
    wire [63:0] _16265;
    wire [63:0] _16266;
    wire [62:0] _16267;
    wire [63:0] _16269;
    wire _16270;
    wire _16271;
    wire _16259;
    wire [63:0] _16256;
    wire [63:0] _16257;
    wire [62:0] _16258;
    wire [63:0] _16260;
    wire _16261;
    wire _16262;
    wire _16250;
    wire [63:0] _16247;
    wire [63:0] _16248;
    wire [62:0] _16249;
    wire [63:0] _16251;
    wire _16252;
    wire _16253;
    wire _16241;
    wire [63:0] _16238;
    wire [63:0] _16239;
    wire [62:0] _16240;
    wire [63:0] _16242;
    wire _16243;
    wire _16244;
    wire _16232;
    wire [63:0] _16229;
    wire [63:0] _16230;
    wire [62:0] _16231;
    wire [63:0] _16233;
    wire _16234;
    wire _16235;
    wire _16223;
    wire [63:0] _16220;
    wire [63:0] _16221;
    wire [62:0] _16222;
    wire [63:0] _16224;
    wire _16225;
    wire _16226;
    wire _16214;
    wire [63:0] _16211;
    wire [63:0] _16212;
    wire [62:0] _16213;
    wire [63:0] _16215;
    wire _16216;
    wire _16217;
    wire _16205;
    wire [63:0] _16202;
    wire [63:0] _16203;
    wire [62:0] _16204;
    wire [63:0] _16206;
    wire _16207;
    wire _16208;
    wire _16196;
    wire [63:0] _16193;
    wire [63:0] _16194;
    wire [62:0] _16195;
    wire [63:0] _16197;
    wire _16198;
    wire _16199;
    wire _16187;
    wire [63:0] _16184;
    wire [63:0] _16185;
    wire [62:0] _16186;
    wire [63:0] _16188;
    wire _16189;
    wire _16190;
    wire _16178;
    wire [63:0] _16175;
    wire [63:0] _16176;
    wire [62:0] _16177;
    wire [63:0] _16179;
    wire _16180;
    wire _16181;
    wire _16169;
    wire [63:0] _16166;
    wire [63:0] _16167;
    wire [62:0] _16168;
    wire [63:0] _16170;
    wire _16171;
    wire _16172;
    wire _16160;
    wire [63:0] _16157;
    wire [63:0] _16158;
    wire [62:0] _16159;
    wire [63:0] _16161;
    wire _16162;
    wire _16163;
    wire _16151;
    wire [63:0] _16148;
    wire [63:0] _16149;
    wire [62:0] _16150;
    wire [63:0] _16152;
    wire _16153;
    wire _16154;
    wire _16142;
    wire [63:0] _16139;
    wire [63:0] _16140;
    wire [62:0] _16141;
    wire [63:0] _16143;
    wire _16144;
    wire _16145;
    wire _16133;
    wire [63:0] _16130;
    wire [63:0] _16131;
    wire [62:0] _16132;
    wire [63:0] _16134;
    wire _16135;
    wire _16136;
    wire _16124;
    wire [63:0] _16121;
    wire [63:0] _16122;
    wire [62:0] _16123;
    wire [63:0] _16125;
    wire _16126;
    wire _16127;
    wire _16115;
    wire [63:0] _16112;
    wire [63:0] _16113;
    wire [62:0] _16114;
    wire [63:0] _16116;
    wire _16117;
    wire _16118;
    wire _16106;
    wire [63:0] _16103;
    wire [63:0] _16104;
    wire [62:0] _16105;
    wire [63:0] _16107;
    wire _16108;
    wire _16109;
    wire _16097;
    wire [63:0] _16094;
    wire [63:0] _16095;
    wire [62:0] _16096;
    wire [63:0] _16098;
    wire _16099;
    wire _16100;
    wire _16088;
    wire [63:0] _16085;
    wire [63:0] _16086;
    wire [62:0] _16087;
    wire [63:0] _16089;
    wire _16090;
    wire _16091;
    wire _16079;
    wire [63:0] _16076;
    wire [63:0] _16077;
    wire [62:0] _16078;
    wire [63:0] _16080;
    wire _16081;
    wire _16082;
    wire _16070;
    wire [63:0] _16067;
    wire [63:0] _16068;
    wire [62:0] _16069;
    wire [63:0] _16071;
    wire _16072;
    wire _16073;
    wire _16061;
    wire [63:0] _16058;
    wire [63:0] _16059;
    wire [62:0] _16060;
    wire [63:0] _16062;
    wire _16063;
    wire _16064;
    wire _16052;
    wire [63:0] _16049;
    wire [63:0] _16050;
    wire [62:0] _16051;
    wire [63:0] _16053;
    wire _16054;
    wire _16055;
    wire _16043;
    wire [63:0] _16040;
    wire [63:0] _16041;
    wire [62:0] _16042;
    wire [63:0] _16044;
    wire _16045;
    wire _16046;
    wire _16034;
    wire [63:0] _16031;
    wire [63:0] _16032;
    wire [62:0] _16033;
    wire [63:0] _16035;
    wire _16036;
    wire _16037;
    wire _16025;
    wire [63:0] _16022;
    wire [63:0] _16023;
    wire [62:0] _16024;
    wire [63:0] _16026;
    wire _16027;
    wire _16028;
    wire _16016;
    wire [63:0] _16013;
    wire [63:0] _16014;
    wire [62:0] _16015;
    wire [63:0] _16017;
    wire _16018;
    wire _16019;
    wire _16007;
    wire [63:0] _16004;
    wire [63:0] _16005;
    wire [62:0] _16006;
    wire [63:0] _16008;
    wire _16009;
    wire _16010;
    wire _15998;
    wire [63:0] _15995;
    wire [63:0] _15996;
    wire [62:0] _15997;
    wire [63:0] _15999;
    wire _16000;
    wire _16001;
    wire _15989;
    wire [63:0] _15986;
    wire [63:0] _15987;
    wire [62:0] _15988;
    wire [63:0] _15990;
    wire _15991;
    wire _15992;
    wire _15980;
    wire [63:0] _15977;
    wire [63:0] _15978;
    wire [62:0] _15979;
    wire [63:0] _15981;
    wire _15982;
    wire _15983;
    wire _15971;
    wire [63:0] _15968;
    wire [63:0] _15969;
    wire [62:0] _15970;
    wire [63:0] _15972;
    wire _15973;
    wire _15974;
    wire _15962;
    wire [63:0] _15959;
    wire [63:0] _15960;
    wire [62:0] _15961;
    wire [63:0] _15963;
    wire _15964;
    wire _15965;
    wire _15953;
    wire [63:0] _15950;
    wire [63:0] _15951;
    wire [62:0] _15952;
    wire [63:0] _15954;
    wire _15955;
    wire _15956;
    wire _15944;
    wire [63:0] _15941;
    wire [63:0] _15942;
    wire [62:0] _15943;
    wire [63:0] _15945;
    wire _15946;
    wire _15947;
    wire _15935;
    wire [63:0] _15932;
    wire [63:0] _15933;
    wire [62:0] _15934;
    wire [63:0] _15936;
    wire _15937;
    wire _15938;
    wire _15926;
    wire [63:0] _15923;
    wire [63:0] _15924;
    wire [62:0] _15925;
    wire [63:0] _15927;
    wire _15928;
    wire _15929;
    wire _15917;
    wire [63:0] _15914;
    wire [63:0] _15915;
    wire [62:0] _15916;
    wire [63:0] _15918;
    wire _15919;
    wire _15920;
    wire _15908;
    wire [63:0] _15905;
    wire [63:0] _15906;
    wire [62:0] _15907;
    wire [63:0] _15909;
    wire _15910;
    wire _15911;
    wire _15899;
    wire [63:0] _15896;
    wire [63:0] _15897;
    wire [62:0] _15898;
    wire [63:0] _15900;
    wire _15901;
    wire _15902;
    wire _15890;
    wire [63:0] _15887;
    wire [63:0] _15888;
    wire [62:0] _15889;
    wire [63:0] _15891;
    wire _15892;
    wire _15893;
    wire _15881;
    wire [63:0] _15878;
    wire [63:0] _15879;
    wire [62:0] _15880;
    wire [63:0] _15882;
    wire _15883;
    wire _15884;
    wire _15872;
    wire [63:0] _15869;
    wire [63:0] _15870;
    wire [62:0] _15871;
    wire [63:0] _15873;
    wire _15874;
    wire _15875;
    wire _15863;
    wire [63:0] _15860;
    wire [63:0] _15861;
    wire [62:0] _15862;
    wire [63:0] _15864;
    wire _15865;
    wire _15866;
    wire _15854;
    wire [63:0] _15851;
    wire [63:0] _15852;
    wire [62:0] _15853;
    wire [63:0] _15855;
    wire _15856;
    wire _15857;
    wire _15845;
    wire [63:0] _15842;
    wire [63:0] _15843;
    wire [62:0] _15844;
    wire [63:0] _15846;
    wire _15847;
    wire _15848;
    wire _15836;
    wire [63:0] _15833;
    wire [63:0] _15834;
    wire [62:0] _15835;
    wire [63:0] _15837;
    wire _15838;
    wire _15839;
    wire _15827;
    wire [63:0] _15824;
    wire [63:0] _15825;
    wire [62:0] _15826;
    wire [63:0] _15828;
    wire _15829;
    wire _15830;
    wire _15818;
    wire [63:0] _15815;
    wire [63:0] _15816;
    wire [62:0] _15817;
    wire [63:0] _15819;
    wire _15820;
    wire _15821;
    wire _15809;
    wire [63:0] _15806;
    wire [63:0] _15807;
    wire [62:0] _15808;
    wire [63:0] _15810;
    wire _15811;
    wire _15812;
    wire _15800;
    wire [63:0] _15797;
    wire [63:0] _15798;
    wire [62:0] _15799;
    wire [63:0] _15801;
    wire _15802;
    wire _15803;
    wire _15791;
    wire [63:0] _15788;
    wire [63:0] _15789;
    wire [62:0] _15790;
    wire [63:0] _15792;
    wire _15793;
    wire _15794;
    wire _15782;
    wire [63:0] _15779;
    wire [63:0] _15780;
    wire [62:0] _15781;
    wire [63:0] _15783;
    wire _15784;
    wire _15785;
    wire [63:0] _15774;
    wire [63:0] _15770;
    wire [63:0] _15771;
    wire _15772;
    wire [63:0] _15773;
    wire _15775;
    wire _15776;
    wire [63:0] _15777;
    wire [62:0] _15778;
    wire [63:0] _15786;
    wire [62:0] _15787;
    wire [63:0] _15795;
    wire [62:0] _15796;
    wire [63:0] _15804;
    wire [62:0] _15805;
    wire [63:0] _15813;
    wire [62:0] _15814;
    wire [63:0] _15822;
    wire [62:0] _15823;
    wire [63:0] _15831;
    wire [62:0] _15832;
    wire [63:0] _15840;
    wire [62:0] _15841;
    wire [63:0] _15849;
    wire [62:0] _15850;
    wire [63:0] _15858;
    wire [62:0] _15859;
    wire [63:0] _15867;
    wire [62:0] _15868;
    wire [63:0] _15876;
    wire [62:0] _15877;
    wire [63:0] _15885;
    wire [62:0] _15886;
    wire [63:0] _15894;
    wire [62:0] _15895;
    wire [63:0] _15903;
    wire [62:0] _15904;
    wire [63:0] _15912;
    wire [62:0] _15913;
    wire [63:0] _15921;
    wire [62:0] _15922;
    wire [63:0] _15930;
    wire [62:0] _15931;
    wire [63:0] _15939;
    wire [62:0] _15940;
    wire [63:0] _15948;
    wire [62:0] _15949;
    wire [63:0] _15957;
    wire [62:0] _15958;
    wire [63:0] _15966;
    wire [62:0] _15967;
    wire [63:0] _15975;
    wire [62:0] _15976;
    wire [63:0] _15984;
    wire [62:0] _15985;
    wire [63:0] _15993;
    wire [62:0] _15994;
    wire [63:0] _16002;
    wire [62:0] _16003;
    wire [63:0] _16011;
    wire [62:0] _16012;
    wire [63:0] _16020;
    wire [62:0] _16021;
    wire [63:0] _16029;
    wire [62:0] _16030;
    wire [63:0] _16038;
    wire [62:0] _16039;
    wire [63:0] _16047;
    wire [62:0] _16048;
    wire [63:0] _16056;
    wire [62:0] _16057;
    wire [63:0] _16065;
    wire [62:0] _16066;
    wire [63:0] _16074;
    wire [62:0] _16075;
    wire [63:0] _16083;
    wire [62:0] _16084;
    wire [63:0] _16092;
    wire [62:0] _16093;
    wire [63:0] _16101;
    wire [62:0] _16102;
    wire [63:0] _16110;
    wire [62:0] _16111;
    wire [63:0] _16119;
    wire [62:0] _16120;
    wire [63:0] _16128;
    wire [62:0] _16129;
    wire [63:0] _16137;
    wire [62:0] _16138;
    wire [63:0] _16146;
    wire [62:0] _16147;
    wire [63:0] _16155;
    wire [62:0] _16156;
    wire [63:0] _16164;
    wire [62:0] _16165;
    wire [63:0] _16173;
    wire [62:0] _16174;
    wire [63:0] _16182;
    wire [62:0] _16183;
    wire [63:0] _16191;
    wire [62:0] _16192;
    wire [63:0] _16200;
    wire [62:0] _16201;
    wire [63:0] _16209;
    wire [62:0] _16210;
    wire [63:0] _16218;
    wire [62:0] _16219;
    wire [63:0] _16227;
    wire [62:0] _16228;
    wire [63:0] _16236;
    wire [62:0] _16237;
    wire [63:0] _16245;
    wire [62:0] _16246;
    wire [63:0] _16254;
    wire [62:0] _16255;
    wire [63:0] _16263;
    wire [62:0] _16264;
    wire [63:0] _16272;
    wire [62:0] _16273;
    wire [63:0] _16281;
    wire [62:0] _16282;
    wire [63:0] _16290;
    wire [62:0] _16291;
    wire [63:0] _16299;
    wire [62:0] _16300;
    wire [63:0] _16308;
    wire [62:0] _16309;
    wire [63:0] _16317;
    wire [62:0] _16318;
    wire [63:0] _16326;
    wire [62:0] _16327;
    wire [63:0] _16335;
    wire [62:0] _16336;
    wire [63:0] _16344;
    wire [127:0] _16345;
    wire [63:0] _16346;
    wire [63:0] _15767;
    wire _16347;
    wire [63:0] _16348;
    wire [63:0] _15764;
    wire _15765;
    wire [63:0] _15766;
    wire _16349;
    wire _16350;
    wire [63:0] _17513;
    wire _15754;
    wire [63:0] _15751;
    wire [63:0] _15752;
    wire [62:0] _15753;
    wire [63:0] _15755;
    wire _15756;
    wire _15757;
    wire _15745;
    wire [63:0] _15742;
    wire [63:0] _15743;
    wire [62:0] _15744;
    wire [63:0] _15746;
    wire _15747;
    wire _15748;
    wire _15736;
    wire [63:0] _15733;
    wire [63:0] _15734;
    wire [62:0] _15735;
    wire [63:0] _15737;
    wire _15738;
    wire _15739;
    wire _15727;
    wire [63:0] _15724;
    wire [63:0] _15725;
    wire [62:0] _15726;
    wire [63:0] _15728;
    wire _15729;
    wire _15730;
    wire _15718;
    wire [63:0] _15715;
    wire [63:0] _15716;
    wire [62:0] _15717;
    wire [63:0] _15719;
    wire _15720;
    wire _15721;
    wire _15709;
    wire [63:0] _15706;
    wire [63:0] _15707;
    wire [62:0] _15708;
    wire [63:0] _15710;
    wire _15711;
    wire _15712;
    wire _15700;
    wire [63:0] _15697;
    wire [63:0] _15698;
    wire [62:0] _15699;
    wire [63:0] _15701;
    wire _15702;
    wire _15703;
    wire _15691;
    wire [63:0] _15688;
    wire [63:0] _15689;
    wire [62:0] _15690;
    wire [63:0] _15692;
    wire _15693;
    wire _15694;
    wire _15682;
    wire [63:0] _15679;
    wire [63:0] _15680;
    wire [62:0] _15681;
    wire [63:0] _15683;
    wire _15684;
    wire _15685;
    wire _15673;
    wire [63:0] _15670;
    wire [63:0] _15671;
    wire [62:0] _15672;
    wire [63:0] _15674;
    wire _15675;
    wire _15676;
    wire _15664;
    wire [63:0] _15661;
    wire [63:0] _15662;
    wire [62:0] _15663;
    wire [63:0] _15665;
    wire _15666;
    wire _15667;
    wire _15655;
    wire [63:0] _15652;
    wire [63:0] _15653;
    wire [62:0] _15654;
    wire [63:0] _15656;
    wire _15657;
    wire _15658;
    wire _15646;
    wire [63:0] _15643;
    wire [63:0] _15644;
    wire [62:0] _15645;
    wire [63:0] _15647;
    wire _15648;
    wire _15649;
    wire _15637;
    wire [63:0] _15634;
    wire [63:0] _15635;
    wire [62:0] _15636;
    wire [63:0] _15638;
    wire _15639;
    wire _15640;
    wire _15628;
    wire [63:0] _15625;
    wire [63:0] _15626;
    wire [62:0] _15627;
    wire [63:0] _15629;
    wire _15630;
    wire _15631;
    wire _15619;
    wire [63:0] _15616;
    wire [63:0] _15617;
    wire [62:0] _15618;
    wire [63:0] _15620;
    wire _15621;
    wire _15622;
    wire _15610;
    wire [63:0] _15607;
    wire [63:0] _15608;
    wire [62:0] _15609;
    wire [63:0] _15611;
    wire _15612;
    wire _15613;
    wire _15601;
    wire [63:0] _15598;
    wire [63:0] _15599;
    wire [62:0] _15600;
    wire [63:0] _15602;
    wire _15603;
    wire _15604;
    wire _15592;
    wire [63:0] _15589;
    wire [63:0] _15590;
    wire [62:0] _15591;
    wire [63:0] _15593;
    wire _15594;
    wire _15595;
    wire _15583;
    wire [63:0] _15580;
    wire [63:0] _15581;
    wire [62:0] _15582;
    wire [63:0] _15584;
    wire _15585;
    wire _15586;
    wire _15574;
    wire [63:0] _15571;
    wire [63:0] _15572;
    wire [62:0] _15573;
    wire [63:0] _15575;
    wire _15576;
    wire _15577;
    wire _15565;
    wire [63:0] _15562;
    wire [63:0] _15563;
    wire [62:0] _15564;
    wire [63:0] _15566;
    wire _15567;
    wire _15568;
    wire _15556;
    wire [63:0] _15553;
    wire [63:0] _15554;
    wire [62:0] _15555;
    wire [63:0] _15557;
    wire _15558;
    wire _15559;
    wire _15547;
    wire [63:0] _15544;
    wire [63:0] _15545;
    wire [62:0] _15546;
    wire [63:0] _15548;
    wire _15549;
    wire _15550;
    wire _15538;
    wire [63:0] _15535;
    wire [63:0] _15536;
    wire [62:0] _15537;
    wire [63:0] _15539;
    wire _15540;
    wire _15541;
    wire _15529;
    wire [63:0] _15526;
    wire [63:0] _15527;
    wire [62:0] _15528;
    wire [63:0] _15530;
    wire _15531;
    wire _15532;
    wire _15520;
    wire [63:0] _15517;
    wire [63:0] _15518;
    wire [62:0] _15519;
    wire [63:0] _15521;
    wire _15522;
    wire _15523;
    wire _15511;
    wire [63:0] _15508;
    wire [63:0] _15509;
    wire [62:0] _15510;
    wire [63:0] _15512;
    wire _15513;
    wire _15514;
    wire _15502;
    wire [63:0] _15499;
    wire [63:0] _15500;
    wire [62:0] _15501;
    wire [63:0] _15503;
    wire _15504;
    wire _15505;
    wire _15493;
    wire [63:0] _15490;
    wire [63:0] _15491;
    wire [62:0] _15492;
    wire [63:0] _15494;
    wire _15495;
    wire _15496;
    wire _15484;
    wire [63:0] _15481;
    wire [63:0] _15482;
    wire [62:0] _15483;
    wire [63:0] _15485;
    wire _15486;
    wire _15487;
    wire _15475;
    wire [63:0] _15472;
    wire [63:0] _15473;
    wire [62:0] _15474;
    wire [63:0] _15476;
    wire _15477;
    wire _15478;
    wire _15466;
    wire [63:0] _15463;
    wire [63:0] _15464;
    wire [62:0] _15465;
    wire [63:0] _15467;
    wire _15468;
    wire _15469;
    wire _15457;
    wire [63:0] _15454;
    wire [63:0] _15455;
    wire [62:0] _15456;
    wire [63:0] _15458;
    wire _15459;
    wire _15460;
    wire _15448;
    wire [63:0] _15445;
    wire [63:0] _15446;
    wire [62:0] _15447;
    wire [63:0] _15449;
    wire _15450;
    wire _15451;
    wire _15439;
    wire [63:0] _15436;
    wire [63:0] _15437;
    wire [62:0] _15438;
    wire [63:0] _15440;
    wire _15441;
    wire _15442;
    wire _15430;
    wire [63:0] _15427;
    wire [63:0] _15428;
    wire [62:0] _15429;
    wire [63:0] _15431;
    wire _15432;
    wire _15433;
    wire _15421;
    wire [63:0] _15418;
    wire [63:0] _15419;
    wire [62:0] _15420;
    wire [63:0] _15422;
    wire _15423;
    wire _15424;
    wire _15412;
    wire [63:0] _15409;
    wire [63:0] _15410;
    wire [62:0] _15411;
    wire [63:0] _15413;
    wire _15414;
    wire _15415;
    wire _15403;
    wire [63:0] _15400;
    wire [63:0] _15401;
    wire [62:0] _15402;
    wire [63:0] _15404;
    wire _15405;
    wire _15406;
    wire _15394;
    wire [63:0] _15391;
    wire [63:0] _15392;
    wire [62:0] _15393;
    wire [63:0] _15395;
    wire _15396;
    wire _15397;
    wire _15385;
    wire [63:0] _15382;
    wire [63:0] _15383;
    wire [62:0] _15384;
    wire [63:0] _15386;
    wire _15387;
    wire _15388;
    wire _15376;
    wire [63:0] _15373;
    wire [63:0] _15374;
    wire [62:0] _15375;
    wire [63:0] _15377;
    wire _15378;
    wire _15379;
    wire _15367;
    wire [63:0] _15364;
    wire [63:0] _15365;
    wire [62:0] _15366;
    wire [63:0] _15368;
    wire _15369;
    wire _15370;
    wire _15358;
    wire [63:0] _15355;
    wire [63:0] _15356;
    wire [62:0] _15357;
    wire [63:0] _15359;
    wire _15360;
    wire _15361;
    wire _15349;
    wire [63:0] _15346;
    wire [63:0] _15347;
    wire [62:0] _15348;
    wire [63:0] _15350;
    wire _15351;
    wire _15352;
    wire _15340;
    wire [63:0] _15337;
    wire [63:0] _15338;
    wire [62:0] _15339;
    wire [63:0] _15341;
    wire _15342;
    wire _15343;
    wire _15331;
    wire [63:0] _15328;
    wire [63:0] _15329;
    wire [62:0] _15330;
    wire [63:0] _15332;
    wire _15333;
    wire _15334;
    wire _15322;
    wire [63:0] _15319;
    wire [63:0] _15320;
    wire [62:0] _15321;
    wire [63:0] _15323;
    wire _15324;
    wire _15325;
    wire _15313;
    wire [63:0] _15310;
    wire [63:0] _15311;
    wire [62:0] _15312;
    wire [63:0] _15314;
    wire _15315;
    wire _15316;
    wire _15304;
    wire [63:0] _15301;
    wire [63:0] _15302;
    wire [62:0] _15303;
    wire [63:0] _15305;
    wire _15306;
    wire _15307;
    wire _15295;
    wire [63:0] _15292;
    wire [63:0] _15293;
    wire [62:0] _15294;
    wire [63:0] _15296;
    wire _15297;
    wire _15298;
    wire _15286;
    wire [63:0] _15283;
    wire [63:0] _15284;
    wire [62:0] _15285;
    wire [63:0] _15287;
    wire _15288;
    wire _15289;
    wire _15277;
    wire [63:0] _15274;
    wire [63:0] _15275;
    wire [62:0] _15276;
    wire [63:0] _15278;
    wire _15279;
    wire _15280;
    wire _15268;
    wire [63:0] _15265;
    wire [63:0] _15266;
    wire [62:0] _15267;
    wire [63:0] _15269;
    wire _15270;
    wire _15271;
    wire _15259;
    wire [63:0] _15256;
    wire [63:0] _15257;
    wire [62:0] _15258;
    wire [63:0] _15260;
    wire _15261;
    wire _15262;
    wire _15250;
    wire [63:0] _15247;
    wire [63:0] _15248;
    wire [62:0] _15249;
    wire [63:0] _15251;
    wire _15252;
    wire _15253;
    wire _15241;
    wire [63:0] _15238;
    wire [63:0] _15239;
    wire [62:0] _15240;
    wire [63:0] _15242;
    wire _15243;
    wire _15244;
    wire _15232;
    wire [63:0] _15229;
    wire [63:0] _15230;
    wire [62:0] _15231;
    wire [63:0] _15233;
    wire _15234;
    wire _15235;
    wire _15223;
    wire [63:0] _15220;
    wire [63:0] _15221;
    wire [62:0] _15222;
    wire [63:0] _15224;
    wire _15225;
    wire _15226;
    wire _15214;
    wire [63:0] _15211;
    wire [63:0] _15212;
    wire [62:0] _15213;
    wire [63:0] _15215;
    wire _15216;
    wire _15217;
    wire _15205;
    wire [63:0] _15202;
    wire [63:0] _15203;
    wire [62:0] _15204;
    wire [63:0] _15206;
    wire _15207;
    wire _15208;
    wire _15196;
    wire [63:0] _15193;
    wire [63:0] _15194;
    wire [62:0] _15195;
    wire [63:0] _15197;
    wire _15198;
    wire _15199;
    wire [63:0] _15183;
    wire [127:0] _15184;
    wire [63:0] _15185;
    wire _15186;
    wire [63:0] _15187;
    wire _15189;
    wire _15190;
    wire [63:0] _15191;
    wire [62:0] _15192;
    wire [63:0] _15200;
    wire [62:0] _15201;
    wire [63:0] _15209;
    wire [62:0] _15210;
    wire [63:0] _15218;
    wire [62:0] _15219;
    wire [63:0] _15227;
    wire [62:0] _15228;
    wire [63:0] _15236;
    wire [62:0] _15237;
    wire [63:0] _15245;
    wire [62:0] _15246;
    wire [63:0] _15254;
    wire [62:0] _15255;
    wire [63:0] _15263;
    wire [62:0] _15264;
    wire [63:0] _15272;
    wire [62:0] _15273;
    wire [63:0] _15281;
    wire [62:0] _15282;
    wire [63:0] _15290;
    wire [62:0] _15291;
    wire [63:0] _15299;
    wire [62:0] _15300;
    wire [63:0] _15308;
    wire [62:0] _15309;
    wire [63:0] _15317;
    wire [62:0] _15318;
    wire [63:0] _15326;
    wire [62:0] _15327;
    wire [63:0] _15335;
    wire [62:0] _15336;
    wire [63:0] _15344;
    wire [62:0] _15345;
    wire [63:0] _15353;
    wire [62:0] _15354;
    wire [63:0] _15362;
    wire [62:0] _15363;
    wire [63:0] _15371;
    wire [62:0] _15372;
    wire [63:0] _15380;
    wire [62:0] _15381;
    wire [63:0] _15389;
    wire [62:0] _15390;
    wire [63:0] _15398;
    wire [62:0] _15399;
    wire [63:0] _15407;
    wire [62:0] _15408;
    wire [63:0] _15416;
    wire [62:0] _15417;
    wire [63:0] _15425;
    wire [62:0] _15426;
    wire [63:0] _15434;
    wire [62:0] _15435;
    wire [63:0] _15443;
    wire [62:0] _15444;
    wire [63:0] _15452;
    wire [62:0] _15453;
    wire [63:0] _15461;
    wire [62:0] _15462;
    wire [63:0] _15470;
    wire [62:0] _15471;
    wire [63:0] _15479;
    wire [62:0] _15480;
    wire [63:0] _15488;
    wire [62:0] _15489;
    wire [63:0] _15497;
    wire [62:0] _15498;
    wire [63:0] _15506;
    wire [62:0] _15507;
    wire [63:0] _15515;
    wire [62:0] _15516;
    wire [63:0] _15524;
    wire [62:0] _15525;
    wire [63:0] _15533;
    wire [62:0] _15534;
    wire [63:0] _15542;
    wire [62:0] _15543;
    wire [63:0] _15551;
    wire [62:0] _15552;
    wire [63:0] _15560;
    wire [62:0] _15561;
    wire [63:0] _15569;
    wire [62:0] _15570;
    wire [63:0] _15578;
    wire [62:0] _15579;
    wire [63:0] _15587;
    wire [62:0] _15588;
    wire [63:0] _15596;
    wire [62:0] _15597;
    wire [63:0] _15605;
    wire [62:0] _15606;
    wire [63:0] _15614;
    wire [62:0] _15615;
    wire [63:0] _15623;
    wire [62:0] _15624;
    wire [63:0] _15632;
    wire [62:0] _15633;
    wire [63:0] _15641;
    wire [62:0] _15642;
    wire [63:0] _15650;
    wire [62:0] _15651;
    wire [63:0] _15659;
    wire [62:0] _15660;
    wire [63:0] _15668;
    wire [62:0] _15669;
    wire [63:0] _15677;
    wire [62:0] _15678;
    wire [63:0] _15686;
    wire [62:0] _15687;
    wire [63:0] _15695;
    wire [62:0] _15696;
    wire [63:0] _15704;
    wire [62:0] _15705;
    wire [63:0] _15713;
    wire [62:0] _15714;
    wire [63:0] _15722;
    wire [62:0] _15723;
    wire [63:0] _15731;
    wire [62:0] _15732;
    wire [63:0] _15740;
    wire [62:0] _15741;
    wire [63:0] _15749;
    wire [62:0] _15750;
    wire [63:0] _15758;
    wire [127:0] _15759;
    wire [63:0] _15760;
    wire _15171;
    wire [63:0] _15168;
    wire [63:0] _15169;
    wire [62:0] _15170;
    wire [63:0] _15172;
    wire _15173;
    wire _15174;
    wire _15162;
    wire [63:0] _15159;
    wire [63:0] _15160;
    wire [62:0] _15161;
    wire [63:0] _15163;
    wire _15164;
    wire _15165;
    wire _15153;
    wire [63:0] _15150;
    wire [63:0] _15151;
    wire [62:0] _15152;
    wire [63:0] _15154;
    wire _15155;
    wire _15156;
    wire _15144;
    wire [63:0] _15141;
    wire [63:0] _15142;
    wire [62:0] _15143;
    wire [63:0] _15145;
    wire _15146;
    wire _15147;
    wire _15135;
    wire [63:0] _15132;
    wire [63:0] _15133;
    wire [62:0] _15134;
    wire [63:0] _15136;
    wire _15137;
    wire _15138;
    wire _15126;
    wire [63:0] _15123;
    wire [63:0] _15124;
    wire [62:0] _15125;
    wire [63:0] _15127;
    wire _15128;
    wire _15129;
    wire _15117;
    wire [63:0] _15114;
    wire [63:0] _15115;
    wire [62:0] _15116;
    wire [63:0] _15118;
    wire _15119;
    wire _15120;
    wire _15108;
    wire [63:0] _15105;
    wire [63:0] _15106;
    wire [62:0] _15107;
    wire [63:0] _15109;
    wire _15110;
    wire _15111;
    wire _15099;
    wire [63:0] _15096;
    wire [63:0] _15097;
    wire [62:0] _15098;
    wire [63:0] _15100;
    wire _15101;
    wire _15102;
    wire _15090;
    wire [63:0] _15087;
    wire [63:0] _15088;
    wire [62:0] _15089;
    wire [63:0] _15091;
    wire _15092;
    wire _15093;
    wire _15081;
    wire [63:0] _15078;
    wire [63:0] _15079;
    wire [62:0] _15080;
    wire [63:0] _15082;
    wire _15083;
    wire _15084;
    wire _15072;
    wire [63:0] _15069;
    wire [63:0] _15070;
    wire [62:0] _15071;
    wire [63:0] _15073;
    wire _15074;
    wire _15075;
    wire _15063;
    wire [63:0] _15060;
    wire [63:0] _15061;
    wire [62:0] _15062;
    wire [63:0] _15064;
    wire _15065;
    wire _15066;
    wire _15054;
    wire [63:0] _15051;
    wire [63:0] _15052;
    wire [62:0] _15053;
    wire [63:0] _15055;
    wire _15056;
    wire _15057;
    wire _15045;
    wire [63:0] _15042;
    wire [63:0] _15043;
    wire [62:0] _15044;
    wire [63:0] _15046;
    wire _15047;
    wire _15048;
    wire _15036;
    wire [63:0] _15033;
    wire [63:0] _15034;
    wire [62:0] _15035;
    wire [63:0] _15037;
    wire _15038;
    wire _15039;
    wire _15027;
    wire [63:0] _15024;
    wire [63:0] _15025;
    wire [62:0] _15026;
    wire [63:0] _15028;
    wire _15029;
    wire _15030;
    wire _15018;
    wire [63:0] _15015;
    wire [63:0] _15016;
    wire [62:0] _15017;
    wire [63:0] _15019;
    wire _15020;
    wire _15021;
    wire _15009;
    wire [63:0] _15006;
    wire [63:0] _15007;
    wire [62:0] _15008;
    wire [63:0] _15010;
    wire _15011;
    wire _15012;
    wire _15000;
    wire [63:0] _14997;
    wire [63:0] _14998;
    wire [62:0] _14999;
    wire [63:0] _15001;
    wire _15002;
    wire _15003;
    wire _14991;
    wire [63:0] _14988;
    wire [63:0] _14989;
    wire [62:0] _14990;
    wire [63:0] _14992;
    wire _14993;
    wire _14994;
    wire _14982;
    wire [63:0] _14979;
    wire [63:0] _14980;
    wire [62:0] _14981;
    wire [63:0] _14983;
    wire _14984;
    wire _14985;
    wire _14973;
    wire [63:0] _14970;
    wire [63:0] _14971;
    wire [62:0] _14972;
    wire [63:0] _14974;
    wire _14975;
    wire _14976;
    wire _14964;
    wire [63:0] _14961;
    wire [63:0] _14962;
    wire [62:0] _14963;
    wire [63:0] _14965;
    wire _14966;
    wire _14967;
    wire _14955;
    wire [63:0] _14952;
    wire [63:0] _14953;
    wire [62:0] _14954;
    wire [63:0] _14956;
    wire _14957;
    wire _14958;
    wire _14946;
    wire [63:0] _14943;
    wire [63:0] _14944;
    wire [62:0] _14945;
    wire [63:0] _14947;
    wire _14948;
    wire _14949;
    wire _14937;
    wire [63:0] _14934;
    wire [63:0] _14935;
    wire [62:0] _14936;
    wire [63:0] _14938;
    wire _14939;
    wire _14940;
    wire _14928;
    wire [63:0] _14925;
    wire [63:0] _14926;
    wire [62:0] _14927;
    wire [63:0] _14929;
    wire _14930;
    wire _14931;
    wire _14919;
    wire [63:0] _14916;
    wire [63:0] _14917;
    wire [62:0] _14918;
    wire [63:0] _14920;
    wire _14921;
    wire _14922;
    wire _14910;
    wire [63:0] _14907;
    wire [63:0] _14908;
    wire [62:0] _14909;
    wire [63:0] _14911;
    wire _14912;
    wire _14913;
    wire _14901;
    wire [63:0] _14898;
    wire [63:0] _14899;
    wire [62:0] _14900;
    wire [63:0] _14902;
    wire _14903;
    wire _14904;
    wire _14892;
    wire [63:0] _14889;
    wire [63:0] _14890;
    wire [62:0] _14891;
    wire [63:0] _14893;
    wire _14894;
    wire _14895;
    wire _14883;
    wire [63:0] _14880;
    wire [63:0] _14881;
    wire [62:0] _14882;
    wire [63:0] _14884;
    wire _14885;
    wire _14886;
    wire _14874;
    wire [63:0] _14871;
    wire [63:0] _14872;
    wire [62:0] _14873;
    wire [63:0] _14875;
    wire _14876;
    wire _14877;
    wire _14865;
    wire [63:0] _14862;
    wire [63:0] _14863;
    wire [62:0] _14864;
    wire [63:0] _14866;
    wire _14867;
    wire _14868;
    wire _14856;
    wire [63:0] _14853;
    wire [63:0] _14854;
    wire [62:0] _14855;
    wire [63:0] _14857;
    wire _14858;
    wire _14859;
    wire _14847;
    wire [63:0] _14844;
    wire [63:0] _14845;
    wire [62:0] _14846;
    wire [63:0] _14848;
    wire _14849;
    wire _14850;
    wire _14838;
    wire [63:0] _14835;
    wire [63:0] _14836;
    wire [62:0] _14837;
    wire [63:0] _14839;
    wire _14840;
    wire _14841;
    wire _14829;
    wire [63:0] _14826;
    wire [63:0] _14827;
    wire [62:0] _14828;
    wire [63:0] _14830;
    wire _14831;
    wire _14832;
    wire _14820;
    wire [63:0] _14817;
    wire [63:0] _14818;
    wire [62:0] _14819;
    wire [63:0] _14821;
    wire _14822;
    wire _14823;
    wire _14811;
    wire [63:0] _14808;
    wire [63:0] _14809;
    wire [62:0] _14810;
    wire [63:0] _14812;
    wire _14813;
    wire _14814;
    wire _14802;
    wire [63:0] _14799;
    wire [63:0] _14800;
    wire [62:0] _14801;
    wire [63:0] _14803;
    wire _14804;
    wire _14805;
    wire _14793;
    wire [63:0] _14790;
    wire [63:0] _14791;
    wire [62:0] _14792;
    wire [63:0] _14794;
    wire _14795;
    wire _14796;
    wire _14784;
    wire [63:0] _14781;
    wire [63:0] _14782;
    wire [62:0] _14783;
    wire [63:0] _14785;
    wire _14786;
    wire _14787;
    wire _14775;
    wire [63:0] _14772;
    wire [63:0] _14773;
    wire [62:0] _14774;
    wire [63:0] _14776;
    wire _14777;
    wire _14778;
    wire _14766;
    wire [63:0] _14763;
    wire [63:0] _14764;
    wire [62:0] _14765;
    wire [63:0] _14767;
    wire _14768;
    wire _14769;
    wire _14757;
    wire [63:0] _14754;
    wire [63:0] _14755;
    wire [62:0] _14756;
    wire [63:0] _14758;
    wire _14759;
    wire _14760;
    wire _14748;
    wire [63:0] _14745;
    wire [63:0] _14746;
    wire [62:0] _14747;
    wire [63:0] _14749;
    wire _14750;
    wire _14751;
    wire _14739;
    wire [63:0] _14736;
    wire [63:0] _14737;
    wire [62:0] _14738;
    wire [63:0] _14740;
    wire _14741;
    wire _14742;
    wire _14730;
    wire [63:0] _14727;
    wire [63:0] _14728;
    wire [62:0] _14729;
    wire [63:0] _14731;
    wire _14732;
    wire _14733;
    wire _14721;
    wire [63:0] _14718;
    wire [63:0] _14719;
    wire [62:0] _14720;
    wire [63:0] _14722;
    wire _14723;
    wire _14724;
    wire _14712;
    wire [63:0] _14709;
    wire [63:0] _14710;
    wire [62:0] _14711;
    wire [63:0] _14713;
    wire _14714;
    wire _14715;
    wire _14703;
    wire [63:0] _14700;
    wire [63:0] _14701;
    wire [62:0] _14702;
    wire [63:0] _14704;
    wire _14705;
    wire _14706;
    wire _14694;
    wire [63:0] _14691;
    wire [63:0] _14692;
    wire [62:0] _14693;
    wire [63:0] _14695;
    wire _14696;
    wire _14697;
    wire _14685;
    wire [63:0] _14682;
    wire [63:0] _14683;
    wire [62:0] _14684;
    wire [63:0] _14686;
    wire _14687;
    wire _14688;
    wire _14676;
    wire [63:0] _14673;
    wire [63:0] _14674;
    wire [62:0] _14675;
    wire [63:0] _14677;
    wire _14678;
    wire _14679;
    wire _14667;
    wire [63:0] _14664;
    wire [63:0] _14665;
    wire [62:0] _14666;
    wire [63:0] _14668;
    wire _14669;
    wire _14670;
    wire _14658;
    wire [63:0] _14655;
    wire [63:0] _14656;
    wire [62:0] _14657;
    wire [63:0] _14659;
    wire _14660;
    wire _14661;
    wire _14649;
    wire [63:0] _14646;
    wire [63:0] _14647;
    wire [62:0] _14648;
    wire [63:0] _14650;
    wire _14651;
    wire _14652;
    wire _14640;
    wire [63:0] _14637;
    wire [63:0] _14638;
    wire [62:0] _14639;
    wire [63:0] _14641;
    wire _14642;
    wire _14643;
    wire _14631;
    wire [63:0] _14628;
    wire [63:0] _14629;
    wire [62:0] _14630;
    wire [63:0] _14632;
    wire _14633;
    wire _14634;
    wire _14622;
    wire [63:0] _14619;
    wire [63:0] _14620;
    wire [62:0] _14621;
    wire [63:0] _14623;
    wire _14624;
    wire _14625;
    wire _14613;
    wire [63:0] _14610;
    wire [63:0] _14611;
    wire [62:0] _14612;
    wire [63:0] _14614;
    wire _14615;
    wire _14616;
    wire [63:0] _14603;
    wire _14604;
    wire [63:0] _14605;
    wire _14606;
    wire _14607;
    wire [63:0] _14608;
    wire [62:0] _14609;
    wire [63:0] _14617;
    wire [62:0] _14618;
    wire [63:0] _14626;
    wire [62:0] _14627;
    wire [63:0] _14635;
    wire [62:0] _14636;
    wire [63:0] _14644;
    wire [62:0] _14645;
    wire [63:0] _14653;
    wire [62:0] _14654;
    wire [63:0] _14662;
    wire [62:0] _14663;
    wire [63:0] _14671;
    wire [62:0] _14672;
    wire [63:0] _14680;
    wire [62:0] _14681;
    wire [63:0] _14689;
    wire [62:0] _14690;
    wire [63:0] _14698;
    wire [62:0] _14699;
    wire [63:0] _14707;
    wire [62:0] _14708;
    wire [63:0] _14716;
    wire [62:0] _14717;
    wire [63:0] _14725;
    wire [62:0] _14726;
    wire [63:0] _14734;
    wire [62:0] _14735;
    wire [63:0] _14743;
    wire [62:0] _14744;
    wire [63:0] _14752;
    wire [62:0] _14753;
    wire [63:0] _14761;
    wire [62:0] _14762;
    wire [63:0] _14770;
    wire [62:0] _14771;
    wire [63:0] _14779;
    wire [62:0] _14780;
    wire [63:0] _14788;
    wire [62:0] _14789;
    wire [63:0] _14797;
    wire [62:0] _14798;
    wire [63:0] _14806;
    wire [62:0] _14807;
    wire [63:0] _14815;
    wire [62:0] _14816;
    wire [63:0] _14824;
    wire [62:0] _14825;
    wire [63:0] _14833;
    wire [62:0] _14834;
    wire [63:0] _14842;
    wire [62:0] _14843;
    wire [63:0] _14851;
    wire [62:0] _14852;
    wire [63:0] _14860;
    wire [62:0] _14861;
    wire [63:0] _14869;
    wire [62:0] _14870;
    wire [63:0] _14878;
    wire [62:0] _14879;
    wire [63:0] _14887;
    wire [62:0] _14888;
    wire [63:0] _14896;
    wire [62:0] _14897;
    wire [63:0] _14905;
    wire [62:0] _14906;
    wire [63:0] _14914;
    wire [62:0] _14915;
    wire [63:0] _14923;
    wire [62:0] _14924;
    wire [63:0] _14932;
    wire [62:0] _14933;
    wire [63:0] _14941;
    wire [62:0] _14942;
    wire [63:0] _14950;
    wire [62:0] _14951;
    wire [63:0] _14959;
    wire [62:0] _14960;
    wire [63:0] _14968;
    wire [62:0] _14969;
    wire [63:0] _14977;
    wire [62:0] _14978;
    wire [63:0] _14986;
    wire [62:0] _14987;
    wire [63:0] _14995;
    wire [62:0] _14996;
    wire [63:0] _15004;
    wire [62:0] _15005;
    wire [63:0] _15013;
    wire [62:0] _15014;
    wire [63:0] _15022;
    wire [62:0] _15023;
    wire [63:0] _15031;
    wire [62:0] _15032;
    wire [63:0] _15040;
    wire [62:0] _15041;
    wire [63:0] _15049;
    wire [62:0] _15050;
    wire [63:0] _15058;
    wire [62:0] _15059;
    wire [63:0] _15067;
    wire [62:0] _15068;
    wire [63:0] _15076;
    wire [62:0] _15077;
    wire [63:0] _15085;
    wire [62:0] _15086;
    wire [63:0] _15094;
    wire [62:0] _15095;
    wire [63:0] _15103;
    wire [62:0] _15104;
    wire [63:0] _15112;
    wire [62:0] _15113;
    wire [63:0] _15121;
    wire [62:0] _15122;
    wire [63:0] _15130;
    wire [62:0] _15131;
    wire [63:0] _15139;
    wire [62:0] _15140;
    wire [63:0] _15148;
    wire [62:0] _15149;
    wire [63:0] _15157;
    wire [62:0] _15158;
    wire [63:0] _15166;
    wire [62:0] _15167;
    wire [63:0] _15175;
    wire [63:0] _15177;
    wire [127:0] _15178;
    wire [63:0] _15179;
    wire [63:0] _15761;
    wire _14589;
    wire [63:0] _14586;
    wire [63:0] _14587;
    wire [62:0] _14588;
    wire [63:0] _14590;
    wire _14591;
    wire _14592;
    wire _14580;
    wire [63:0] _14577;
    wire [63:0] _14578;
    wire [62:0] _14579;
    wire [63:0] _14581;
    wire _14582;
    wire _14583;
    wire _14571;
    wire [63:0] _14568;
    wire [63:0] _14569;
    wire [62:0] _14570;
    wire [63:0] _14572;
    wire _14573;
    wire _14574;
    wire _14562;
    wire [63:0] _14559;
    wire [63:0] _14560;
    wire [62:0] _14561;
    wire [63:0] _14563;
    wire _14564;
    wire _14565;
    wire _14553;
    wire [63:0] _14550;
    wire [63:0] _14551;
    wire [62:0] _14552;
    wire [63:0] _14554;
    wire _14555;
    wire _14556;
    wire _14544;
    wire [63:0] _14541;
    wire [63:0] _14542;
    wire [62:0] _14543;
    wire [63:0] _14545;
    wire _14546;
    wire _14547;
    wire _14535;
    wire [63:0] _14532;
    wire [63:0] _14533;
    wire [62:0] _14534;
    wire [63:0] _14536;
    wire _14537;
    wire _14538;
    wire _14526;
    wire [63:0] _14523;
    wire [63:0] _14524;
    wire [62:0] _14525;
    wire [63:0] _14527;
    wire _14528;
    wire _14529;
    wire _14517;
    wire [63:0] _14514;
    wire [63:0] _14515;
    wire [62:0] _14516;
    wire [63:0] _14518;
    wire _14519;
    wire _14520;
    wire _14508;
    wire [63:0] _14505;
    wire [63:0] _14506;
    wire [62:0] _14507;
    wire [63:0] _14509;
    wire _14510;
    wire _14511;
    wire _14499;
    wire [63:0] _14496;
    wire [63:0] _14497;
    wire [62:0] _14498;
    wire [63:0] _14500;
    wire _14501;
    wire _14502;
    wire _14490;
    wire [63:0] _14487;
    wire [63:0] _14488;
    wire [62:0] _14489;
    wire [63:0] _14491;
    wire _14492;
    wire _14493;
    wire _14481;
    wire [63:0] _14478;
    wire [63:0] _14479;
    wire [62:0] _14480;
    wire [63:0] _14482;
    wire _14483;
    wire _14484;
    wire _14472;
    wire [63:0] _14469;
    wire [63:0] _14470;
    wire [62:0] _14471;
    wire [63:0] _14473;
    wire _14474;
    wire _14475;
    wire _14463;
    wire [63:0] _14460;
    wire [63:0] _14461;
    wire [62:0] _14462;
    wire [63:0] _14464;
    wire _14465;
    wire _14466;
    wire _14454;
    wire [63:0] _14451;
    wire [63:0] _14452;
    wire [62:0] _14453;
    wire [63:0] _14455;
    wire _14456;
    wire _14457;
    wire _14445;
    wire [63:0] _14442;
    wire [63:0] _14443;
    wire [62:0] _14444;
    wire [63:0] _14446;
    wire _14447;
    wire _14448;
    wire _14436;
    wire [63:0] _14433;
    wire [63:0] _14434;
    wire [62:0] _14435;
    wire [63:0] _14437;
    wire _14438;
    wire _14439;
    wire _14427;
    wire [63:0] _14424;
    wire [63:0] _14425;
    wire [62:0] _14426;
    wire [63:0] _14428;
    wire _14429;
    wire _14430;
    wire _14418;
    wire [63:0] _14415;
    wire [63:0] _14416;
    wire [62:0] _14417;
    wire [63:0] _14419;
    wire _14420;
    wire _14421;
    wire _14409;
    wire [63:0] _14406;
    wire [63:0] _14407;
    wire [62:0] _14408;
    wire [63:0] _14410;
    wire _14411;
    wire _14412;
    wire _14400;
    wire [63:0] _14397;
    wire [63:0] _14398;
    wire [62:0] _14399;
    wire [63:0] _14401;
    wire _14402;
    wire _14403;
    wire _14391;
    wire [63:0] _14388;
    wire [63:0] _14389;
    wire [62:0] _14390;
    wire [63:0] _14392;
    wire _14393;
    wire _14394;
    wire _14382;
    wire [63:0] _14379;
    wire [63:0] _14380;
    wire [62:0] _14381;
    wire [63:0] _14383;
    wire _14384;
    wire _14385;
    wire _14373;
    wire [63:0] _14370;
    wire [63:0] _14371;
    wire [62:0] _14372;
    wire [63:0] _14374;
    wire _14375;
    wire _14376;
    wire _14364;
    wire [63:0] _14361;
    wire [63:0] _14362;
    wire [62:0] _14363;
    wire [63:0] _14365;
    wire _14366;
    wire _14367;
    wire _14355;
    wire [63:0] _14352;
    wire [63:0] _14353;
    wire [62:0] _14354;
    wire [63:0] _14356;
    wire _14357;
    wire _14358;
    wire _14346;
    wire [63:0] _14343;
    wire [63:0] _14344;
    wire [62:0] _14345;
    wire [63:0] _14347;
    wire _14348;
    wire _14349;
    wire _14337;
    wire [63:0] _14334;
    wire [63:0] _14335;
    wire [62:0] _14336;
    wire [63:0] _14338;
    wire _14339;
    wire _14340;
    wire _14328;
    wire [63:0] _14325;
    wire [63:0] _14326;
    wire [62:0] _14327;
    wire [63:0] _14329;
    wire _14330;
    wire _14331;
    wire _14319;
    wire [63:0] _14316;
    wire [63:0] _14317;
    wire [62:0] _14318;
    wire [63:0] _14320;
    wire _14321;
    wire _14322;
    wire _14310;
    wire [63:0] _14307;
    wire [63:0] _14308;
    wire [62:0] _14309;
    wire [63:0] _14311;
    wire _14312;
    wire _14313;
    wire _14301;
    wire [63:0] _14298;
    wire [63:0] _14299;
    wire [62:0] _14300;
    wire [63:0] _14302;
    wire _14303;
    wire _14304;
    wire _14292;
    wire [63:0] _14289;
    wire [63:0] _14290;
    wire [62:0] _14291;
    wire [63:0] _14293;
    wire _14294;
    wire _14295;
    wire _14283;
    wire [63:0] _14280;
    wire [63:0] _14281;
    wire [62:0] _14282;
    wire [63:0] _14284;
    wire _14285;
    wire _14286;
    wire _14274;
    wire [63:0] _14271;
    wire [63:0] _14272;
    wire [62:0] _14273;
    wire [63:0] _14275;
    wire _14276;
    wire _14277;
    wire _14265;
    wire [63:0] _14262;
    wire [63:0] _14263;
    wire [62:0] _14264;
    wire [63:0] _14266;
    wire _14267;
    wire _14268;
    wire _14256;
    wire [63:0] _14253;
    wire [63:0] _14254;
    wire [62:0] _14255;
    wire [63:0] _14257;
    wire _14258;
    wire _14259;
    wire _14247;
    wire [63:0] _14244;
    wire [63:0] _14245;
    wire [62:0] _14246;
    wire [63:0] _14248;
    wire _14249;
    wire _14250;
    wire _14238;
    wire [63:0] _14235;
    wire [63:0] _14236;
    wire [62:0] _14237;
    wire [63:0] _14239;
    wire _14240;
    wire _14241;
    wire _14229;
    wire [63:0] _14226;
    wire [63:0] _14227;
    wire [62:0] _14228;
    wire [63:0] _14230;
    wire _14231;
    wire _14232;
    wire _14220;
    wire [63:0] _14217;
    wire [63:0] _14218;
    wire [62:0] _14219;
    wire [63:0] _14221;
    wire _14222;
    wire _14223;
    wire _14211;
    wire [63:0] _14208;
    wire [63:0] _14209;
    wire [62:0] _14210;
    wire [63:0] _14212;
    wire _14213;
    wire _14214;
    wire _14202;
    wire [63:0] _14199;
    wire [63:0] _14200;
    wire [62:0] _14201;
    wire [63:0] _14203;
    wire _14204;
    wire _14205;
    wire _14193;
    wire [63:0] _14190;
    wire [63:0] _14191;
    wire [62:0] _14192;
    wire [63:0] _14194;
    wire _14195;
    wire _14196;
    wire _14184;
    wire [63:0] _14181;
    wire [63:0] _14182;
    wire [62:0] _14183;
    wire [63:0] _14185;
    wire _14186;
    wire _14187;
    wire _14175;
    wire [63:0] _14172;
    wire [63:0] _14173;
    wire [62:0] _14174;
    wire [63:0] _14176;
    wire _14177;
    wire _14178;
    wire _14166;
    wire [63:0] _14163;
    wire [63:0] _14164;
    wire [62:0] _14165;
    wire [63:0] _14167;
    wire _14168;
    wire _14169;
    wire _14157;
    wire [63:0] _14154;
    wire [63:0] _14155;
    wire [62:0] _14156;
    wire [63:0] _14158;
    wire _14159;
    wire _14160;
    wire _14148;
    wire [63:0] _14145;
    wire [63:0] _14146;
    wire [62:0] _14147;
    wire [63:0] _14149;
    wire _14150;
    wire _14151;
    wire _14139;
    wire [63:0] _14136;
    wire [63:0] _14137;
    wire [62:0] _14138;
    wire [63:0] _14140;
    wire _14141;
    wire _14142;
    wire _14130;
    wire [63:0] _14127;
    wire [63:0] _14128;
    wire [62:0] _14129;
    wire [63:0] _14131;
    wire _14132;
    wire _14133;
    wire _14121;
    wire [63:0] _14118;
    wire [63:0] _14119;
    wire [62:0] _14120;
    wire [63:0] _14122;
    wire _14123;
    wire _14124;
    wire _14112;
    wire [63:0] _14109;
    wire [63:0] _14110;
    wire [62:0] _14111;
    wire [63:0] _14113;
    wire _14114;
    wire _14115;
    wire _14103;
    wire [63:0] _14100;
    wire [63:0] _14101;
    wire [62:0] _14102;
    wire [63:0] _14104;
    wire _14105;
    wire _14106;
    wire _14094;
    wire [63:0] _14091;
    wire [63:0] _14092;
    wire [62:0] _14093;
    wire [63:0] _14095;
    wire _14096;
    wire _14097;
    wire _14085;
    wire [63:0] _14082;
    wire [63:0] _14083;
    wire [62:0] _14084;
    wire [63:0] _14086;
    wire _14087;
    wire _14088;
    wire _14076;
    wire [63:0] _14073;
    wire [63:0] _14074;
    wire [62:0] _14075;
    wire [63:0] _14077;
    wire _14078;
    wire _14079;
    wire _14067;
    wire [63:0] _14064;
    wire [63:0] _14065;
    wire [62:0] _14066;
    wire [63:0] _14068;
    wire _14069;
    wire _14070;
    wire _14058;
    wire [63:0] _14055;
    wire [63:0] _14056;
    wire [62:0] _14057;
    wire [63:0] _14059;
    wire _14060;
    wire _14061;
    wire _14049;
    wire [63:0] _14046;
    wire [63:0] _14047;
    wire [62:0] _14048;
    wire [63:0] _14050;
    wire _14051;
    wire _14052;
    wire _14040;
    wire [63:0] _14037;
    wire [63:0] _14038;
    wire [62:0] _14039;
    wire [63:0] _14041;
    wire _14042;
    wire _14043;
    wire _14031;
    wire [63:0] _14028;
    wire [63:0] _14029;
    wire [62:0] _14030;
    wire [63:0] _14032;
    wire _14033;
    wire _14034;
    wire [63:0] _14023;
    wire [63:0] _14019;
    wire [63:0] _14020;
    wire _14021;
    wire [63:0] _14022;
    wire _14024;
    wire _14025;
    wire [63:0] _14026;
    wire [62:0] _14027;
    wire [63:0] _14035;
    wire [62:0] _14036;
    wire [63:0] _14044;
    wire [62:0] _14045;
    wire [63:0] _14053;
    wire [62:0] _14054;
    wire [63:0] _14062;
    wire [62:0] _14063;
    wire [63:0] _14071;
    wire [62:0] _14072;
    wire [63:0] _14080;
    wire [62:0] _14081;
    wire [63:0] _14089;
    wire [62:0] _14090;
    wire [63:0] _14098;
    wire [62:0] _14099;
    wire [63:0] _14107;
    wire [62:0] _14108;
    wire [63:0] _14116;
    wire [62:0] _14117;
    wire [63:0] _14125;
    wire [62:0] _14126;
    wire [63:0] _14134;
    wire [62:0] _14135;
    wire [63:0] _14143;
    wire [62:0] _14144;
    wire [63:0] _14152;
    wire [62:0] _14153;
    wire [63:0] _14161;
    wire [62:0] _14162;
    wire [63:0] _14170;
    wire [62:0] _14171;
    wire [63:0] _14179;
    wire [62:0] _14180;
    wire [63:0] _14188;
    wire [62:0] _14189;
    wire [63:0] _14197;
    wire [62:0] _14198;
    wire [63:0] _14206;
    wire [62:0] _14207;
    wire [63:0] _14215;
    wire [62:0] _14216;
    wire [63:0] _14224;
    wire [62:0] _14225;
    wire [63:0] _14233;
    wire [62:0] _14234;
    wire [63:0] _14242;
    wire [62:0] _14243;
    wire [63:0] _14251;
    wire [62:0] _14252;
    wire [63:0] _14260;
    wire [62:0] _14261;
    wire [63:0] _14269;
    wire [62:0] _14270;
    wire [63:0] _14278;
    wire [62:0] _14279;
    wire [63:0] _14287;
    wire [62:0] _14288;
    wire [63:0] _14296;
    wire [62:0] _14297;
    wire [63:0] _14305;
    wire [62:0] _14306;
    wire [63:0] _14314;
    wire [62:0] _14315;
    wire [63:0] _14323;
    wire [62:0] _14324;
    wire [63:0] _14332;
    wire [62:0] _14333;
    wire [63:0] _14341;
    wire [62:0] _14342;
    wire [63:0] _14350;
    wire [62:0] _14351;
    wire [63:0] _14359;
    wire [62:0] _14360;
    wire [63:0] _14368;
    wire [62:0] _14369;
    wire [63:0] _14377;
    wire [62:0] _14378;
    wire [63:0] _14386;
    wire [62:0] _14387;
    wire [63:0] _14395;
    wire [62:0] _14396;
    wire [63:0] _14404;
    wire [62:0] _14405;
    wire [63:0] _14413;
    wire [62:0] _14414;
    wire [63:0] _14422;
    wire [62:0] _14423;
    wire [63:0] _14431;
    wire [62:0] _14432;
    wire [63:0] _14440;
    wire [62:0] _14441;
    wire [63:0] _14449;
    wire [62:0] _14450;
    wire [63:0] _14458;
    wire [62:0] _14459;
    wire [63:0] _14467;
    wire [62:0] _14468;
    wire [63:0] _14476;
    wire [62:0] _14477;
    wire [63:0] _14485;
    wire [62:0] _14486;
    wire [63:0] _14494;
    wire [62:0] _14495;
    wire [63:0] _14503;
    wire [62:0] _14504;
    wire [63:0] _14512;
    wire [62:0] _14513;
    wire [63:0] _14521;
    wire [62:0] _14522;
    wire [63:0] _14530;
    wire [62:0] _14531;
    wire [63:0] _14539;
    wire [62:0] _14540;
    wire [63:0] _14548;
    wire [62:0] _14549;
    wire [63:0] _14557;
    wire [62:0] _14558;
    wire [63:0] _14566;
    wire [62:0] _14567;
    wire [63:0] _14575;
    wire [62:0] _14576;
    wire [63:0] _14584;
    wire [62:0] _14585;
    wire [63:0] _14593;
    wire [127:0] _14594;
    wire [63:0] _14595;
    wire _14596;
    wire [63:0] _14597;
    wire [63:0] _14013;
    wire _14014;
    wire [63:0] _14015;
    wire _14598;
    wire _14599;
    wire [63:0] _15762;
    wire _14003;
    wire [63:0] _14000;
    wire [63:0] _14001;
    wire [62:0] _14002;
    wire [63:0] _14004;
    wire _14005;
    wire _14006;
    wire _13994;
    wire [63:0] _13991;
    wire [63:0] _13992;
    wire [62:0] _13993;
    wire [63:0] _13995;
    wire _13996;
    wire _13997;
    wire _13985;
    wire [63:0] _13982;
    wire [63:0] _13983;
    wire [62:0] _13984;
    wire [63:0] _13986;
    wire _13987;
    wire _13988;
    wire _13976;
    wire [63:0] _13973;
    wire [63:0] _13974;
    wire [62:0] _13975;
    wire [63:0] _13977;
    wire _13978;
    wire _13979;
    wire _13967;
    wire [63:0] _13964;
    wire [63:0] _13965;
    wire [62:0] _13966;
    wire [63:0] _13968;
    wire _13969;
    wire _13970;
    wire _13958;
    wire [63:0] _13955;
    wire [63:0] _13956;
    wire [62:0] _13957;
    wire [63:0] _13959;
    wire _13960;
    wire _13961;
    wire _13949;
    wire [63:0] _13946;
    wire [63:0] _13947;
    wire [62:0] _13948;
    wire [63:0] _13950;
    wire _13951;
    wire _13952;
    wire _13940;
    wire [63:0] _13937;
    wire [63:0] _13938;
    wire [62:0] _13939;
    wire [63:0] _13941;
    wire _13942;
    wire _13943;
    wire _13931;
    wire [63:0] _13928;
    wire [63:0] _13929;
    wire [62:0] _13930;
    wire [63:0] _13932;
    wire _13933;
    wire _13934;
    wire _13922;
    wire [63:0] _13919;
    wire [63:0] _13920;
    wire [62:0] _13921;
    wire [63:0] _13923;
    wire _13924;
    wire _13925;
    wire _13913;
    wire [63:0] _13910;
    wire [63:0] _13911;
    wire [62:0] _13912;
    wire [63:0] _13914;
    wire _13915;
    wire _13916;
    wire _13904;
    wire [63:0] _13901;
    wire [63:0] _13902;
    wire [62:0] _13903;
    wire [63:0] _13905;
    wire _13906;
    wire _13907;
    wire _13895;
    wire [63:0] _13892;
    wire [63:0] _13893;
    wire [62:0] _13894;
    wire [63:0] _13896;
    wire _13897;
    wire _13898;
    wire _13886;
    wire [63:0] _13883;
    wire [63:0] _13884;
    wire [62:0] _13885;
    wire [63:0] _13887;
    wire _13888;
    wire _13889;
    wire _13877;
    wire [63:0] _13874;
    wire [63:0] _13875;
    wire [62:0] _13876;
    wire [63:0] _13878;
    wire _13879;
    wire _13880;
    wire _13868;
    wire [63:0] _13865;
    wire [63:0] _13866;
    wire [62:0] _13867;
    wire [63:0] _13869;
    wire _13870;
    wire _13871;
    wire _13859;
    wire [63:0] _13856;
    wire [63:0] _13857;
    wire [62:0] _13858;
    wire [63:0] _13860;
    wire _13861;
    wire _13862;
    wire _13850;
    wire [63:0] _13847;
    wire [63:0] _13848;
    wire [62:0] _13849;
    wire [63:0] _13851;
    wire _13852;
    wire _13853;
    wire _13841;
    wire [63:0] _13838;
    wire [63:0] _13839;
    wire [62:0] _13840;
    wire [63:0] _13842;
    wire _13843;
    wire _13844;
    wire _13832;
    wire [63:0] _13829;
    wire [63:0] _13830;
    wire [62:0] _13831;
    wire [63:0] _13833;
    wire _13834;
    wire _13835;
    wire _13823;
    wire [63:0] _13820;
    wire [63:0] _13821;
    wire [62:0] _13822;
    wire [63:0] _13824;
    wire _13825;
    wire _13826;
    wire _13814;
    wire [63:0] _13811;
    wire [63:0] _13812;
    wire [62:0] _13813;
    wire [63:0] _13815;
    wire _13816;
    wire _13817;
    wire _13805;
    wire [63:0] _13802;
    wire [63:0] _13803;
    wire [62:0] _13804;
    wire [63:0] _13806;
    wire _13807;
    wire _13808;
    wire _13796;
    wire [63:0] _13793;
    wire [63:0] _13794;
    wire [62:0] _13795;
    wire [63:0] _13797;
    wire _13798;
    wire _13799;
    wire _13787;
    wire [63:0] _13784;
    wire [63:0] _13785;
    wire [62:0] _13786;
    wire [63:0] _13788;
    wire _13789;
    wire _13790;
    wire _13778;
    wire [63:0] _13775;
    wire [63:0] _13776;
    wire [62:0] _13777;
    wire [63:0] _13779;
    wire _13780;
    wire _13781;
    wire _13769;
    wire [63:0] _13766;
    wire [63:0] _13767;
    wire [62:0] _13768;
    wire [63:0] _13770;
    wire _13771;
    wire _13772;
    wire _13760;
    wire [63:0] _13757;
    wire [63:0] _13758;
    wire [62:0] _13759;
    wire [63:0] _13761;
    wire _13762;
    wire _13763;
    wire _13751;
    wire [63:0] _13748;
    wire [63:0] _13749;
    wire [62:0] _13750;
    wire [63:0] _13752;
    wire _13753;
    wire _13754;
    wire _13742;
    wire [63:0] _13739;
    wire [63:0] _13740;
    wire [62:0] _13741;
    wire [63:0] _13743;
    wire _13744;
    wire _13745;
    wire _13733;
    wire [63:0] _13730;
    wire [63:0] _13731;
    wire [62:0] _13732;
    wire [63:0] _13734;
    wire _13735;
    wire _13736;
    wire _13724;
    wire [63:0] _13721;
    wire [63:0] _13722;
    wire [62:0] _13723;
    wire [63:0] _13725;
    wire _13726;
    wire _13727;
    wire _13715;
    wire [63:0] _13712;
    wire [63:0] _13713;
    wire [62:0] _13714;
    wire [63:0] _13716;
    wire _13717;
    wire _13718;
    wire _13706;
    wire [63:0] _13703;
    wire [63:0] _13704;
    wire [62:0] _13705;
    wire [63:0] _13707;
    wire _13708;
    wire _13709;
    wire _13697;
    wire [63:0] _13694;
    wire [63:0] _13695;
    wire [62:0] _13696;
    wire [63:0] _13698;
    wire _13699;
    wire _13700;
    wire _13688;
    wire [63:0] _13685;
    wire [63:0] _13686;
    wire [62:0] _13687;
    wire [63:0] _13689;
    wire _13690;
    wire _13691;
    wire _13679;
    wire [63:0] _13676;
    wire [63:0] _13677;
    wire [62:0] _13678;
    wire [63:0] _13680;
    wire _13681;
    wire _13682;
    wire _13670;
    wire [63:0] _13667;
    wire [63:0] _13668;
    wire [62:0] _13669;
    wire [63:0] _13671;
    wire _13672;
    wire _13673;
    wire _13661;
    wire [63:0] _13658;
    wire [63:0] _13659;
    wire [62:0] _13660;
    wire [63:0] _13662;
    wire _13663;
    wire _13664;
    wire _13652;
    wire [63:0] _13649;
    wire [63:0] _13650;
    wire [62:0] _13651;
    wire [63:0] _13653;
    wire _13654;
    wire _13655;
    wire _13643;
    wire [63:0] _13640;
    wire [63:0] _13641;
    wire [62:0] _13642;
    wire [63:0] _13644;
    wire _13645;
    wire _13646;
    wire _13634;
    wire [63:0] _13631;
    wire [63:0] _13632;
    wire [62:0] _13633;
    wire [63:0] _13635;
    wire _13636;
    wire _13637;
    wire _13625;
    wire [63:0] _13622;
    wire [63:0] _13623;
    wire [62:0] _13624;
    wire [63:0] _13626;
    wire _13627;
    wire _13628;
    wire _13616;
    wire [63:0] _13613;
    wire [63:0] _13614;
    wire [62:0] _13615;
    wire [63:0] _13617;
    wire _13618;
    wire _13619;
    wire _13607;
    wire [63:0] _13604;
    wire [63:0] _13605;
    wire [62:0] _13606;
    wire [63:0] _13608;
    wire _13609;
    wire _13610;
    wire _13598;
    wire [63:0] _13595;
    wire [63:0] _13596;
    wire [62:0] _13597;
    wire [63:0] _13599;
    wire _13600;
    wire _13601;
    wire _13589;
    wire [63:0] _13586;
    wire [63:0] _13587;
    wire [62:0] _13588;
    wire [63:0] _13590;
    wire _13591;
    wire _13592;
    wire _13580;
    wire [63:0] _13577;
    wire [63:0] _13578;
    wire [62:0] _13579;
    wire [63:0] _13581;
    wire _13582;
    wire _13583;
    wire _13571;
    wire [63:0] _13568;
    wire [63:0] _13569;
    wire [62:0] _13570;
    wire [63:0] _13572;
    wire _13573;
    wire _13574;
    wire _13562;
    wire [63:0] _13559;
    wire [63:0] _13560;
    wire [62:0] _13561;
    wire [63:0] _13563;
    wire _13564;
    wire _13565;
    wire _13553;
    wire [63:0] _13550;
    wire [63:0] _13551;
    wire [62:0] _13552;
    wire [63:0] _13554;
    wire _13555;
    wire _13556;
    wire _13544;
    wire [63:0] _13541;
    wire [63:0] _13542;
    wire [62:0] _13543;
    wire [63:0] _13545;
    wire _13546;
    wire _13547;
    wire _13535;
    wire [63:0] _13532;
    wire [63:0] _13533;
    wire [62:0] _13534;
    wire [63:0] _13536;
    wire _13537;
    wire _13538;
    wire _13526;
    wire [63:0] _13523;
    wire [63:0] _13524;
    wire [62:0] _13525;
    wire [63:0] _13527;
    wire _13528;
    wire _13529;
    wire _13517;
    wire [63:0] _13514;
    wire [63:0] _13515;
    wire [62:0] _13516;
    wire [63:0] _13518;
    wire _13519;
    wire _13520;
    wire _13508;
    wire [63:0] _13505;
    wire [63:0] _13506;
    wire [62:0] _13507;
    wire [63:0] _13509;
    wire _13510;
    wire _13511;
    wire _13499;
    wire [63:0] _13496;
    wire [63:0] _13497;
    wire [62:0] _13498;
    wire [63:0] _13500;
    wire _13501;
    wire _13502;
    wire _13490;
    wire [63:0] _13487;
    wire [63:0] _13488;
    wire [62:0] _13489;
    wire [63:0] _13491;
    wire _13492;
    wire _13493;
    wire _13481;
    wire [63:0] _13478;
    wire [63:0] _13479;
    wire [62:0] _13480;
    wire [63:0] _13482;
    wire _13483;
    wire _13484;
    wire _13472;
    wire [63:0] _13469;
    wire [63:0] _13470;
    wire [62:0] _13471;
    wire [63:0] _13473;
    wire _13474;
    wire _13475;
    wire _13463;
    wire [63:0] _13460;
    wire [63:0] _13461;
    wire [62:0] _13462;
    wire [63:0] _13464;
    wire _13465;
    wire _13466;
    wire _13454;
    wire [63:0] _13451;
    wire [63:0] _13452;
    wire [62:0] _13453;
    wire [63:0] _13455;
    wire _13456;
    wire _13457;
    wire _13445;
    wire [63:0] _13442;
    wire [63:0] _13443;
    wire [62:0] _13444;
    wire [63:0] _13446;
    wire _13447;
    wire _13448;
    wire [63:0] _13432;
    wire [127:0] _13433;
    wire [63:0] _13434;
    wire _13435;
    wire [63:0] _13436;
    wire _13438;
    wire _13439;
    wire [63:0] _13440;
    wire [62:0] _13441;
    wire [63:0] _13449;
    wire [62:0] _13450;
    wire [63:0] _13458;
    wire [62:0] _13459;
    wire [63:0] _13467;
    wire [62:0] _13468;
    wire [63:0] _13476;
    wire [62:0] _13477;
    wire [63:0] _13485;
    wire [62:0] _13486;
    wire [63:0] _13494;
    wire [62:0] _13495;
    wire [63:0] _13503;
    wire [62:0] _13504;
    wire [63:0] _13512;
    wire [62:0] _13513;
    wire [63:0] _13521;
    wire [62:0] _13522;
    wire [63:0] _13530;
    wire [62:0] _13531;
    wire [63:0] _13539;
    wire [62:0] _13540;
    wire [63:0] _13548;
    wire [62:0] _13549;
    wire [63:0] _13557;
    wire [62:0] _13558;
    wire [63:0] _13566;
    wire [62:0] _13567;
    wire [63:0] _13575;
    wire [62:0] _13576;
    wire [63:0] _13584;
    wire [62:0] _13585;
    wire [63:0] _13593;
    wire [62:0] _13594;
    wire [63:0] _13602;
    wire [62:0] _13603;
    wire [63:0] _13611;
    wire [62:0] _13612;
    wire [63:0] _13620;
    wire [62:0] _13621;
    wire [63:0] _13629;
    wire [62:0] _13630;
    wire [63:0] _13638;
    wire [62:0] _13639;
    wire [63:0] _13647;
    wire [62:0] _13648;
    wire [63:0] _13656;
    wire [62:0] _13657;
    wire [63:0] _13665;
    wire [62:0] _13666;
    wire [63:0] _13674;
    wire [62:0] _13675;
    wire [63:0] _13683;
    wire [62:0] _13684;
    wire [63:0] _13692;
    wire [62:0] _13693;
    wire [63:0] _13701;
    wire [62:0] _13702;
    wire [63:0] _13710;
    wire [62:0] _13711;
    wire [63:0] _13719;
    wire [62:0] _13720;
    wire [63:0] _13728;
    wire [62:0] _13729;
    wire [63:0] _13737;
    wire [62:0] _13738;
    wire [63:0] _13746;
    wire [62:0] _13747;
    wire [63:0] _13755;
    wire [62:0] _13756;
    wire [63:0] _13764;
    wire [62:0] _13765;
    wire [63:0] _13773;
    wire [62:0] _13774;
    wire [63:0] _13782;
    wire [62:0] _13783;
    wire [63:0] _13791;
    wire [62:0] _13792;
    wire [63:0] _13800;
    wire [62:0] _13801;
    wire [63:0] _13809;
    wire [62:0] _13810;
    wire [63:0] _13818;
    wire [62:0] _13819;
    wire [63:0] _13827;
    wire [62:0] _13828;
    wire [63:0] _13836;
    wire [62:0] _13837;
    wire [63:0] _13845;
    wire [62:0] _13846;
    wire [63:0] _13854;
    wire [62:0] _13855;
    wire [63:0] _13863;
    wire [62:0] _13864;
    wire [63:0] _13872;
    wire [62:0] _13873;
    wire [63:0] _13881;
    wire [62:0] _13882;
    wire [63:0] _13890;
    wire [62:0] _13891;
    wire [63:0] _13899;
    wire [62:0] _13900;
    wire [63:0] _13908;
    wire [62:0] _13909;
    wire [63:0] _13917;
    wire [62:0] _13918;
    wire [63:0] _13926;
    wire [62:0] _13927;
    wire [63:0] _13935;
    wire [62:0] _13936;
    wire [63:0] _13944;
    wire [62:0] _13945;
    wire [63:0] _13953;
    wire [62:0] _13954;
    wire [63:0] _13962;
    wire [62:0] _13963;
    wire [63:0] _13971;
    wire [62:0] _13972;
    wire [63:0] _13980;
    wire [62:0] _13981;
    wire [63:0] _13989;
    wire [62:0] _13990;
    wire [63:0] _13998;
    wire [62:0] _13999;
    wire [63:0] _14007;
    wire [127:0] _14008;
    wire [63:0] _14009;
    wire _13420;
    wire [63:0] _13417;
    wire [63:0] _13418;
    wire [62:0] _13419;
    wire [63:0] _13421;
    wire _13422;
    wire _13423;
    wire _13411;
    wire [63:0] _13408;
    wire [63:0] _13409;
    wire [62:0] _13410;
    wire [63:0] _13412;
    wire _13413;
    wire _13414;
    wire _13402;
    wire [63:0] _13399;
    wire [63:0] _13400;
    wire [62:0] _13401;
    wire [63:0] _13403;
    wire _13404;
    wire _13405;
    wire _13393;
    wire [63:0] _13390;
    wire [63:0] _13391;
    wire [62:0] _13392;
    wire [63:0] _13394;
    wire _13395;
    wire _13396;
    wire _13384;
    wire [63:0] _13381;
    wire [63:0] _13382;
    wire [62:0] _13383;
    wire [63:0] _13385;
    wire _13386;
    wire _13387;
    wire _13375;
    wire [63:0] _13372;
    wire [63:0] _13373;
    wire [62:0] _13374;
    wire [63:0] _13376;
    wire _13377;
    wire _13378;
    wire _13366;
    wire [63:0] _13363;
    wire [63:0] _13364;
    wire [62:0] _13365;
    wire [63:0] _13367;
    wire _13368;
    wire _13369;
    wire _13357;
    wire [63:0] _13354;
    wire [63:0] _13355;
    wire [62:0] _13356;
    wire [63:0] _13358;
    wire _13359;
    wire _13360;
    wire _13348;
    wire [63:0] _13345;
    wire [63:0] _13346;
    wire [62:0] _13347;
    wire [63:0] _13349;
    wire _13350;
    wire _13351;
    wire _13339;
    wire [63:0] _13336;
    wire [63:0] _13337;
    wire [62:0] _13338;
    wire [63:0] _13340;
    wire _13341;
    wire _13342;
    wire _13330;
    wire [63:0] _13327;
    wire [63:0] _13328;
    wire [62:0] _13329;
    wire [63:0] _13331;
    wire _13332;
    wire _13333;
    wire _13321;
    wire [63:0] _13318;
    wire [63:0] _13319;
    wire [62:0] _13320;
    wire [63:0] _13322;
    wire _13323;
    wire _13324;
    wire _13312;
    wire [63:0] _13309;
    wire [63:0] _13310;
    wire [62:0] _13311;
    wire [63:0] _13313;
    wire _13314;
    wire _13315;
    wire _13303;
    wire [63:0] _13300;
    wire [63:0] _13301;
    wire [62:0] _13302;
    wire [63:0] _13304;
    wire _13305;
    wire _13306;
    wire _13294;
    wire [63:0] _13291;
    wire [63:0] _13292;
    wire [62:0] _13293;
    wire [63:0] _13295;
    wire _13296;
    wire _13297;
    wire _13285;
    wire [63:0] _13282;
    wire [63:0] _13283;
    wire [62:0] _13284;
    wire [63:0] _13286;
    wire _13287;
    wire _13288;
    wire _13276;
    wire [63:0] _13273;
    wire [63:0] _13274;
    wire [62:0] _13275;
    wire [63:0] _13277;
    wire _13278;
    wire _13279;
    wire _13267;
    wire [63:0] _13264;
    wire [63:0] _13265;
    wire [62:0] _13266;
    wire [63:0] _13268;
    wire _13269;
    wire _13270;
    wire _13258;
    wire [63:0] _13255;
    wire [63:0] _13256;
    wire [62:0] _13257;
    wire [63:0] _13259;
    wire _13260;
    wire _13261;
    wire _13249;
    wire [63:0] _13246;
    wire [63:0] _13247;
    wire [62:0] _13248;
    wire [63:0] _13250;
    wire _13251;
    wire _13252;
    wire _13240;
    wire [63:0] _13237;
    wire [63:0] _13238;
    wire [62:0] _13239;
    wire [63:0] _13241;
    wire _13242;
    wire _13243;
    wire _13231;
    wire [63:0] _13228;
    wire [63:0] _13229;
    wire [62:0] _13230;
    wire [63:0] _13232;
    wire _13233;
    wire _13234;
    wire _13222;
    wire [63:0] _13219;
    wire [63:0] _13220;
    wire [62:0] _13221;
    wire [63:0] _13223;
    wire _13224;
    wire _13225;
    wire _13213;
    wire [63:0] _13210;
    wire [63:0] _13211;
    wire [62:0] _13212;
    wire [63:0] _13214;
    wire _13215;
    wire _13216;
    wire _13204;
    wire [63:0] _13201;
    wire [63:0] _13202;
    wire [62:0] _13203;
    wire [63:0] _13205;
    wire _13206;
    wire _13207;
    wire _13195;
    wire [63:0] _13192;
    wire [63:0] _13193;
    wire [62:0] _13194;
    wire [63:0] _13196;
    wire _13197;
    wire _13198;
    wire _13186;
    wire [63:0] _13183;
    wire [63:0] _13184;
    wire [62:0] _13185;
    wire [63:0] _13187;
    wire _13188;
    wire _13189;
    wire _13177;
    wire [63:0] _13174;
    wire [63:0] _13175;
    wire [62:0] _13176;
    wire [63:0] _13178;
    wire _13179;
    wire _13180;
    wire _13168;
    wire [63:0] _13165;
    wire [63:0] _13166;
    wire [62:0] _13167;
    wire [63:0] _13169;
    wire _13170;
    wire _13171;
    wire _13159;
    wire [63:0] _13156;
    wire [63:0] _13157;
    wire [62:0] _13158;
    wire [63:0] _13160;
    wire _13161;
    wire _13162;
    wire _13150;
    wire [63:0] _13147;
    wire [63:0] _13148;
    wire [62:0] _13149;
    wire [63:0] _13151;
    wire _13152;
    wire _13153;
    wire _13141;
    wire [63:0] _13138;
    wire [63:0] _13139;
    wire [62:0] _13140;
    wire [63:0] _13142;
    wire _13143;
    wire _13144;
    wire _13132;
    wire [63:0] _13129;
    wire [63:0] _13130;
    wire [62:0] _13131;
    wire [63:0] _13133;
    wire _13134;
    wire _13135;
    wire _13123;
    wire [63:0] _13120;
    wire [63:0] _13121;
    wire [62:0] _13122;
    wire [63:0] _13124;
    wire _13125;
    wire _13126;
    wire _13114;
    wire [63:0] _13111;
    wire [63:0] _13112;
    wire [62:0] _13113;
    wire [63:0] _13115;
    wire _13116;
    wire _13117;
    wire _13105;
    wire [63:0] _13102;
    wire [63:0] _13103;
    wire [62:0] _13104;
    wire [63:0] _13106;
    wire _13107;
    wire _13108;
    wire _13096;
    wire [63:0] _13093;
    wire [63:0] _13094;
    wire [62:0] _13095;
    wire [63:0] _13097;
    wire _13098;
    wire _13099;
    wire _13087;
    wire [63:0] _13084;
    wire [63:0] _13085;
    wire [62:0] _13086;
    wire [63:0] _13088;
    wire _13089;
    wire _13090;
    wire _13078;
    wire [63:0] _13075;
    wire [63:0] _13076;
    wire [62:0] _13077;
    wire [63:0] _13079;
    wire _13080;
    wire _13081;
    wire _13069;
    wire [63:0] _13066;
    wire [63:0] _13067;
    wire [62:0] _13068;
    wire [63:0] _13070;
    wire _13071;
    wire _13072;
    wire _13060;
    wire [63:0] _13057;
    wire [63:0] _13058;
    wire [62:0] _13059;
    wire [63:0] _13061;
    wire _13062;
    wire _13063;
    wire _13051;
    wire [63:0] _13048;
    wire [63:0] _13049;
    wire [62:0] _13050;
    wire [63:0] _13052;
    wire _13053;
    wire _13054;
    wire _13042;
    wire [63:0] _13039;
    wire [63:0] _13040;
    wire [62:0] _13041;
    wire [63:0] _13043;
    wire _13044;
    wire _13045;
    wire _13033;
    wire [63:0] _13030;
    wire [63:0] _13031;
    wire [62:0] _13032;
    wire [63:0] _13034;
    wire _13035;
    wire _13036;
    wire _13024;
    wire [63:0] _13021;
    wire [63:0] _13022;
    wire [62:0] _13023;
    wire [63:0] _13025;
    wire _13026;
    wire _13027;
    wire _13015;
    wire [63:0] _13012;
    wire [63:0] _13013;
    wire [62:0] _13014;
    wire [63:0] _13016;
    wire _13017;
    wire _13018;
    wire _13006;
    wire [63:0] _13003;
    wire [63:0] _13004;
    wire [62:0] _13005;
    wire [63:0] _13007;
    wire _13008;
    wire _13009;
    wire _12997;
    wire [63:0] _12994;
    wire [63:0] _12995;
    wire [62:0] _12996;
    wire [63:0] _12998;
    wire _12999;
    wire _13000;
    wire _12988;
    wire [63:0] _12985;
    wire [63:0] _12986;
    wire [62:0] _12987;
    wire [63:0] _12989;
    wire _12990;
    wire _12991;
    wire _12979;
    wire [63:0] _12976;
    wire [63:0] _12977;
    wire [62:0] _12978;
    wire [63:0] _12980;
    wire _12981;
    wire _12982;
    wire _12970;
    wire [63:0] _12967;
    wire [63:0] _12968;
    wire [62:0] _12969;
    wire [63:0] _12971;
    wire _12972;
    wire _12973;
    wire _12961;
    wire [63:0] _12958;
    wire [63:0] _12959;
    wire [62:0] _12960;
    wire [63:0] _12962;
    wire _12963;
    wire _12964;
    wire _12952;
    wire [63:0] _12949;
    wire [63:0] _12950;
    wire [62:0] _12951;
    wire [63:0] _12953;
    wire _12954;
    wire _12955;
    wire _12943;
    wire [63:0] _12940;
    wire [63:0] _12941;
    wire [62:0] _12942;
    wire [63:0] _12944;
    wire _12945;
    wire _12946;
    wire _12934;
    wire [63:0] _12931;
    wire [63:0] _12932;
    wire [62:0] _12933;
    wire [63:0] _12935;
    wire _12936;
    wire _12937;
    wire _12925;
    wire [63:0] _12922;
    wire [63:0] _12923;
    wire [62:0] _12924;
    wire [63:0] _12926;
    wire _12927;
    wire _12928;
    wire _12916;
    wire [63:0] _12913;
    wire [63:0] _12914;
    wire [62:0] _12915;
    wire [63:0] _12917;
    wire _12918;
    wire _12919;
    wire _12907;
    wire [63:0] _12904;
    wire [63:0] _12905;
    wire [62:0] _12906;
    wire [63:0] _12908;
    wire _12909;
    wire _12910;
    wire _12898;
    wire [63:0] _12895;
    wire [63:0] _12896;
    wire [62:0] _12897;
    wire [63:0] _12899;
    wire _12900;
    wire _12901;
    wire _12889;
    wire [63:0] _12886;
    wire [63:0] _12887;
    wire [62:0] _12888;
    wire [63:0] _12890;
    wire _12891;
    wire _12892;
    wire _12880;
    wire [63:0] _12877;
    wire [63:0] _12878;
    wire [62:0] _12879;
    wire [63:0] _12881;
    wire _12882;
    wire _12883;
    wire _12871;
    wire [63:0] _12868;
    wire [63:0] _12869;
    wire [62:0] _12870;
    wire [63:0] _12872;
    wire _12873;
    wire _12874;
    wire _12862;
    wire [63:0] _12859;
    wire [63:0] _12860;
    wire [62:0] _12861;
    wire [63:0] _12863;
    wire _12864;
    wire _12865;
    wire [63:0] _12852;
    wire _12853;
    wire [63:0] _12854;
    wire _12855;
    wire _12856;
    wire [63:0] _12857;
    wire [62:0] _12858;
    wire [63:0] _12866;
    wire [62:0] _12867;
    wire [63:0] _12875;
    wire [62:0] _12876;
    wire [63:0] _12884;
    wire [62:0] _12885;
    wire [63:0] _12893;
    wire [62:0] _12894;
    wire [63:0] _12902;
    wire [62:0] _12903;
    wire [63:0] _12911;
    wire [62:0] _12912;
    wire [63:0] _12920;
    wire [62:0] _12921;
    wire [63:0] _12929;
    wire [62:0] _12930;
    wire [63:0] _12938;
    wire [62:0] _12939;
    wire [63:0] _12947;
    wire [62:0] _12948;
    wire [63:0] _12956;
    wire [62:0] _12957;
    wire [63:0] _12965;
    wire [62:0] _12966;
    wire [63:0] _12974;
    wire [62:0] _12975;
    wire [63:0] _12983;
    wire [62:0] _12984;
    wire [63:0] _12992;
    wire [62:0] _12993;
    wire [63:0] _13001;
    wire [62:0] _13002;
    wire [63:0] _13010;
    wire [62:0] _13011;
    wire [63:0] _13019;
    wire [62:0] _13020;
    wire [63:0] _13028;
    wire [62:0] _13029;
    wire [63:0] _13037;
    wire [62:0] _13038;
    wire [63:0] _13046;
    wire [62:0] _13047;
    wire [63:0] _13055;
    wire [62:0] _13056;
    wire [63:0] _13064;
    wire [62:0] _13065;
    wire [63:0] _13073;
    wire [62:0] _13074;
    wire [63:0] _13082;
    wire [62:0] _13083;
    wire [63:0] _13091;
    wire [62:0] _13092;
    wire [63:0] _13100;
    wire [62:0] _13101;
    wire [63:0] _13109;
    wire [62:0] _13110;
    wire [63:0] _13118;
    wire [62:0] _13119;
    wire [63:0] _13127;
    wire [62:0] _13128;
    wire [63:0] _13136;
    wire [62:0] _13137;
    wire [63:0] _13145;
    wire [62:0] _13146;
    wire [63:0] _13154;
    wire [62:0] _13155;
    wire [63:0] _13163;
    wire [62:0] _13164;
    wire [63:0] _13172;
    wire [62:0] _13173;
    wire [63:0] _13181;
    wire [62:0] _13182;
    wire [63:0] _13190;
    wire [62:0] _13191;
    wire [63:0] _13199;
    wire [62:0] _13200;
    wire [63:0] _13208;
    wire [62:0] _13209;
    wire [63:0] _13217;
    wire [62:0] _13218;
    wire [63:0] _13226;
    wire [62:0] _13227;
    wire [63:0] _13235;
    wire [62:0] _13236;
    wire [63:0] _13244;
    wire [62:0] _13245;
    wire [63:0] _13253;
    wire [62:0] _13254;
    wire [63:0] _13262;
    wire [62:0] _13263;
    wire [63:0] _13271;
    wire [62:0] _13272;
    wire [63:0] _13280;
    wire [62:0] _13281;
    wire [63:0] _13289;
    wire [62:0] _13290;
    wire [63:0] _13298;
    wire [62:0] _13299;
    wire [63:0] _13307;
    wire [62:0] _13308;
    wire [63:0] _13316;
    wire [62:0] _13317;
    wire [63:0] _13325;
    wire [62:0] _13326;
    wire [63:0] _13334;
    wire [62:0] _13335;
    wire [63:0] _13343;
    wire [62:0] _13344;
    wire [63:0] _13352;
    wire [62:0] _13353;
    wire [63:0] _13361;
    wire [62:0] _13362;
    wire [63:0] _13370;
    wire [62:0] _13371;
    wire [63:0] _13379;
    wire [62:0] _13380;
    wire [63:0] _13388;
    wire [62:0] _13389;
    wire [63:0] _13397;
    wire [62:0] _13398;
    wire [63:0] _13406;
    wire [62:0] _13407;
    wire [63:0] _13415;
    wire [62:0] _13416;
    wire [63:0] _13424;
    wire [63:0] _13426;
    wire [127:0] _13427;
    wire [63:0] _13428;
    wire [63:0] _14010;
    wire _12838;
    wire [63:0] _12835;
    wire [63:0] _12836;
    wire [62:0] _12837;
    wire [63:0] _12839;
    wire _12840;
    wire _12841;
    wire _12829;
    wire [63:0] _12826;
    wire [63:0] _12827;
    wire [62:0] _12828;
    wire [63:0] _12830;
    wire _12831;
    wire _12832;
    wire _12820;
    wire [63:0] _12817;
    wire [63:0] _12818;
    wire [62:0] _12819;
    wire [63:0] _12821;
    wire _12822;
    wire _12823;
    wire _12811;
    wire [63:0] _12808;
    wire [63:0] _12809;
    wire [62:0] _12810;
    wire [63:0] _12812;
    wire _12813;
    wire _12814;
    wire _12802;
    wire [63:0] _12799;
    wire [63:0] _12800;
    wire [62:0] _12801;
    wire [63:0] _12803;
    wire _12804;
    wire _12805;
    wire _12793;
    wire [63:0] _12790;
    wire [63:0] _12791;
    wire [62:0] _12792;
    wire [63:0] _12794;
    wire _12795;
    wire _12796;
    wire _12784;
    wire [63:0] _12781;
    wire [63:0] _12782;
    wire [62:0] _12783;
    wire [63:0] _12785;
    wire _12786;
    wire _12787;
    wire _12775;
    wire [63:0] _12772;
    wire [63:0] _12773;
    wire [62:0] _12774;
    wire [63:0] _12776;
    wire _12777;
    wire _12778;
    wire _12766;
    wire [63:0] _12763;
    wire [63:0] _12764;
    wire [62:0] _12765;
    wire [63:0] _12767;
    wire _12768;
    wire _12769;
    wire _12757;
    wire [63:0] _12754;
    wire [63:0] _12755;
    wire [62:0] _12756;
    wire [63:0] _12758;
    wire _12759;
    wire _12760;
    wire _12748;
    wire [63:0] _12745;
    wire [63:0] _12746;
    wire [62:0] _12747;
    wire [63:0] _12749;
    wire _12750;
    wire _12751;
    wire _12739;
    wire [63:0] _12736;
    wire [63:0] _12737;
    wire [62:0] _12738;
    wire [63:0] _12740;
    wire _12741;
    wire _12742;
    wire _12730;
    wire [63:0] _12727;
    wire [63:0] _12728;
    wire [62:0] _12729;
    wire [63:0] _12731;
    wire _12732;
    wire _12733;
    wire _12721;
    wire [63:0] _12718;
    wire [63:0] _12719;
    wire [62:0] _12720;
    wire [63:0] _12722;
    wire _12723;
    wire _12724;
    wire _12712;
    wire [63:0] _12709;
    wire [63:0] _12710;
    wire [62:0] _12711;
    wire [63:0] _12713;
    wire _12714;
    wire _12715;
    wire _12703;
    wire [63:0] _12700;
    wire [63:0] _12701;
    wire [62:0] _12702;
    wire [63:0] _12704;
    wire _12705;
    wire _12706;
    wire _12694;
    wire [63:0] _12691;
    wire [63:0] _12692;
    wire [62:0] _12693;
    wire [63:0] _12695;
    wire _12696;
    wire _12697;
    wire _12685;
    wire [63:0] _12682;
    wire [63:0] _12683;
    wire [62:0] _12684;
    wire [63:0] _12686;
    wire _12687;
    wire _12688;
    wire _12676;
    wire [63:0] _12673;
    wire [63:0] _12674;
    wire [62:0] _12675;
    wire [63:0] _12677;
    wire _12678;
    wire _12679;
    wire _12667;
    wire [63:0] _12664;
    wire [63:0] _12665;
    wire [62:0] _12666;
    wire [63:0] _12668;
    wire _12669;
    wire _12670;
    wire _12658;
    wire [63:0] _12655;
    wire [63:0] _12656;
    wire [62:0] _12657;
    wire [63:0] _12659;
    wire _12660;
    wire _12661;
    wire _12649;
    wire [63:0] _12646;
    wire [63:0] _12647;
    wire [62:0] _12648;
    wire [63:0] _12650;
    wire _12651;
    wire _12652;
    wire _12640;
    wire [63:0] _12637;
    wire [63:0] _12638;
    wire [62:0] _12639;
    wire [63:0] _12641;
    wire _12642;
    wire _12643;
    wire _12631;
    wire [63:0] _12628;
    wire [63:0] _12629;
    wire [62:0] _12630;
    wire [63:0] _12632;
    wire _12633;
    wire _12634;
    wire _12622;
    wire [63:0] _12619;
    wire [63:0] _12620;
    wire [62:0] _12621;
    wire [63:0] _12623;
    wire _12624;
    wire _12625;
    wire _12613;
    wire [63:0] _12610;
    wire [63:0] _12611;
    wire [62:0] _12612;
    wire [63:0] _12614;
    wire _12615;
    wire _12616;
    wire _12604;
    wire [63:0] _12601;
    wire [63:0] _12602;
    wire [62:0] _12603;
    wire [63:0] _12605;
    wire _12606;
    wire _12607;
    wire _12595;
    wire [63:0] _12592;
    wire [63:0] _12593;
    wire [62:0] _12594;
    wire [63:0] _12596;
    wire _12597;
    wire _12598;
    wire _12586;
    wire [63:0] _12583;
    wire [63:0] _12584;
    wire [62:0] _12585;
    wire [63:0] _12587;
    wire _12588;
    wire _12589;
    wire _12577;
    wire [63:0] _12574;
    wire [63:0] _12575;
    wire [62:0] _12576;
    wire [63:0] _12578;
    wire _12579;
    wire _12580;
    wire _12568;
    wire [63:0] _12565;
    wire [63:0] _12566;
    wire [62:0] _12567;
    wire [63:0] _12569;
    wire _12570;
    wire _12571;
    wire _12559;
    wire [63:0] _12556;
    wire [63:0] _12557;
    wire [62:0] _12558;
    wire [63:0] _12560;
    wire _12561;
    wire _12562;
    wire _12550;
    wire [63:0] _12547;
    wire [63:0] _12548;
    wire [62:0] _12549;
    wire [63:0] _12551;
    wire _12552;
    wire _12553;
    wire _12541;
    wire [63:0] _12538;
    wire [63:0] _12539;
    wire [62:0] _12540;
    wire [63:0] _12542;
    wire _12543;
    wire _12544;
    wire _12532;
    wire [63:0] _12529;
    wire [63:0] _12530;
    wire [62:0] _12531;
    wire [63:0] _12533;
    wire _12534;
    wire _12535;
    wire _12523;
    wire [63:0] _12520;
    wire [63:0] _12521;
    wire [62:0] _12522;
    wire [63:0] _12524;
    wire _12525;
    wire _12526;
    wire _12514;
    wire [63:0] _12511;
    wire [63:0] _12512;
    wire [62:0] _12513;
    wire [63:0] _12515;
    wire _12516;
    wire _12517;
    wire _12505;
    wire [63:0] _12502;
    wire [63:0] _12503;
    wire [62:0] _12504;
    wire [63:0] _12506;
    wire _12507;
    wire _12508;
    wire _12496;
    wire [63:0] _12493;
    wire [63:0] _12494;
    wire [62:0] _12495;
    wire [63:0] _12497;
    wire _12498;
    wire _12499;
    wire _12487;
    wire [63:0] _12484;
    wire [63:0] _12485;
    wire [62:0] _12486;
    wire [63:0] _12488;
    wire _12489;
    wire _12490;
    wire _12478;
    wire [63:0] _12475;
    wire [63:0] _12476;
    wire [62:0] _12477;
    wire [63:0] _12479;
    wire _12480;
    wire _12481;
    wire _12469;
    wire [63:0] _12466;
    wire [63:0] _12467;
    wire [62:0] _12468;
    wire [63:0] _12470;
    wire _12471;
    wire _12472;
    wire _12460;
    wire [63:0] _12457;
    wire [63:0] _12458;
    wire [62:0] _12459;
    wire [63:0] _12461;
    wire _12462;
    wire _12463;
    wire _12451;
    wire [63:0] _12448;
    wire [63:0] _12449;
    wire [62:0] _12450;
    wire [63:0] _12452;
    wire _12453;
    wire _12454;
    wire _12442;
    wire [63:0] _12439;
    wire [63:0] _12440;
    wire [62:0] _12441;
    wire [63:0] _12443;
    wire _12444;
    wire _12445;
    wire _12433;
    wire [63:0] _12430;
    wire [63:0] _12431;
    wire [62:0] _12432;
    wire [63:0] _12434;
    wire _12435;
    wire _12436;
    wire _12424;
    wire [63:0] _12421;
    wire [63:0] _12422;
    wire [62:0] _12423;
    wire [63:0] _12425;
    wire _12426;
    wire _12427;
    wire _12415;
    wire [63:0] _12412;
    wire [63:0] _12413;
    wire [62:0] _12414;
    wire [63:0] _12416;
    wire _12417;
    wire _12418;
    wire _12406;
    wire [63:0] _12403;
    wire [63:0] _12404;
    wire [62:0] _12405;
    wire [63:0] _12407;
    wire _12408;
    wire _12409;
    wire _12397;
    wire [63:0] _12394;
    wire [63:0] _12395;
    wire [62:0] _12396;
    wire [63:0] _12398;
    wire _12399;
    wire _12400;
    wire _12388;
    wire [63:0] _12385;
    wire [63:0] _12386;
    wire [62:0] _12387;
    wire [63:0] _12389;
    wire _12390;
    wire _12391;
    wire _12379;
    wire [63:0] _12376;
    wire [63:0] _12377;
    wire [62:0] _12378;
    wire [63:0] _12380;
    wire _12381;
    wire _12382;
    wire _12370;
    wire [63:0] _12367;
    wire [63:0] _12368;
    wire [62:0] _12369;
    wire [63:0] _12371;
    wire _12372;
    wire _12373;
    wire _12361;
    wire [63:0] _12358;
    wire [63:0] _12359;
    wire [62:0] _12360;
    wire [63:0] _12362;
    wire _12363;
    wire _12364;
    wire _12352;
    wire [63:0] _12349;
    wire [63:0] _12350;
    wire [62:0] _12351;
    wire [63:0] _12353;
    wire _12354;
    wire _12355;
    wire _12343;
    wire [63:0] _12340;
    wire [63:0] _12341;
    wire [62:0] _12342;
    wire [63:0] _12344;
    wire _12345;
    wire _12346;
    wire _12334;
    wire [63:0] _12331;
    wire [63:0] _12332;
    wire [62:0] _12333;
    wire [63:0] _12335;
    wire _12336;
    wire _12337;
    wire _12325;
    wire [63:0] _12322;
    wire [63:0] _12323;
    wire [62:0] _12324;
    wire [63:0] _12326;
    wire _12327;
    wire _12328;
    wire _12316;
    wire [63:0] _12313;
    wire [63:0] _12314;
    wire [62:0] _12315;
    wire [63:0] _12317;
    wire _12318;
    wire _12319;
    wire _12307;
    wire [63:0] _12304;
    wire [63:0] _12305;
    wire [62:0] _12306;
    wire [63:0] _12308;
    wire _12309;
    wire _12310;
    wire _12298;
    wire [63:0] _12295;
    wire [63:0] _12296;
    wire [62:0] _12297;
    wire [63:0] _12299;
    wire _12300;
    wire _12301;
    wire _12289;
    wire [63:0] _12286;
    wire [63:0] _12287;
    wire [62:0] _12288;
    wire [63:0] _12290;
    wire _12291;
    wire _12292;
    wire _12280;
    wire [63:0] _12277;
    wire [63:0] _12278;
    wire [62:0] _12279;
    wire [63:0] _12281;
    wire _12282;
    wire _12283;
    wire [63:0] _12272;
    wire [63:0] _12268;
    wire [63:0] _12269;
    wire _12270;
    wire [63:0] _12271;
    wire _12273;
    wire _12274;
    wire [63:0] _12275;
    wire [62:0] _12276;
    wire [63:0] _12284;
    wire [62:0] _12285;
    wire [63:0] _12293;
    wire [62:0] _12294;
    wire [63:0] _12302;
    wire [62:0] _12303;
    wire [63:0] _12311;
    wire [62:0] _12312;
    wire [63:0] _12320;
    wire [62:0] _12321;
    wire [63:0] _12329;
    wire [62:0] _12330;
    wire [63:0] _12338;
    wire [62:0] _12339;
    wire [63:0] _12347;
    wire [62:0] _12348;
    wire [63:0] _12356;
    wire [62:0] _12357;
    wire [63:0] _12365;
    wire [62:0] _12366;
    wire [63:0] _12374;
    wire [62:0] _12375;
    wire [63:0] _12383;
    wire [62:0] _12384;
    wire [63:0] _12392;
    wire [62:0] _12393;
    wire [63:0] _12401;
    wire [62:0] _12402;
    wire [63:0] _12410;
    wire [62:0] _12411;
    wire [63:0] _12419;
    wire [62:0] _12420;
    wire [63:0] _12428;
    wire [62:0] _12429;
    wire [63:0] _12437;
    wire [62:0] _12438;
    wire [63:0] _12446;
    wire [62:0] _12447;
    wire [63:0] _12455;
    wire [62:0] _12456;
    wire [63:0] _12464;
    wire [62:0] _12465;
    wire [63:0] _12473;
    wire [62:0] _12474;
    wire [63:0] _12482;
    wire [62:0] _12483;
    wire [63:0] _12491;
    wire [62:0] _12492;
    wire [63:0] _12500;
    wire [62:0] _12501;
    wire [63:0] _12509;
    wire [62:0] _12510;
    wire [63:0] _12518;
    wire [62:0] _12519;
    wire [63:0] _12527;
    wire [62:0] _12528;
    wire [63:0] _12536;
    wire [62:0] _12537;
    wire [63:0] _12545;
    wire [62:0] _12546;
    wire [63:0] _12554;
    wire [62:0] _12555;
    wire [63:0] _12563;
    wire [62:0] _12564;
    wire [63:0] _12572;
    wire [62:0] _12573;
    wire [63:0] _12581;
    wire [62:0] _12582;
    wire [63:0] _12590;
    wire [62:0] _12591;
    wire [63:0] _12599;
    wire [62:0] _12600;
    wire [63:0] _12608;
    wire [62:0] _12609;
    wire [63:0] _12617;
    wire [62:0] _12618;
    wire [63:0] _12626;
    wire [62:0] _12627;
    wire [63:0] _12635;
    wire [62:0] _12636;
    wire [63:0] _12644;
    wire [62:0] _12645;
    wire [63:0] _12653;
    wire [62:0] _12654;
    wire [63:0] _12662;
    wire [62:0] _12663;
    wire [63:0] _12671;
    wire [62:0] _12672;
    wire [63:0] _12680;
    wire [62:0] _12681;
    wire [63:0] _12689;
    wire [62:0] _12690;
    wire [63:0] _12698;
    wire [62:0] _12699;
    wire [63:0] _12707;
    wire [62:0] _12708;
    wire [63:0] _12716;
    wire [62:0] _12717;
    wire [63:0] _12725;
    wire [62:0] _12726;
    wire [63:0] _12734;
    wire [62:0] _12735;
    wire [63:0] _12743;
    wire [62:0] _12744;
    wire [63:0] _12752;
    wire [62:0] _12753;
    wire [63:0] _12761;
    wire [62:0] _12762;
    wire [63:0] _12770;
    wire [62:0] _12771;
    wire [63:0] _12779;
    wire [62:0] _12780;
    wire [63:0] _12788;
    wire [62:0] _12789;
    wire [63:0] _12797;
    wire [62:0] _12798;
    wire [63:0] _12806;
    wire [62:0] _12807;
    wire [63:0] _12815;
    wire [62:0] _12816;
    wire [63:0] _12824;
    wire [62:0] _12825;
    wire [63:0] _12833;
    wire [62:0] _12834;
    wire [63:0] _12842;
    wire [127:0] _12843;
    wire [63:0] _12844;
    wire [63:0] _12265;
    wire _12845;
    wire [63:0] _12846;
    wire _12263;
    wire [63:0] _12264;
    wire _12847;
    wire _12848;
    wire [63:0] _14011;
    wire _12252;
    wire [63:0] _12249;
    wire [63:0] _12250;
    wire [62:0] _12251;
    wire [63:0] _12253;
    wire _12254;
    wire _12255;
    wire _12243;
    wire [63:0] _12240;
    wire [63:0] _12241;
    wire [62:0] _12242;
    wire [63:0] _12244;
    wire _12245;
    wire _12246;
    wire _12234;
    wire [63:0] _12231;
    wire [63:0] _12232;
    wire [62:0] _12233;
    wire [63:0] _12235;
    wire _12236;
    wire _12237;
    wire _12225;
    wire [63:0] _12222;
    wire [63:0] _12223;
    wire [62:0] _12224;
    wire [63:0] _12226;
    wire _12227;
    wire _12228;
    wire _12216;
    wire [63:0] _12213;
    wire [63:0] _12214;
    wire [62:0] _12215;
    wire [63:0] _12217;
    wire _12218;
    wire _12219;
    wire _12207;
    wire [63:0] _12204;
    wire [63:0] _12205;
    wire [62:0] _12206;
    wire [63:0] _12208;
    wire _12209;
    wire _12210;
    wire _12198;
    wire [63:0] _12195;
    wire [63:0] _12196;
    wire [62:0] _12197;
    wire [63:0] _12199;
    wire _12200;
    wire _12201;
    wire _12189;
    wire [63:0] _12186;
    wire [63:0] _12187;
    wire [62:0] _12188;
    wire [63:0] _12190;
    wire _12191;
    wire _12192;
    wire _12180;
    wire [63:0] _12177;
    wire [63:0] _12178;
    wire [62:0] _12179;
    wire [63:0] _12181;
    wire _12182;
    wire _12183;
    wire _12171;
    wire [63:0] _12168;
    wire [63:0] _12169;
    wire [62:0] _12170;
    wire [63:0] _12172;
    wire _12173;
    wire _12174;
    wire _12162;
    wire [63:0] _12159;
    wire [63:0] _12160;
    wire [62:0] _12161;
    wire [63:0] _12163;
    wire _12164;
    wire _12165;
    wire _12153;
    wire [63:0] _12150;
    wire [63:0] _12151;
    wire [62:0] _12152;
    wire [63:0] _12154;
    wire _12155;
    wire _12156;
    wire _12144;
    wire [63:0] _12141;
    wire [63:0] _12142;
    wire [62:0] _12143;
    wire [63:0] _12145;
    wire _12146;
    wire _12147;
    wire _12135;
    wire [63:0] _12132;
    wire [63:0] _12133;
    wire [62:0] _12134;
    wire [63:0] _12136;
    wire _12137;
    wire _12138;
    wire _12126;
    wire [63:0] _12123;
    wire [63:0] _12124;
    wire [62:0] _12125;
    wire [63:0] _12127;
    wire _12128;
    wire _12129;
    wire _12117;
    wire [63:0] _12114;
    wire [63:0] _12115;
    wire [62:0] _12116;
    wire [63:0] _12118;
    wire _12119;
    wire _12120;
    wire _12108;
    wire [63:0] _12105;
    wire [63:0] _12106;
    wire [62:0] _12107;
    wire [63:0] _12109;
    wire _12110;
    wire _12111;
    wire _12099;
    wire [63:0] _12096;
    wire [63:0] _12097;
    wire [62:0] _12098;
    wire [63:0] _12100;
    wire _12101;
    wire _12102;
    wire _12090;
    wire [63:0] _12087;
    wire [63:0] _12088;
    wire [62:0] _12089;
    wire [63:0] _12091;
    wire _12092;
    wire _12093;
    wire _12081;
    wire [63:0] _12078;
    wire [63:0] _12079;
    wire [62:0] _12080;
    wire [63:0] _12082;
    wire _12083;
    wire _12084;
    wire _12072;
    wire [63:0] _12069;
    wire [63:0] _12070;
    wire [62:0] _12071;
    wire [63:0] _12073;
    wire _12074;
    wire _12075;
    wire _12063;
    wire [63:0] _12060;
    wire [63:0] _12061;
    wire [62:0] _12062;
    wire [63:0] _12064;
    wire _12065;
    wire _12066;
    wire _12054;
    wire [63:0] _12051;
    wire [63:0] _12052;
    wire [62:0] _12053;
    wire [63:0] _12055;
    wire _12056;
    wire _12057;
    wire _12045;
    wire [63:0] _12042;
    wire [63:0] _12043;
    wire [62:0] _12044;
    wire [63:0] _12046;
    wire _12047;
    wire _12048;
    wire _12036;
    wire [63:0] _12033;
    wire [63:0] _12034;
    wire [62:0] _12035;
    wire [63:0] _12037;
    wire _12038;
    wire _12039;
    wire _12027;
    wire [63:0] _12024;
    wire [63:0] _12025;
    wire [62:0] _12026;
    wire [63:0] _12028;
    wire _12029;
    wire _12030;
    wire _12018;
    wire [63:0] _12015;
    wire [63:0] _12016;
    wire [62:0] _12017;
    wire [63:0] _12019;
    wire _12020;
    wire _12021;
    wire _12009;
    wire [63:0] _12006;
    wire [63:0] _12007;
    wire [62:0] _12008;
    wire [63:0] _12010;
    wire _12011;
    wire _12012;
    wire _12000;
    wire [63:0] _11997;
    wire [63:0] _11998;
    wire [62:0] _11999;
    wire [63:0] _12001;
    wire _12002;
    wire _12003;
    wire _11991;
    wire [63:0] _11988;
    wire [63:0] _11989;
    wire [62:0] _11990;
    wire [63:0] _11992;
    wire _11993;
    wire _11994;
    wire _11982;
    wire [63:0] _11979;
    wire [63:0] _11980;
    wire [62:0] _11981;
    wire [63:0] _11983;
    wire _11984;
    wire _11985;
    wire _11973;
    wire [63:0] _11970;
    wire [63:0] _11971;
    wire [62:0] _11972;
    wire [63:0] _11974;
    wire _11975;
    wire _11976;
    wire _11964;
    wire [63:0] _11961;
    wire [63:0] _11962;
    wire [62:0] _11963;
    wire [63:0] _11965;
    wire _11966;
    wire _11967;
    wire _11955;
    wire [63:0] _11952;
    wire [63:0] _11953;
    wire [62:0] _11954;
    wire [63:0] _11956;
    wire _11957;
    wire _11958;
    wire _11946;
    wire [63:0] _11943;
    wire [63:0] _11944;
    wire [62:0] _11945;
    wire [63:0] _11947;
    wire _11948;
    wire _11949;
    wire _11937;
    wire [63:0] _11934;
    wire [63:0] _11935;
    wire [62:0] _11936;
    wire [63:0] _11938;
    wire _11939;
    wire _11940;
    wire _11928;
    wire [63:0] _11925;
    wire [63:0] _11926;
    wire [62:0] _11927;
    wire [63:0] _11929;
    wire _11930;
    wire _11931;
    wire _11919;
    wire [63:0] _11916;
    wire [63:0] _11917;
    wire [62:0] _11918;
    wire [63:0] _11920;
    wire _11921;
    wire _11922;
    wire _11910;
    wire [63:0] _11907;
    wire [63:0] _11908;
    wire [62:0] _11909;
    wire [63:0] _11911;
    wire _11912;
    wire _11913;
    wire _11901;
    wire [63:0] _11898;
    wire [63:0] _11899;
    wire [62:0] _11900;
    wire [63:0] _11902;
    wire _11903;
    wire _11904;
    wire _11892;
    wire [63:0] _11889;
    wire [63:0] _11890;
    wire [62:0] _11891;
    wire [63:0] _11893;
    wire _11894;
    wire _11895;
    wire _11883;
    wire [63:0] _11880;
    wire [63:0] _11881;
    wire [62:0] _11882;
    wire [63:0] _11884;
    wire _11885;
    wire _11886;
    wire _11874;
    wire [63:0] _11871;
    wire [63:0] _11872;
    wire [62:0] _11873;
    wire [63:0] _11875;
    wire _11876;
    wire _11877;
    wire _11865;
    wire [63:0] _11862;
    wire [63:0] _11863;
    wire [62:0] _11864;
    wire [63:0] _11866;
    wire _11867;
    wire _11868;
    wire _11856;
    wire [63:0] _11853;
    wire [63:0] _11854;
    wire [62:0] _11855;
    wire [63:0] _11857;
    wire _11858;
    wire _11859;
    wire _11847;
    wire [63:0] _11844;
    wire [63:0] _11845;
    wire [62:0] _11846;
    wire [63:0] _11848;
    wire _11849;
    wire _11850;
    wire _11838;
    wire [63:0] _11835;
    wire [63:0] _11836;
    wire [62:0] _11837;
    wire [63:0] _11839;
    wire _11840;
    wire _11841;
    wire _11829;
    wire [63:0] _11826;
    wire [63:0] _11827;
    wire [62:0] _11828;
    wire [63:0] _11830;
    wire _11831;
    wire _11832;
    wire _11820;
    wire [63:0] _11817;
    wire [63:0] _11818;
    wire [62:0] _11819;
    wire [63:0] _11821;
    wire _11822;
    wire _11823;
    wire _11811;
    wire [63:0] _11808;
    wire [63:0] _11809;
    wire [62:0] _11810;
    wire [63:0] _11812;
    wire _11813;
    wire _11814;
    wire _11802;
    wire [63:0] _11799;
    wire [63:0] _11800;
    wire [62:0] _11801;
    wire [63:0] _11803;
    wire _11804;
    wire _11805;
    wire _11793;
    wire [63:0] _11790;
    wire [63:0] _11791;
    wire [62:0] _11792;
    wire [63:0] _11794;
    wire _11795;
    wire _11796;
    wire _11784;
    wire [63:0] _11781;
    wire [63:0] _11782;
    wire [62:0] _11783;
    wire [63:0] _11785;
    wire _11786;
    wire _11787;
    wire _11775;
    wire [63:0] _11772;
    wire [63:0] _11773;
    wire [62:0] _11774;
    wire [63:0] _11776;
    wire _11777;
    wire _11778;
    wire _11766;
    wire [63:0] _11763;
    wire [63:0] _11764;
    wire [62:0] _11765;
    wire [63:0] _11767;
    wire _11768;
    wire _11769;
    wire _11757;
    wire [63:0] _11754;
    wire [63:0] _11755;
    wire [62:0] _11756;
    wire [63:0] _11758;
    wire _11759;
    wire _11760;
    wire _11748;
    wire [63:0] _11745;
    wire [63:0] _11746;
    wire [62:0] _11747;
    wire [63:0] _11749;
    wire _11750;
    wire _11751;
    wire _11739;
    wire [63:0] _11736;
    wire [63:0] _11737;
    wire [62:0] _11738;
    wire [63:0] _11740;
    wire _11741;
    wire _11742;
    wire _11730;
    wire [63:0] _11727;
    wire [63:0] _11728;
    wire [62:0] _11729;
    wire [63:0] _11731;
    wire _11732;
    wire _11733;
    wire _11721;
    wire [63:0] _11718;
    wire [63:0] _11719;
    wire [62:0] _11720;
    wire [63:0] _11722;
    wire _11723;
    wire _11724;
    wire _11712;
    wire [63:0] _11709;
    wire [63:0] _11710;
    wire [62:0] _11711;
    wire [63:0] _11713;
    wire _11714;
    wire _11715;
    wire _11703;
    wire [63:0] _11700;
    wire [63:0] _11701;
    wire [62:0] _11702;
    wire [63:0] _11704;
    wire _11705;
    wire _11706;
    wire _11694;
    wire [63:0] _11691;
    wire [63:0] _11692;
    wire [62:0] _11693;
    wire [63:0] _11695;
    wire _11696;
    wire _11697;
    wire [63:0] _11681;
    wire [127:0] _11682;
    wire [63:0] _11683;
    wire _11684;
    wire [63:0] _11685;
    wire _11687;
    wire _11688;
    wire [63:0] _11689;
    wire [62:0] _11690;
    wire [63:0] _11698;
    wire [62:0] _11699;
    wire [63:0] _11707;
    wire [62:0] _11708;
    wire [63:0] _11716;
    wire [62:0] _11717;
    wire [63:0] _11725;
    wire [62:0] _11726;
    wire [63:0] _11734;
    wire [62:0] _11735;
    wire [63:0] _11743;
    wire [62:0] _11744;
    wire [63:0] _11752;
    wire [62:0] _11753;
    wire [63:0] _11761;
    wire [62:0] _11762;
    wire [63:0] _11770;
    wire [62:0] _11771;
    wire [63:0] _11779;
    wire [62:0] _11780;
    wire [63:0] _11788;
    wire [62:0] _11789;
    wire [63:0] _11797;
    wire [62:0] _11798;
    wire [63:0] _11806;
    wire [62:0] _11807;
    wire [63:0] _11815;
    wire [62:0] _11816;
    wire [63:0] _11824;
    wire [62:0] _11825;
    wire [63:0] _11833;
    wire [62:0] _11834;
    wire [63:0] _11842;
    wire [62:0] _11843;
    wire [63:0] _11851;
    wire [62:0] _11852;
    wire [63:0] _11860;
    wire [62:0] _11861;
    wire [63:0] _11869;
    wire [62:0] _11870;
    wire [63:0] _11878;
    wire [62:0] _11879;
    wire [63:0] _11887;
    wire [62:0] _11888;
    wire [63:0] _11896;
    wire [62:0] _11897;
    wire [63:0] _11905;
    wire [62:0] _11906;
    wire [63:0] _11914;
    wire [62:0] _11915;
    wire [63:0] _11923;
    wire [62:0] _11924;
    wire [63:0] _11932;
    wire [62:0] _11933;
    wire [63:0] _11941;
    wire [62:0] _11942;
    wire [63:0] _11950;
    wire [62:0] _11951;
    wire [63:0] _11959;
    wire [62:0] _11960;
    wire [63:0] _11968;
    wire [62:0] _11969;
    wire [63:0] _11977;
    wire [62:0] _11978;
    wire [63:0] _11986;
    wire [62:0] _11987;
    wire [63:0] _11995;
    wire [62:0] _11996;
    wire [63:0] _12004;
    wire [62:0] _12005;
    wire [63:0] _12013;
    wire [62:0] _12014;
    wire [63:0] _12022;
    wire [62:0] _12023;
    wire [63:0] _12031;
    wire [62:0] _12032;
    wire [63:0] _12040;
    wire [62:0] _12041;
    wire [63:0] _12049;
    wire [62:0] _12050;
    wire [63:0] _12058;
    wire [62:0] _12059;
    wire [63:0] _12067;
    wire [62:0] _12068;
    wire [63:0] _12076;
    wire [62:0] _12077;
    wire [63:0] _12085;
    wire [62:0] _12086;
    wire [63:0] _12094;
    wire [62:0] _12095;
    wire [63:0] _12103;
    wire [62:0] _12104;
    wire [63:0] _12112;
    wire [62:0] _12113;
    wire [63:0] _12121;
    wire [62:0] _12122;
    wire [63:0] _12130;
    wire [62:0] _12131;
    wire [63:0] _12139;
    wire [62:0] _12140;
    wire [63:0] _12148;
    wire [62:0] _12149;
    wire [63:0] _12157;
    wire [62:0] _12158;
    wire [63:0] _12166;
    wire [62:0] _12167;
    wire [63:0] _12175;
    wire [62:0] _12176;
    wire [63:0] _12184;
    wire [62:0] _12185;
    wire [63:0] _12193;
    wire [62:0] _12194;
    wire [63:0] _12202;
    wire [62:0] _12203;
    wire [63:0] _12211;
    wire [62:0] _12212;
    wire [63:0] _12220;
    wire [62:0] _12221;
    wire [63:0] _12229;
    wire [62:0] _12230;
    wire [63:0] _12238;
    wire [62:0] _12239;
    wire [63:0] _12247;
    wire [62:0] _12248;
    wire [63:0] _12256;
    wire [127:0] _12257;
    wire [63:0] _12258;
    wire _11669;
    wire [63:0] _11666;
    wire [63:0] _11667;
    wire [62:0] _11668;
    wire [63:0] _11670;
    wire _11671;
    wire _11672;
    wire _11660;
    wire [63:0] _11657;
    wire [63:0] _11658;
    wire [62:0] _11659;
    wire [63:0] _11661;
    wire _11662;
    wire _11663;
    wire _11651;
    wire [63:0] _11648;
    wire [63:0] _11649;
    wire [62:0] _11650;
    wire [63:0] _11652;
    wire _11653;
    wire _11654;
    wire _11642;
    wire [63:0] _11639;
    wire [63:0] _11640;
    wire [62:0] _11641;
    wire [63:0] _11643;
    wire _11644;
    wire _11645;
    wire _11633;
    wire [63:0] _11630;
    wire [63:0] _11631;
    wire [62:0] _11632;
    wire [63:0] _11634;
    wire _11635;
    wire _11636;
    wire _11624;
    wire [63:0] _11621;
    wire [63:0] _11622;
    wire [62:0] _11623;
    wire [63:0] _11625;
    wire _11626;
    wire _11627;
    wire _11615;
    wire [63:0] _11612;
    wire [63:0] _11613;
    wire [62:0] _11614;
    wire [63:0] _11616;
    wire _11617;
    wire _11618;
    wire _11606;
    wire [63:0] _11603;
    wire [63:0] _11604;
    wire [62:0] _11605;
    wire [63:0] _11607;
    wire _11608;
    wire _11609;
    wire _11597;
    wire [63:0] _11594;
    wire [63:0] _11595;
    wire [62:0] _11596;
    wire [63:0] _11598;
    wire _11599;
    wire _11600;
    wire _11588;
    wire [63:0] _11585;
    wire [63:0] _11586;
    wire [62:0] _11587;
    wire [63:0] _11589;
    wire _11590;
    wire _11591;
    wire _11579;
    wire [63:0] _11576;
    wire [63:0] _11577;
    wire [62:0] _11578;
    wire [63:0] _11580;
    wire _11581;
    wire _11582;
    wire _11570;
    wire [63:0] _11567;
    wire [63:0] _11568;
    wire [62:0] _11569;
    wire [63:0] _11571;
    wire _11572;
    wire _11573;
    wire _11561;
    wire [63:0] _11558;
    wire [63:0] _11559;
    wire [62:0] _11560;
    wire [63:0] _11562;
    wire _11563;
    wire _11564;
    wire _11552;
    wire [63:0] _11549;
    wire [63:0] _11550;
    wire [62:0] _11551;
    wire [63:0] _11553;
    wire _11554;
    wire _11555;
    wire _11543;
    wire [63:0] _11540;
    wire [63:0] _11541;
    wire [62:0] _11542;
    wire [63:0] _11544;
    wire _11545;
    wire _11546;
    wire _11534;
    wire [63:0] _11531;
    wire [63:0] _11532;
    wire [62:0] _11533;
    wire [63:0] _11535;
    wire _11536;
    wire _11537;
    wire _11525;
    wire [63:0] _11522;
    wire [63:0] _11523;
    wire [62:0] _11524;
    wire [63:0] _11526;
    wire _11527;
    wire _11528;
    wire _11516;
    wire [63:0] _11513;
    wire [63:0] _11514;
    wire [62:0] _11515;
    wire [63:0] _11517;
    wire _11518;
    wire _11519;
    wire _11507;
    wire [63:0] _11504;
    wire [63:0] _11505;
    wire [62:0] _11506;
    wire [63:0] _11508;
    wire _11509;
    wire _11510;
    wire _11498;
    wire [63:0] _11495;
    wire [63:0] _11496;
    wire [62:0] _11497;
    wire [63:0] _11499;
    wire _11500;
    wire _11501;
    wire _11489;
    wire [63:0] _11486;
    wire [63:0] _11487;
    wire [62:0] _11488;
    wire [63:0] _11490;
    wire _11491;
    wire _11492;
    wire _11480;
    wire [63:0] _11477;
    wire [63:0] _11478;
    wire [62:0] _11479;
    wire [63:0] _11481;
    wire _11482;
    wire _11483;
    wire _11471;
    wire [63:0] _11468;
    wire [63:0] _11469;
    wire [62:0] _11470;
    wire [63:0] _11472;
    wire _11473;
    wire _11474;
    wire _11462;
    wire [63:0] _11459;
    wire [63:0] _11460;
    wire [62:0] _11461;
    wire [63:0] _11463;
    wire _11464;
    wire _11465;
    wire _11453;
    wire [63:0] _11450;
    wire [63:0] _11451;
    wire [62:0] _11452;
    wire [63:0] _11454;
    wire _11455;
    wire _11456;
    wire _11444;
    wire [63:0] _11441;
    wire [63:0] _11442;
    wire [62:0] _11443;
    wire [63:0] _11445;
    wire _11446;
    wire _11447;
    wire _11435;
    wire [63:0] _11432;
    wire [63:0] _11433;
    wire [62:0] _11434;
    wire [63:0] _11436;
    wire _11437;
    wire _11438;
    wire _11426;
    wire [63:0] _11423;
    wire [63:0] _11424;
    wire [62:0] _11425;
    wire [63:0] _11427;
    wire _11428;
    wire _11429;
    wire _11417;
    wire [63:0] _11414;
    wire [63:0] _11415;
    wire [62:0] _11416;
    wire [63:0] _11418;
    wire _11419;
    wire _11420;
    wire _11408;
    wire [63:0] _11405;
    wire [63:0] _11406;
    wire [62:0] _11407;
    wire [63:0] _11409;
    wire _11410;
    wire _11411;
    wire _11399;
    wire [63:0] _11396;
    wire [63:0] _11397;
    wire [62:0] _11398;
    wire [63:0] _11400;
    wire _11401;
    wire _11402;
    wire _11390;
    wire [63:0] _11387;
    wire [63:0] _11388;
    wire [62:0] _11389;
    wire [63:0] _11391;
    wire _11392;
    wire _11393;
    wire _11381;
    wire [63:0] _11378;
    wire [63:0] _11379;
    wire [62:0] _11380;
    wire [63:0] _11382;
    wire _11383;
    wire _11384;
    wire _11372;
    wire [63:0] _11369;
    wire [63:0] _11370;
    wire [62:0] _11371;
    wire [63:0] _11373;
    wire _11374;
    wire _11375;
    wire _11363;
    wire [63:0] _11360;
    wire [63:0] _11361;
    wire [62:0] _11362;
    wire [63:0] _11364;
    wire _11365;
    wire _11366;
    wire _11354;
    wire [63:0] _11351;
    wire [63:0] _11352;
    wire [62:0] _11353;
    wire [63:0] _11355;
    wire _11356;
    wire _11357;
    wire _11345;
    wire [63:0] _11342;
    wire [63:0] _11343;
    wire [62:0] _11344;
    wire [63:0] _11346;
    wire _11347;
    wire _11348;
    wire _11336;
    wire [63:0] _11333;
    wire [63:0] _11334;
    wire [62:0] _11335;
    wire [63:0] _11337;
    wire _11338;
    wire _11339;
    wire _11327;
    wire [63:0] _11324;
    wire [63:0] _11325;
    wire [62:0] _11326;
    wire [63:0] _11328;
    wire _11329;
    wire _11330;
    wire _11318;
    wire [63:0] _11315;
    wire [63:0] _11316;
    wire [62:0] _11317;
    wire [63:0] _11319;
    wire _11320;
    wire _11321;
    wire _11309;
    wire [63:0] _11306;
    wire [63:0] _11307;
    wire [62:0] _11308;
    wire [63:0] _11310;
    wire _11311;
    wire _11312;
    wire _11300;
    wire [63:0] _11297;
    wire [63:0] _11298;
    wire [62:0] _11299;
    wire [63:0] _11301;
    wire _11302;
    wire _11303;
    wire _11291;
    wire [63:0] _11288;
    wire [63:0] _11289;
    wire [62:0] _11290;
    wire [63:0] _11292;
    wire _11293;
    wire _11294;
    wire _11282;
    wire [63:0] _11279;
    wire [63:0] _11280;
    wire [62:0] _11281;
    wire [63:0] _11283;
    wire _11284;
    wire _11285;
    wire _11273;
    wire [63:0] _11270;
    wire [63:0] _11271;
    wire [62:0] _11272;
    wire [63:0] _11274;
    wire _11275;
    wire _11276;
    wire _11264;
    wire [63:0] _11261;
    wire [63:0] _11262;
    wire [62:0] _11263;
    wire [63:0] _11265;
    wire _11266;
    wire _11267;
    wire _11255;
    wire [63:0] _11252;
    wire [63:0] _11253;
    wire [62:0] _11254;
    wire [63:0] _11256;
    wire _11257;
    wire _11258;
    wire _11246;
    wire [63:0] _11243;
    wire [63:0] _11244;
    wire [62:0] _11245;
    wire [63:0] _11247;
    wire _11248;
    wire _11249;
    wire _11237;
    wire [63:0] _11234;
    wire [63:0] _11235;
    wire [62:0] _11236;
    wire [63:0] _11238;
    wire _11239;
    wire _11240;
    wire _11228;
    wire [63:0] _11225;
    wire [63:0] _11226;
    wire [62:0] _11227;
    wire [63:0] _11229;
    wire _11230;
    wire _11231;
    wire _11219;
    wire [63:0] _11216;
    wire [63:0] _11217;
    wire [62:0] _11218;
    wire [63:0] _11220;
    wire _11221;
    wire _11222;
    wire _11210;
    wire [63:0] _11207;
    wire [63:0] _11208;
    wire [62:0] _11209;
    wire [63:0] _11211;
    wire _11212;
    wire _11213;
    wire _11201;
    wire [63:0] _11198;
    wire [63:0] _11199;
    wire [62:0] _11200;
    wire [63:0] _11202;
    wire _11203;
    wire _11204;
    wire _11192;
    wire [63:0] _11189;
    wire [63:0] _11190;
    wire [62:0] _11191;
    wire [63:0] _11193;
    wire _11194;
    wire _11195;
    wire _11183;
    wire [63:0] _11180;
    wire [63:0] _11181;
    wire [62:0] _11182;
    wire [63:0] _11184;
    wire _11185;
    wire _11186;
    wire _11174;
    wire [63:0] _11171;
    wire [63:0] _11172;
    wire [62:0] _11173;
    wire [63:0] _11175;
    wire _11176;
    wire _11177;
    wire _11165;
    wire [63:0] _11162;
    wire [63:0] _11163;
    wire [62:0] _11164;
    wire [63:0] _11166;
    wire _11167;
    wire _11168;
    wire _11156;
    wire [63:0] _11153;
    wire [63:0] _11154;
    wire [62:0] _11155;
    wire [63:0] _11157;
    wire _11158;
    wire _11159;
    wire _11147;
    wire [63:0] _11144;
    wire [63:0] _11145;
    wire [62:0] _11146;
    wire [63:0] _11148;
    wire _11149;
    wire _11150;
    wire _11138;
    wire [63:0] _11135;
    wire [63:0] _11136;
    wire [62:0] _11137;
    wire [63:0] _11139;
    wire _11140;
    wire _11141;
    wire _11129;
    wire [63:0] _11126;
    wire [63:0] _11127;
    wire [62:0] _11128;
    wire [63:0] _11130;
    wire _11131;
    wire _11132;
    wire _11120;
    wire [63:0] _11117;
    wire [63:0] _11118;
    wire [62:0] _11119;
    wire [63:0] _11121;
    wire _11122;
    wire _11123;
    wire _11111;
    wire [63:0] _11108;
    wire [63:0] _11109;
    wire [62:0] _11110;
    wire [63:0] _11112;
    wire _11113;
    wire _11114;
    wire [63:0] _11101;
    wire _11102;
    wire [63:0] _11103;
    wire _11104;
    wire _11105;
    wire [63:0] _11106;
    wire [62:0] _11107;
    wire [63:0] _11115;
    wire [62:0] _11116;
    wire [63:0] _11124;
    wire [62:0] _11125;
    wire [63:0] _11133;
    wire [62:0] _11134;
    wire [63:0] _11142;
    wire [62:0] _11143;
    wire [63:0] _11151;
    wire [62:0] _11152;
    wire [63:0] _11160;
    wire [62:0] _11161;
    wire [63:0] _11169;
    wire [62:0] _11170;
    wire [63:0] _11178;
    wire [62:0] _11179;
    wire [63:0] _11187;
    wire [62:0] _11188;
    wire [63:0] _11196;
    wire [62:0] _11197;
    wire [63:0] _11205;
    wire [62:0] _11206;
    wire [63:0] _11214;
    wire [62:0] _11215;
    wire [63:0] _11223;
    wire [62:0] _11224;
    wire [63:0] _11232;
    wire [62:0] _11233;
    wire [63:0] _11241;
    wire [62:0] _11242;
    wire [63:0] _11250;
    wire [62:0] _11251;
    wire [63:0] _11259;
    wire [62:0] _11260;
    wire [63:0] _11268;
    wire [62:0] _11269;
    wire [63:0] _11277;
    wire [62:0] _11278;
    wire [63:0] _11286;
    wire [62:0] _11287;
    wire [63:0] _11295;
    wire [62:0] _11296;
    wire [63:0] _11304;
    wire [62:0] _11305;
    wire [63:0] _11313;
    wire [62:0] _11314;
    wire [63:0] _11322;
    wire [62:0] _11323;
    wire [63:0] _11331;
    wire [62:0] _11332;
    wire [63:0] _11340;
    wire [62:0] _11341;
    wire [63:0] _11349;
    wire [62:0] _11350;
    wire [63:0] _11358;
    wire [62:0] _11359;
    wire [63:0] _11367;
    wire [62:0] _11368;
    wire [63:0] _11376;
    wire [62:0] _11377;
    wire [63:0] _11385;
    wire [62:0] _11386;
    wire [63:0] _11394;
    wire [62:0] _11395;
    wire [63:0] _11403;
    wire [62:0] _11404;
    wire [63:0] _11412;
    wire [62:0] _11413;
    wire [63:0] _11421;
    wire [62:0] _11422;
    wire [63:0] _11430;
    wire [62:0] _11431;
    wire [63:0] _11439;
    wire [62:0] _11440;
    wire [63:0] _11448;
    wire [62:0] _11449;
    wire [63:0] _11457;
    wire [62:0] _11458;
    wire [63:0] _11466;
    wire [62:0] _11467;
    wire [63:0] _11475;
    wire [62:0] _11476;
    wire [63:0] _11484;
    wire [62:0] _11485;
    wire [63:0] _11493;
    wire [62:0] _11494;
    wire [63:0] _11502;
    wire [62:0] _11503;
    wire [63:0] _11511;
    wire [62:0] _11512;
    wire [63:0] _11520;
    wire [62:0] _11521;
    wire [63:0] _11529;
    wire [62:0] _11530;
    wire [63:0] _11538;
    wire [62:0] _11539;
    wire [63:0] _11547;
    wire [62:0] _11548;
    wire [63:0] _11556;
    wire [62:0] _11557;
    wire [63:0] _11565;
    wire [62:0] _11566;
    wire [63:0] _11574;
    wire [62:0] _11575;
    wire [63:0] _11583;
    wire [62:0] _11584;
    wire [63:0] _11592;
    wire [62:0] _11593;
    wire [63:0] _11601;
    wire [62:0] _11602;
    wire [63:0] _11610;
    wire [62:0] _11611;
    wire [63:0] _11619;
    wire [62:0] _11620;
    wire [63:0] _11628;
    wire [62:0] _11629;
    wire [63:0] _11637;
    wire [62:0] _11638;
    wire [63:0] _11646;
    wire [62:0] _11647;
    wire [63:0] _11655;
    wire [62:0] _11656;
    wire [63:0] _11664;
    wire [62:0] _11665;
    wire [63:0] _11673;
    wire [63:0] _11675;
    wire [127:0] _11676;
    wire [63:0] _11677;
    wire [63:0] _12259;
    wire _11087;
    wire [63:0] _11084;
    wire [63:0] _11085;
    wire [62:0] _11086;
    wire [63:0] _11088;
    wire _11089;
    wire _11090;
    wire _11078;
    wire [63:0] _11075;
    wire [63:0] _11076;
    wire [62:0] _11077;
    wire [63:0] _11079;
    wire _11080;
    wire _11081;
    wire _11069;
    wire [63:0] _11066;
    wire [63:0] _11067;
    wire [62:0] _11068;
    wire [63:0] _11070;
    wire _11071;
    wire _11072;
    wire _11060;
    wire [63:0] _11057;
    wire [63:0] _11058;
    wire [62:0] _11059;
    wire [63:0] _11061;
    wire _11062;
    wire _11063;
    wire _11051;
    wire [63:0] _11048;
    wire [63:0] _11049;
    wire [62:0] _11050;
    wire [63:0] _11052;
    wire _11053;
    wire _11054;
    wire _11042;
    wire [63:0] _11039;
    wire [63:0] _11040;
    wire [62:0] _11041;
    wire [63:0] _11043;
    wire _11044;
    wire _11045;
    wire _11033;
    wire [63:0] _11030;
    wire [63:0] _11031;
    wire [62:0] _11032;
    wire [63:0] _11034;
    wire _11035;
    wire _11036;
    wire _11024;
    wire [63:0] _11021;
    wire [63:0] _11022;
    wire [62:0] _11023;
    wire [63:0] _11025;
    wire _11026;
    wire _11027;
    wire _11015;
    wire [63:0] _11012;
    wire [63:0] _11013;
    wire [62:0] _11014;
    wire [63:0] _11016;
    wire _11017;
    wire _11018;
    wire _11006;
    wire [63:0] _11003;
    wire [63:0] _11004;
    wire [62:0] _11005;
    wire [63:0] _11007;
    wire _11008;
    wire _11009;
    wire _10997;
    wire [63:0] _10994;
    wire [63:0] _10995;
    wire [62:0] _10996;
    wire [63:0] _10998;
    wire _10999;
    wire _11000;
    wire _10988;
    wire [63:0] _10985;
    wire [63:0] _10986;
    wire [62:0] _10987;
    wire [63:0] _10989;
    wire _10990;
    wire _10991;
    wire _10979;
    wire [63:0] _10976;
    wire [63:0] _10977;
    wire [62:0] _10978;
    wire [63:0] _10980;
    wire _10981;
    wire _10982;
    wire _10970;
    wire [63:0] _10967;
    wire [63:0] _10968;
    wire [62:0] _10969;
    wire [63:0] _10971;
    wire _10972;
    wire _10973;
    wire _10961;
    wire [63:0] _10958;
    wire [63:0] _10959;
    wire [62:0] _10960;
    wire [63:0] _10962;
    wire _10963;
    wire _10964;
    wire _10952;
    wire [63:0] _10949;
    wire [63:0] _10950;
    wire [62:0] _10951;
    wire [63:0] _10953;
    wire _10954;
    wire _10955;
    wire _10943;
    wire [63:0] _10940;
    wire [63:0] _10941;
    wire [62:0] _10942;
    wire [63:0] _10944;
    wire _10945;
    wire _10946;
    wire _10934;
    wire [63:0] _10931;
    wire [63:0] _10932;
    wire [62:0] _10933;
    wire [63:0] _10935;
    wire _10936;
    wire _10937;
    wire _10925;
    wire [63:0] _10922;
    wire [63:0] _10923;
    wire [62:0] _10924;
    wire [63:0] _10926;
    wire _10927;
    wire _10928;
    wire _10916;
    wire [63:0] _10913;
    wire [63:0] _10914;
    wire [62:0] _10915;
    wire [63:0] _10917;
    wire _10918;
    wire _10919;
    wire _10907;
    wire [63:0] _10904;
    wire [63:0] _10905;
    wire [62:0] _10906;
    wire [63:0] _10908;
    wire _10909;
    wire _10910;
    wire _10898;
    wire [63:0] _10895;
    wire [63:0] _10896;
    wire [62:0] _10897;
    wire [63:0] _10899;
    wire _10900;
    wire _10901;
    wire _10889;
    wire [63:0] _10886;
    wire [63:0] _10887;
    wire [62:0] _10888;
    wire [63:0] _10890;
    wire _10891;
    wire _10892;
    wire _10880;
    wire [63:0] _10877;
    wire [63:0] _10878;
    wire [62:0] _10879;
    wire [63:0] _10881;
    wire _10882;
    wire _10883;
    wire _10871;
    wire [63:0] _10868;
    wire [63:0] _10869;
    wire [62:0] _10870;
    wire [63:0] _10872;
    wire _10873;
    wire _10874;
    wire _10862;
    wire [63:0] _10859;
    wire [63:0] _10860;
    wire [62:0] _10861;
    wire [63:0] _10863;
    wire _10864;
    wire _10865;
    wire _10853;
    wire [63:0] _10850;
    wire [63:0] _10851;
    wire [62:0] _10852;
    wire [63:0] _10854;
    wire _10855;
    wire _10856;
    wire _10844;
    wire [63:0] _10841;
    wire [63:0] _10842;
    wire [62:0] _10843;
    wire [63:0] _10845;
    wire _10846;
    wire _10847;
    wire _10835;
    wire [63:0] _10832;
    wire [63:0] _10833;
    wire [62:0] _10834;
    wire [63:0] _10836;
    wire _10837;
    wire _10838;
    wire _10826;
    wire [63:0] _10823;
    wire [63:0] _10824;
    wire [62:0] _10825;
    wire [63:0] _10827;
    wire _10828;
    wire _10829;
    wire _10817;
    wire [63:0] _10814;
    wire [63:0] _10815;
    wire [62:0] _10816;
    wire [63:0] _10818;
    wire _10819;
    wire _10820;
    wire _10808;
    wire [63:0] _10805;
    wire [63:0] _10806;
    wire [62:0] _10807;
    wire [63:0] _10809;
    wire _10810;
    wire _10811;
    wire _10799;
    wire [63:0] _10796;
    wire [63:0] _10797;
    wire [62:0] _10798;
    wire [63:0] _10800;
    wire _10801;
    wire _10802;
    wire _10790;
    wire [63:0] _10787;
    wire [63:0] _10788;
    wire [62:0] _10789;
    wire [63:0] _10791;
    wire _10792;
    wire _10793;
    wire _10781;
    wire [63:0] _10778;
    wire [63:0] _10779;
    wire [62:0] _10780;
    wire [63:0] _10782;
    wire _10783;
    wire _10784;
    wire _10772;
    wire [63:0] _10769;
    wire [63:0] _10770;
    wire [62:0] _10771;
    wire [63:0] _10773;
    wire _10774;
    wire _10775;
    wire _10763;
    wire [63:0] _10760;
    wire [63:0] _10761;
    wire [62:0] _10762;
    wire [63:0] _10764;
    wire _10765;
    wire _10766;
    wire _10754;
    wire [63:0] _10751;
    wire [63:0] _10752;
    wire [62:0] _10753;
    wire [63:0] _10755;
    wire _10756;
    wire _10757;
    wire _10745;
    wire [63:0] _10742;
    wire [63:0] _10743;
    wire [62:0] _10744;
    wire [63:0] _10746;
    wire _10747;
    wire _10748;
    wire _10736;
    wire [63:0] _10733;
    wire [63:0] _10734;
    wire [62:0] _10735;
    wire [63:0] _10737;
    wire _10738;
    wire _10739;
    wire _10727;
    wire [63:0] _10724;
    wire [63:0] _10725;
    wire [62:0] _10726;
    wire [63:0] _10728;
    wire _10729;
    wire _10730;
    wire _10718;
    wire [63:0] _10715;
    wire [63:0] _10716;
    wire [62:0] _10717;
    wire [63:0] _10719;
    wire _10720;
    wire _10721;
    wire _10709;
    wire [63:0] _10706;
    wire [63:0] _10707;
    wire [62:0] _10708;
    wire [63:0] _10710;
    wire _10711;
    wire _10712;
    wire _10700;
    wire [63:0] _10697;
    wire [63:0] _10698;
    wire [62:0] _10699;
    wire [63:0] _10701;
    wire _10702;
    wire _10703;
    wire _10691;
    wire [63:0] _10688;
    wire [63:0] _10689;
    wire [62:0] _10690;
    wire [63:0] _10692;
    wire _10693;
    wire _10694;
    wire _10682;
    wire [63:0] _10679;
    wire [63:0] _10680;
    wire [62:0] _10681;
    wire [63:0] _10683;
    wire _10684;
    wire _10685;
    wire _10673;
    wire [63:0] _10670;
    wire [63:0] _10671;
    wire [62:0] _10672;
    wire [63:0] _10674;
    wire _10675;
    wire _10676;
    wire _10664;
    wire [63:0] _10661;
    wire [63:0] _10662;
    wire [62:0] _10663;
    wire [63:0] _10665;
    wire _10666;
    wire _10667;
    wire _10655;
    wire [63:0] _10652;
    wire [63:0] _10653;
    wire [62:0] _10654;
    wire [63:0] _10656;
    wire _10657;
    wire _10658;
    wire _10646;
    wire [63:0] _10643;
    wire [63:0] _10644;
    wire [62:0] _10645;
    wire [63:0] _10647;
    wire _10648;
    wire _10649;
    wire _10637;
    wire [63:0] _10634;
    wire [63:0] _10635;
    wire [62:0] _10636;
    wire [63:0] _10638;
    wire _10639;
    wire _10640;
    wire _10628;
    wire [63:0] _10625;
    wire [63:0] _10626;
    wire [62:0] _10627;
    wire [63:0] _10629;
    wire _10630;
    wire _10631;
    wire _10619;
    wire [63:0] _10616;
    wire [63:0] _10617;
    wire [62:0] _10618;
    wire [63:0] _10620;
    wire _10621;
    wire _10622;
    wire _10610;
    wire [63:0] _10607;
    wire [63:0] _10608;
    wire [62:0] _10609;
    wire [63:0] _10611;
    wire _10612;
    wire _10613;
    wire _10601;
    wire [63:0] _10598;
    wire [63:0] _10599;
    wire [62:0] _10600;
    wire [63:0] _10602;
    wire _10603;
    wire _10604;
    wire _10592;
    wire [63:0] _10589;
    wire [63:0] _10590;
    wire [62:0] _10591;
    wire [63:0] _10593;
    wire _10594;
    wire _10595;
    wire _10583;
    wire [63:0] _10580;
    wire [63:0] _10581;
    wire [62:0] _10582;
    wire [63:0] _10584;
    wire _10585;
    wire _10586;
    wire _10574;
    wire [63:0] _10571;
    wire [63:0] _10572;
    wire [62:0] _10573;
    wire [63:0] _10575;
    wire _10576;
    wire _10577;
    wire _10565;
    wire [63:0] _10562;
    wire [63:0] _10563;
    wire [62:0] _10564;
    wire [63:0] _10566;
    wire _10567;
    wire _10568;
    wire _10556;
    wire [63:0] _10553;
    wire [63:0] _10554;
    wire [62:0] _10555;
    wire [63:0] _10557;
    wire _10558;
    wire _10559;
    wire _10547;
    wire [63:0] _10544;
    wire [63:0] _10545;
    wire [62:0] _10546;
    wire [63:0] _10548;
    wire _10549;
    wire _10550;
    wire _10538;
    wire [63:0] _10535;
    wire [63:0] _10536;
    wire [62:0] _10537;
    wire [63:0] _10539;
    wire _10540;
    wire _10541;
    wire _10529;
    wire [63:0] _10526;
    wire [63:0] _10527;
    wire [62:0] _10528;
    wire [63:0] _10530;
    wire _10531;
    wire _10532;
    wire [63:0] _10521;
    wire [63:0] _10517;
    wire [63:0] _10518;
    wire _10519;
    wire [63:0] _10520;
    wire _10522;
    wire _10523;
    wire [63:0] _10524;
    wire [62:0] _10525;
    wire [63:0] _10533;
    wire [62:0] _10534;
    wire [63:0] _10542;
    wire [62:0] _10543;
    wire [63:0] _10551;
    wire [62:0] _10552;
    wire [63:0] _10560;
    wire [62:0] _10561;
    wire [63:0] _10569;
    wire [62:0] _10570;
    wire [63:0] _10578;
    wire [62:0] _10579;
    wire [63:0] _10587;
    wire [62:0] _10588;
    wire [63:0] _10596;
    wire [62:0] _10597;
    wire [63:0] _10605;
    wire [62:0] _10606;
    wire [63:0] _10614;
    wire [62:0] _10615;
    wire [63:0] _10623;
    wire [62:0] _10624;
    wire [63:0] _10632;
    wire [62:0] _10633;
    wire [63:0] _10641;
    wire [62:0] _10642;
    wire [63:0] _10650;
    wire [62:0] _10651;
    wire [63:0] _10659;
    wire [62:0] _10660;
    wire [63:0] _10668;
    wire [62:0] _10669;
    wire [63:0] _10677;
    wire [62:0] _10678;
    wire [63:0] _10686;
    wire [62:0] _10687;
    wire [63:0] _10695;
    wire [62:0] _10696;
    wire [63:0] _10704;
    wire [62:0] _10705;
    wire [63:0] _10713;
    wire [62:0] _10714;
    wire [63:0] _10722;
    wire [62:0] _10723;
    wire [63:0] _10731;
    wire [62:0] _10732;
    wire [63:0] _10740;
    wire [62:0] _10741;
    wire [63:0] _10749;
    wire [62:0] _10750;
    wire [63:0] _10758;
    wire [62:0] _10759;
    wire [63:0] _10767;
    wire [62:0] _10768;
    wire [63:0] _10776;
    wire [62:0] _10777;
    wire [63:0] _10785;
    wire [62:0] _10786;
    wire [63:0] _10794;
    wire [62:0] _10795;
    wire [63:0] _10803;
    wire [62:0] _10804;
    wire [63:0] _10812;
    wire [62:0] _10813;
    wire [63:0] _10821;
    wire [62:0] _10822;
    wire [63:0] _10830;
    wire [62:0] _10831;
    wire [63:0] _10839;
    wire [62:0] _10840;
    wire [63:0] _10848;
    wire [62:0] _10849;
    wire [63:0] _10857;
    wire [62:0] _10858;
    wire [63:0] _10866;
    wire [62:0] _10867;
    wire [63:0] _10875;
    wire [62:0] _10876;
    wire [63:0] _10884;
    wire [62:0] _10885;
    wire [63:0] _10893;
    wire [62:0] _10894;
    wire [63:0] _10902;
    wire [62:0] _10903;
    wire [63:0] _10911;
    wire [62:0] _10912;
    wire [63:0] _10920;
    wire [62:0] _10921;
    wire [63:0] _10929;
    wire [62:0] _10930;
    wire [63:0] _10938;
    wire [62:0] _10939;
    wire [63:0] _10947;
    wire [62:0] _10948;
    wire [63:0] _10956;
    wire [62:0] _10957;
    wire [63:0] _10965;
    wire [62:0] _10966;
    wire [63:0] _10974;
    wire [62:0] _10975;
    wire [63:0] _10983;
    wire [62:0] _10984;
    wire [63:0] _10992;
    wire [62:0] _10993;
    wire [63:0] _11001;
    wire [62:0] _11002;
    wire [63:0] _11010;
    wire [62:0] _11011;
    wire [63:0] _11019;
    wire [62:0] _11020;
    wire [63:0] _11028;
    wire [62:0] _11029;
    wire [63:0] _11037;
    wire [62:0] _11038;
    wire [63:0] _11046;
    wire [62:0] _11047;
    wire [63:0] _11055;
    wire [62:0] _11056;
    wire [63:0] _11064;
    wire [62:0] _11065;
    wire [63:0] _11073;
    wire [62:0] _11074;
    wire [63:0] _11082;
    wire [62:0] _11083;
    wire [63:0] _11091;
    wire [127:0] _11092;
    wire [63:0] _11093;
    wire _11094;
    wire [63:0] _11095;
    wire [63:0] _10511;
    wire _10512;
    wire [63:0] _10513;
    wire _11096;
    wire _11097;
    wire [63:0] _12260;
    wire _10502;
    wire [63:0] _10499;
    wire [63:0] _10500;
    wire [62:0] _10501;
    wire [63:0] _10503;
    wire _10504;
    wire _10505;
    wire _10493;
    wire [63:0] _10490;
    wire [63:0] _10491;
    wire [62:0] _10492;
    wire [63:0] _10494;
    wire _10495;
    wire _10496;
    wire _10484;
    wire [63:0] _10481;
    wire [63:0] _10482;
    wire [62:0] _10483;
    wire [63:0] _10485;
    wire _10486;
    wire _10487;
    wire _10475;
    wire [63:0] _10472;
    wire [63:0] _10473;
    wire [62:0] _10474;
    wire [63:0] _10476;
    wire _10477;
    wire _10478;
    wire _10466;
    wire [63:0] _10463;
    wire [63:0] _10464;
    wire [62:0] _10465;
    wire [63:0] _10467;
    wire _10468;
    wire _10469;
    wire _10457;
    wire [63:0] _10454;
    wire [63:0] _10455;
    wire [62:0] _10456;
    wire [63:0] _10458;
    wire _10459;
    wire _10460;
    wire _10448;
    wire [63:0] _10445;
    wire [63:0] _10446;
    wire [62:0] _10447;
    wire [63:0] _10449;
    wire _10450;
    wire _10451;
    wire _10439;
    wire [63:0] _10436;
    wire [63:0] _10437;
    wire [62:0] _10438;
    wire [63:0] _10440;
    wire _10441;
    wire _10442;
    wire _10430;
    wire [63:0] _10427;
    wire [63:0] _10428;
    wire [62:0] _10429;
    wire [63:0] _10431;
    wire _10432;
    wire _10433;
    wire _10421;
    wire [63:0] _10418;
    wire [63:0] _10419;
    wire [62:0] _10420;
    wire [63:0] _10422;
    wire _10423;
    wire _10424;
    wire _10412;
    wire [63:0] _10409;
    wire [63:0] _10410;
    wire [62:0] _10411;
    wire [63:0] _10413;
    wire _10414;
    wire _10415;
    wire _10403;
    wire [63:0] _10400;
    wire [63:0] _10401;
    wire [62:0] _10402;
    wire [63:0] _10404;
    wire _10405;
    wire _10406;
    wire _10394;
    wire [63:0] _10391;
    wire [63:0] _10392;
    wire [62:0] _10393;
    wire [63:0] _10395;
    wire _10396;
    wire _10397;
    wire _10385;
    wire [63:0] _10382;
    wire [63:0] _10383;
    wire [62:0] _10384;
    wire [63:0] _10386;
    wire _10387;
    wire _10388;
    wire _10376;
    wire [63:0] _10373;
    wire [63:0] _10374;
    wire [62:0] _10375;
    wire [63:0] _10377;
    wire _10378;
    wire _10379;
    wire _10367;
    wire [63:0] _10364;
    wire [63:0] _10365;
    wire [62:0] _10366;
    wire [63:0] _10368;
    wire _10369;
    wire _10370;
    wire _10358;
    wire [63:0] _10355;
    wire [63:0] _10356;
    wire [62:0] _10357;
    wire [63:0] _10359;
    wire _10360;
    wire _10361;
    wire _10349;
    wire [63:0] _10346;
    wire [63:0] _10347;
    wire [62:0] _10348;
    wire [63:0] _10350;
    wire _10351;
    wire _10352;
    wire _10340;
    wire [63:0] _10337;
    wire [63:0] _10338;
    wire [62:0] _10339;
    wire [63:0] _10341;
    wire _10342;
    wire _10343;
    wire _10331;
    wire [63:0] _10328;
    wire [63:0] _10329;
    wire [62:0] _10330;
    wire [63:0] _10332;
    wire _10333;
    wire _10334;
    wire _10322;
    wire [63:0] _10319;
    wire [63:0] _10320;
    wire [62:0] _10321;
    wire [63:0] _10323;
    wire _10324;
    wire _10325;
    wire _10313;
    wire [63:0] _10310;
    wire [63:0] _10311;
    wire [62:0] _10312;
    wire [63:0] _10314;
    wire _10315;
    wire _10316;
    wire _10304;
    wire [63:0] _10301;
    wire [63:0] _10302;
    wire [62:0] _10303;
    wire [63:0] _10305;
    wire _10306;
    wire _10307;
    wire _10295;
    wire [63:0] _10292;
    wire [63:0] _10293;
    wire [62:0] _10294;
    wire [63:0] _10296;
    wire _10297;
    wire _10298;
    wire _10286;
    wire [63:0] _10283;
    wire [63:0] _10284;
    wire [62:0] _10285;
    wire [63:0] _10287;
    wire _10288;
    wire _10289;
    wire _10277;
    wire [63:0] _10274;
    wire [63:0] _10275;
    wire [62:0] _10276;
    wire [63:0] _10278;
    wire _10279;
    wire _10280;
    wire _10268;
    wire [63:0] _10265;
    wire [63:0] _10266;
    wire [62:0] _10267;
    wire [63:0] _10269;
    wire _10270;
    wire _10271;
    wire _10259;
    wire [63:0] _10256;
    wire [63:0] _10257;
    wire [62:0] _10258;
    wire [63:0] _10260;
    wire _10261;
    wire _10262;
    wire _10250;
    wire [63:0] _10247;
    wire [63:0] _10248;
    wire [62:0] _10249;
    wire [63:0] _10251;
    wire _10252;
    wire _10253;
    wire _10241;
    wire [63:0] _10238;
    wire [63:0] _10239;
    wire [62:0] _10240;
    wire [63:0] _10242;
    wire _10243;
    wire _10244;
    wire _10232;
    wire [63:0] _10229;
    wire [63:0] _10230;
    wire [62:0] _10231;
    wire [63:0] _10233;
    wire _10234;
    wire _10235;
    wire _10223;
    wire [63:0] _10220;
    wire [63:0] _10221;
    wire [62:0] _10222;
    wire [63:0] _10224;
    wire _10225;
    wire _10226;
    wire _10214;
    wire [63:0] _10211;
    wire [63:0] _10212;
    wire [62:0] _10213;
    wire [63:0] _10215;
    wire _10216;
    wire _10217;
    wire _10205;
    wire [63:0] _10202;
    wire [63:0] _10203;
    wire [62:0] _10204;
    wire [63:0] _10206;
    wire _10207;
    wire _10208;
    wire _10196;
    wire [63:0] _10193;
    wire [63:0] _10194;
    wire [62:0] _10195;
    wire [63:0] _10197;
    wire _10198;
    wire _10199;
    wire _10187;
    wire [63:0] _10184;
    wire [63:0] _10185;
    wire [62:0] _10186;
    wire [63:0] _10188;
    wire _10189;
    wire _10190;
    wire _10178;
    wire [63:0] _10175;
    wire [63:0] _10176;
    wire [62:0] _10177;
    wire [63:0] _10179;
    wire _10180;
    wire _10181;
    wire _10169;
    wire [63:0] _10166;
    wire [63:0] _10167;
    wire [62:0] _10168;
    wire [63:0] _10170;
    wire _10171;
    wire _10172;
    wire _10160;
    wire [63:0] _10157;
    wire [63:0] _10158;
    wire [62:0] _10159;
    wire [63:0] _10161;
    wire _10162;
    wire _10163;
    wire _10151;
    wire [63:0] _10148;
    wire [63:0] _10149;
    wire [62:0] _10150;
    wire [63:0] _10152;
    wire _10153;
    wire _10154;
    wire _10142;
    wire [63:0] _10139;
    wire [63:0] _10140;
    wire [62:0] _10141;
    wire [63:0] _10143;
    wire _10144;
    wire _10145;
    wire _10133;
    wire [63:0] _10130;
    wire [63:0] _10131;
    wire [62:0] _10132;
    wire [63:0] _10134;
    wire _10135;
    wire _10136;
    wire _10124;
    wire [63:0] _10121;
    wire [63:0] _10122;
    wire [62:0] _10123;
    wire [63:0] _10125;
    wire _10126;
    wire _10127;
    wire _10115;
    wire [63:0] _10112;
    wire [63:0] _10113;
    wire [62:0] _10114;
    wire [63:0] _10116;
    wire _10117;
    wire _10118;
    wire _10106;
    wire [63:0] _10103;
    wire [63:0] _10104;
    wire [62:0] _10105;
    wire [63:0] _10107;
    wire _10108;
    wire _10109;
    wire _10097;
    wire [63:0] _10094;
    wire [63:0] _10095;
    wire [62:0] _10096;
    wire [63:0] _10098;
    wire _10099;
    wire _10100;
    wire _10088;
    wire [63:0] _10085;
    wire [63:0] _10086;
    wire [62:0] _10087;
    wire [63:0] _10089;
    wire _10090;
    wire _10091;
    wire _10079;
    wire [63:0] _10076;
    wire [63:0] _10077;
    wire [62:0] _10078;
    wire [63:0] _10080;
    wire _10081;
    wire _10082;
    wire _10070;
    wire [63:0] _10067;
    wire [63:0] _10068;
    wire [62:0] _10069;
    wire [63:0] _10071;
    wire _10072;
    wire _10073;
    wire _10061;
    wire [63:0] _10058;
    wire [63:0] _10059;
    wire [62:0] _10060;
    wire [63:0] _10062;
    wire _10063;
    wire _10064;
    wire _10052;
    wire [63:0] _10049;
    wire [63:0] _10050;
    wire [62:0] _10051;
    wire [63:0] _10053;
    wire _10054;
    wire _10055;
    wire _10043;
    wire [63:0] _10040;
    wire [63:0] _10041;
    wire [62:0] _10042;
    wire [63:0] _10044;
    wire _10045;
    wire _10046;
    wire _10034;
    wire [63:0] _10031;
    wire [63:0] _10032;
    wire [62:0] _10033;
    wire [63:0] _10035;
    wire _10036;
    wire _10037;
    wire _10025;
    wire [63:0] _10022;
    wire [63:0] _10023;
    wire [62:0] _10024;
    wire [63:0] _10026;
    wire _10027;
    wire _10028;
    wire _10016;
    wire [63:0] _10013;
    wire [63:0] _10014;
    wire [62:0] _10015;
    wire [63:0] _10017;
    wire _10018;
    wire _10019;
    wire _10007;
    wire [63:0] _10004;
    wire [63:0] _10005;
    wire [62:0] _10006;
    wire [63:0] _10008;
    wire _10009;
    wire _10010;
    wire _9998;
    wire [63:0] _9995;
    wire [63:0] _9996;
    wire [62:0] _9997;
    wire [63:0] _9999;
    wire _10000;
    wire _10001;
    wire _9989;
    wire [63:0] _9986;
    wire [63:0] _9987;
    wire [62:0] _9988;
    wire [63:0] _9990;
    wire _9991;
    wire _9992;
    wire _9980;
    wire [63:0] _9977;
    wire [63:0] _9978;
    wire [62:0] _9979;
    wire [63:0] _9981;
    wire _9982;
    wire _9983;
    wire _9971;
    wire [63:0] _9968;
    wire [63:0] _9969;
    wire [62:0] _9970;
    wire [63:0] _9972;
    wire _9973;
    wire _9974;
    wire _9962;
    wire [63:0] _9959;
    wire [63:0] _9960;
    wire [62:0] _9961;
    wire [63:0] _9963;
    wire _9964;
    wire _9965;
    wire _9953;
    wire [63:0] _9950;
    wire [63:0] _9951;
    wire [62:0] _9952;
    wire [63:0] _9954;
    wire _9955;
    wire _9956;
    wire _9944;
    wire [63:0] _9941;
    wire [63:0] _9942;
    wire [62:0] _9943;
    wire [63:0] _9945;
    wire _9946;
    wire _9947;
    wire [63:0] _9931;
    wire [127:0] _9932;
    wire [63:0] _9933;
    wire _9934;
    wire [63:0] _9935;
    wire _9937;
    wire _9938;
    wire [63:0] _9939;
    wire [62:0] _9940;
    wire [63:0] _9948;
    wire [62:0] _9949;
    wire [63:0] _9957;
    wire [62:0] _9958;
    wire [63:0] _9966;
    wire [62:0] _9967;
    wire [63:0] _9975;
    wire [62:0] _9976;
    wire [63:0] _9984;
    wire [62:0] _9985;
    wire [63:0] _9993;
    wire [62:0] _9994;
    wire [63:0] _10002;
    wire [62:0] _10003;
    wire [63:0] _10011;
    wire [62:0] _10012;
    wire [63:0] _10020;
    wire [62:0] _10021;
    wire [63:0] _10029;
    wire [62:0] _10030;
    wire [63:0] _10038;
    wire [62:0] _10039;
    wire [63:0] _10047;
    wire [62:0] _10048;
    wire [63:0] _10056;
    wire [62:0] _10057;
    wire [63:0] _10065;
    wire [62:0] _10066;
    wire [63:0] _10074;
    wire [62:0] _10075;
    wire [63:0] _10083;
    wire [62:0] _10084;
    wire [63:0] _10092;
    wire [62:0] _10093;
    wire [63:0] _10101;
    wire [62:0] _10102;
    wire [63:0] _10110;
    wire [62:0] _10111;
    wire [63:0] _10119;
    wire [62:0] _10120;
    wire [63:0] _10128;
    wire [62:0] _10129;
    wire [63:0] _10137;
    wire [62:0] _10138;
    wire [63:0] _10146;
    wire [62:0] _10147;
    wire [63:0] _10155;
    wire [62:0] _10156;
    wire [63:0] _10164;
    wire [62:0] _10165;
    wire [63:0] _10173;
    wire [62:0] _10174;
    wire [63:0] _10182;
    wire [62:0] _10183;
    wire [63:0] _10191;
    wire [62:0] _10192;
    wire [63:0] _10200;
    wire [62:0] _10201;
    wire [63:0] _10209;
    wire [62:0] _10210;
    wire [63:0] _10218;
    wire [62:0] _10219;
    wire [63:0] _10227;
    wire [62:0] _10228;
    wire [63:0] _10236;
    wire [62:0] _10237;
    wire [63:0] _10245;
    wire [62:0] _10246;
    wire [63:0] _10254;
    wire [62:0] _10255;
    wire [63:0] _10263;
    wire [62:0] _10264;
    wire [63:0] _10272;
    wire [62:0] _10273;
    wire [63:0] _10281;
    wire [62:0] _10282;
    wire [63:0] _10290;
    wire [62:0] _10291;
    wire [63:0] _10299;
    wire [62:0] _10300;
    wire [63:0] _10308;
    wire [62:0] _10309;
    wire [63:0] _10317;
    wire [62:0] _10318;
    wire [63:0] _10326;
    wire [62:0] _10327;
    wire [63:0] _10335;
    wire [62:0] _10336;
    wire [63:0] _10344;
    wire [62:0] _10345;
    wire [63:0] _10353;
    wire [62:0] _10354;
    wire [63:0] _10362;
    wire [62:0] _10363;
    wire [63:0] _10371;
    wire [62:0] _10372;
    wire [63:0] _10380;
    wire [62:0] _10381;
    wire [63:0] _10389;
    wire [62:0] _10390;
    wire [63:0] _10398;
    wire [62:0] _10399;
    wire [63:0] _10407;
    wire [62:0] _10408;
    wire [63:0] _10416;
    wire [62:0] _10417;
    wire [63:0] _10425;
    wire [62:0] _10426;
    wire [63:0] _10434;
    wire [62:0] _10435;
    wire [63:0] _10443;
    wire [62:0] _10444;
    wire [63:0] _10452;
    wire [62:0] _10453;
    wire [63:0] _10461;
    wire [62:0] _10462;
    wire [63:0] _10470;
    wire [62:0] _10471;
    wire [63:0] _10479;
    wire [62:0] _10480;
    wire [63:0] _10488;
    wire [62:0] _10489;
    wire [63:0] _10497;
    wire [62:0] _10498;
    wire [63:0] _10506;
    wire [127:0] _10507;
    wire [63:0] _10508;
    wire _9919;
    wire [63:0] _9916;
    wire [63:0] _9917;
    wire [62:0] _9918;
    wire [63:0] _9920;
    wire _9921;
    wire _9922;
    wire _9910;
    wire [63:0] _9907;
    wire [63:0] _9908;
    wire [62:0] _9909;
    wire [63:0] _9911;
    wire _9912;
    wire _9913;
    wire _9901;
    wire [63:0] _9898;
    wire [63:0] _9899;
    wire [62:0] _9900;
    wire [63:0] _9902;
    wire _9903;
    wire _9904;
    wire _9892;
    wire [63:0] _9889;
    wire [63:0] _9890;
    wire [62:0] _9891;
    wire [63:0] _9893;
    wire _9894;
    wire _9895;
    wire _9883;
    wire [63:0] _9880;
    wire [63:0] _9881;
    wire [62:0] _9882;
    wire [63:0] _9884;
    wire _9885;
    wire _9886;
    wire _9874;
    wire [63:0] _9871;
    wire [63:0] _9872;
    wire [62:0] _9873;
    wire [63:0] _9875;
    wire _9876;
    wire _9877;
    wire _9865;
    wire [63:0] _9862;
    wire [63:0] _9863;
    wire [62:0] _9864;
    wire [63:0] _9866;
    wire _9867;
    wire _9868;
    wire _9856;
    wire [63:0] _9853;
    wire [63:0] _9854;
    wire [62:0] _9855;
    wire [63:0] _9857;
    wire _9858;
    wire _9859;
    wire _9847;
    wire [63:0] _9844;
    wire [63:0] _9845;
    wire [62:0] _9846;
    wire [63:0] _9848;
    wire _9849;
    wire _9850;
    wire _9838;
    wire [63:0] _9835;
    wire [63:0] _9836;
    wire [62:0] _9837;
    wire [63:0] _9839;
    wire _9840;
    wire _9841;
    wire _9829;
    wire [63:0] _9826;
    wire [63:0] _9827;
    wire [62:0] _9828;
    wire [63:0] _9830;
    wire _9831;
    wire _9832;
    wire _9820;
    wire [63:0] _9817;
    wire [63:0] _9818;
    wire [62:0] _9819;
    wire [63:0] _9821;
    wire _9822;
    wire _9823;
    wire _9811;
    wire [63:0] _9808;
    wire [63:0] _9809;
    wire [62:0] _9810;
    wire [63:0] _9812;
    wire _9813;
    wire _9814;
    wire _9802;
    wire [63:0] _9799;
    wire [63:0] _9800;
    wire [62:0] _9801;
    wire [63:0] _9803;
    wire _9804;
    wire _9805;
    wire _9793;
    wire [63:0] _9790;
    wire [63:0] _9791;
    wire [62:0] _9792;
    wire [63:0] _9794;
    wire _9795;
    wire _9796;
    wire _9784;
    wire [63:0] _9781;
    wire [63:0] _9782;
    wire [62:0] _9783;
    wire [63:0] _9785;
    wire _9786;
    wire _9787;
    wire _9775;
    wire [63:0] _9772;
    wire [63:0] _9773;
    wire [62:0] _9774;
    wire [63:0] _9776;
    wire _9777;
    wire _9778;
    wire _9766;
    wire [63:0] _9763;
    wire [63:0] _9764;
    wire [62:0] _9765;
    wire [63:0] _9767;
    wire _9768;
    wire _9769;
    wire _9757;
    wire [63:0] _9754;
    wire [63:0] _9755;
    wire [62:0] _9756;
    wire [63:0] _9758;
    wire _9759;
    wire _9760;
    wire _9748;
    wire [63:0] _9745;
    wire [63:0] _9746;
    wire [62:0] _9747;
    wire [63:0] _9749;
    wire _9750;
    wire _9751;
    wire _9739;
    wire [63:0] _9736;
    wire [63:0] _9737;
    wire [62:0] _9738;
    wire [63:0] _9740;
    wire _9741;
    wire _9742;
    wire _9730;
    wire [63:0] _9727;
    wire [63:0] _9728;
    wire [62:0] _9729;
    wire [63:0] _9731;
    wire _9732;
    wire _9733;
    wire _9721;
    wire [63:0] _9718;
    wire [63:0] _9719;
    wire [62:0] _9720;
    wire [63:0] _9722;
    wire _9723;
    wire _9724;
    wire _9712;
    wire [63:0] _9709;
    wire [63:0] _9710;
    wire [62:0] _9711;
    wire [63:0] _9713;
    wire _9714;
    wire _9715;
    wire _9703;
    wire [63:0] _9700;
    wire [63:0] _9701;
    wire [62:0] _9702;
    wire [63:0] _9704;
    wire _9705;
    wire _9706;
    wire _9694;
    wire [63:0] _9691;
    wire [63:0] _9692;
    wire [62:0] _9693;
    wire [63:0] _9695;
    wire _9696;
    wire _9697;
    wire _9685;
    wire [63:0] _9682;
    wire [63:0] _9683;
    wire [62:0] _9684;
    wire [63:0] _9686;
    wire _9687;
    wire _9688;
    wire _9676;
    wire [63:0] _9673;
    wire [63:0] _9674;
    wire [62:0] _9675;
    wire [63:0] _9677;
    wire _9678;
    wire _9679;
    wire _9667;
    wire [63:0] _9664;
    wire [63:0] _9665;
    wire [62:0] _9666;
    wire [63:0] _9668;
    wire _9669;
    wire _9670;
    wire _9658;
    wire [63:0] _9655;
    wire [63:0] _9656;
    wire [62:0] _9657;
    wire [63:0] _9659;
    wire _9660;
    wire _9661;
    wire _9649;
    wire [63:0] _9646;
    wire [63:0] _9647;
    wire [62:0] _9648;
    wire [63:0] _9650;
    wire _9651;
    wire _9652;
    wire _9640;
    wire [63:0] _9637;
    wire [63:0] _9638;
    wire [62:0] _9639;
    wire [63:0] _9641;
    wire _9642;
    wire _9643;
    wire _9631;
    wire [63:0] _9628;
    wire [63:0] _9629;
    wire [62:0] _9630;
    wire [63:0] _9632;
    wire _9633;
    wire _9634;
    wire _9622;
    wire [63:0] _9619;
    wire [63:0] _9620;
    wire [62:0] _9621;
    wire [63:0] _9623;
    wire _9624;
    wire _9625;
    wire _9613;
    wire [63:0] _9610;
    wire [63:0] _9611;
    wire [62:0] _9612;
    wire [63:0] _9614;
    wire _9615;
    wire _9616;
    wire _9604;
    wire [63:0] _9601;
    wire [63:0] _9602;
    wire [62:0] _9603;
    wire [63:0] _9605;
    wire _9606;
    wire _9607;
    wire _9595;
    wire [63:0] _9592;
    wire [63:0] _9593;
    wire [62:0] _9594;
    wire [63:0] _9596;
    wire _9597;
    wire _9598;
    wire _9586;
    wire [63:0] _9583;
    wire [63:0] _9584;
    wire [62:0] _9585;
    wire [63:0] _9587;
    wire _9588;
    wire _9589;
    wire _9577;
    wire [63:0] _9574;
    wire [63:0] _9575;
    wire [62:0] _9576;
    wire [63:0] _9578;
    wire _9579;
    wire _9580;
    wire _9568;
    wire [63:0] _9565;
    wire [63:0] _9566;
    wire [62:0] _9567;
    wire [63:0] _9569;
    wire _9570;
    wire _9571;
    wire _9559;
    wire [63:0] _9556;
    wire [63:0] _9557;
    wire [62:0] _9558;
    wire [63:0] _9560;
    wire _9561;
    wire _9562;
    wire _9550;
    wire [63:0] _9547;
    wire [63:0] _9548;
    wire [62:0] _9549;
    wire [63:0] _9551;
    wire _9552;
    wire _9553;
    wire _9541;
    wire [63:0] _9538;
    wire [63:0] _9539;
    wire [62:0] _9540;
    wire [63:0] _9542;
    wire _9543;
    wire _9544;
    wire _9532;
    wire [63:0] _9529;
    wire [63:0] _9530;
    wire [62:0] _9531;
    wire [63:0] _9533;
    wire _9534;
    wire _9535;
    wire _9523;
    wire [63:0] _9520;
    wire [63:0] _9521;
    wire [62:0] _9522;
    wire [63:0] _9524;
    wire _9525;
    wire _9526;
    wire _9514;
    wire [63:0] _9511;
    wire [63:0] _9512;
    wire [62:0] _9513;
    wire [63:0] _9515;
    wire _9516;
    wire _9517;
    wire _9505;
    wire [63:0] _9502;
    wire [63:0] _9503;
    wire [62:0] _9504;
    wire [63:0] _9506;
    wire _9507;
    wire _9508;
    wire _9496;
    wire [63:0] _9493;
    wire [63:0] _9494;
    wire [62:0] _9495;
    wire [63:0] _9497;
    wire _9498;
    wire _9499;
    wire _9487;
    wire [63:0] _9484;
    wire [63:0] _9485;
    wire [62:0] _9486;
    wire [63:0] _9488;
    wire _9489;
    wire _9490;
    wire _9478;
    wire [63:0] _9475;
    wire [63:0] _9476;
    wire [62:0] _9477;
    wire [63:0] _9479;
    wire _9480;
    wire _9481;
    wire _9469;
    wire [63:0] _9466;
    wire [63:0] _9467;
    wire [62:0] _9468;
    wire [63:0] _9470;
    wire _9471;
    wire _9472;
    wire _9460;
    wire [63:0] _9457;
    wire [63:0] _9458;
    wire [62:0] _9459;
    wire [63:0] _9461;
    wire _9462;
    wire _9463;
    wire _9451;
    wire [63:0] _9448;
    wire [63:0] _9449;
    wire [62:0] _9450;
    wire [63:0] _9452;
    wire _9453;
    wire _9454;
    wire _9442;
    wire [63:0] _9439;
    wire [63:0] _9440;
    wire [62:0] _9441;
    wire [63:0] _9443;
    wire _9444;
    wire _9445;
    wire _9433;
    wire [63:0] _9430;
    wire [63:0] _9431;
    wire [62:0] _9432;
    wire [63:0] _9434;
    wire _9435;
    wire _9436;
    wire _9424;
    wire [63:0] _9421;
    wire [63:0] _9422;
    wire [62:0] _9423;
    wire [63:0] _9425;
    wire _9426;
    wire _9427;
    wire _9415;
    wire [63:0] _9412;
    wire [63:0] _9413;
    wire [62:0] _9414;
    wire [63:0] _9416;
    wire _9417;
    wire _9418;
    wire _9406;
    wire [63:0] _9403;
    wire [63:0] _9404;
    wire [62:0] _9405;
    wire [63:0] _9407;
    wire _9408;
    wire _9409;
    wire _9397;
    wire [63:0] _9394;
    wire [63:0] _9395;
    wire [62:0] _9396;
    wire [63:0] _9398;
    wire _9399;
    wire _9400;
    wire _9388;
    wire [63:0] _9385;
    wire [63:0] _9386;
    wire [62:0] _9387;
    wire [63:0] _9389;
    wire _9390;
    wire _9391;
    wire _9379;
    wire [63:0] _9376;
    wire [63:0] _9377;
    wire [62:0] _9378;
    wire [63:0] _9380;
    wire _9381;
    wire _9382;
    wire _9370;
    wire [63:0] _9367;
    wire [63:0] _9368;
    wire [62:0] _9369;
    wire [63:0] _9371;
    wire _9372;
    wire _9373;
    wire _9361;
    wire [63:0] _9358;
    wire [63:0] _9359;
    wire [62:0] _9360;
    wire [63:0] _9362;
    wire _9363;
    wire _9364;
    wire [63:0] _9351;
    wire _9352;
    wire [63:0] _9353;
    wire _9354;
    wire _9355;
    wire [63:0] _9356;
    wire [62:0] _9357;
    wire [63:0] _9365;
    wire [62:0] _9366;
    wire [63:0] _9374;
    wire [62:0] _9375;
    wire [63:0] _9383;
    wire [62:0] _9384;
    wire [63:0] _9392;
    wire [62:0] _9393;
    wire [63:0] _9401;
    wire [62:0] _9402;
    wire [63:0] _9410;
    wire [62:0] _9411;
    wire [63:0] _9419;
    wire [62:0] _9420;
    wire [63:0] _9428;
    wire [62:0] _9429;
    wire [63:0] _9437;
    wire [62:0] _9438;
    wire [63:0] _9446;
    wire [62:0] _9447;
    wire [63:0] _9455;
    wire [62:0] _9456;
    wire [63:0] _9464;
    wire [62:0] _9465;
    wire [63:0] _9473;
    wire [62:0] _9474;
    wire [63:0] _9482;
    wire [62:0] _9483;
    wire [63:0] _9491;
    wire [62:0] _9492;
    wire [63:0] _9500;
    wire [62:0] _9501;
    wire [63:0] _9509;
    wire [62:0] _9510;
    wire [63:0] _9518;
    wire [62:0] _9519;
    wire [63:0] _9527;
    wire [62:0] _9528;
    wire [63:0] _9536;
    wire [62:0] _9537;
    wire [63:0] _9545;
    wire [62:0] _9546;
    wire [63:0] _9554;
    wire [62:0] _9555;
    wire [63:0] _9563;
    wire [62:0] _9564;
    wire [63:0] _9572;
    wire [62:0] _9573;
    wire [63:0] _9581;
    wire [62:0] _9582;
    wire [63:0] _9590;
    wire [62:0] _9591;
    wire [63:0] _9599;
    wire [62:0] _9600;
    wire [63:0] _9608;
    wire [62:0] _9609;
    wire [63:0] _9617;
    wire [62:0] _9618;
    wire [63:0] _9626;
    wire [62:0] _9627;
    wire [63:0] _9635;
    wire [62:0] _9636;
    wire [63:0] _9644;
    wire [62:0] _9645;
    wire [63:0] _9653;
    wire [62:0] _9654;
    wire [63:0] _9662;
    wire [62:0] _9663;
    wire [63:0] _9671;
    wire [62:0] _9672;
    wire [63:0] _9680;
    wire [62:0] _9681;
    wire [63:0] _9689;
    wire [62:0] _9690;
    wire [63:0] _9698;
    wire [62:0] _9699;
    wire [63:0] _9707;
    wire [62:0] _9708;
    wire [63:0] _9716;
    wire [62:0] _9717;
    wire [63:0] _9725;
    wire [62:0] _9726;
    wire [63:0] _9734;
    wire [62:0] _9735;
    wire [63:0] _9743;
    wire [62:0] _9744;
    wire [63:0] _9752;
    wire [62:0] _9753;
    wire [63:0] _9761;
    wire [62:0] _9762;
    wire [63:0] _9770;
    wire [62:0] _9771;
    wire [63:0] _9779;
    wire [62:0] _9780;
    wire [63:0] _9788;
    wire [62:0] _9789;
    wire [63:0] _9797;
    wire [62:0] _9798;
    wire [63:0] _9806;
    wire [62:0] _9807;
    wire [63:0] _9815;
    wire [62:0] _9816;
    wire [63:0] _9824;
    wire [62:0] _9825;
    wire [63:0] _9833;
    wire [62:0] _9834;
    wire [63:0] _9842;
    wire [62:0] _9843;
    wire [63:0] _9851;
    wire [62:0] _9852;
    wire [63:0] _9860;
    wire [62:0] _9861;
    wire [63:0] _9869;
    wire [62:0] _9870;
    wire [63:0] _9878;
    wire [62:0] _9879;
    wire [63:0] _9887;
    wire [62:0] _9888;
    wire [63:0] _9896;
    wire [62:0] _9897;
    wire [63:0] _9905;
    wire [62:0] _9906;
    wire [63:0] _9914;
    wire [62:0] _9915;
    wire [63:0] _9923;
    wire [63:0] _9925;
    wire [127:0] _9926;
    wire [63:0] _9927;
    wire [63:0] _10509;
    wire _9337;
    wire [63:0] _9334;
    wire [63:0] _9335;
    wire [62:0] _9336;
    wire [63:0] _9338;
    wire _9339;
    wire _9340;
    wire _9328;
    wire [63:0] _9325;
    wire [63:0] _9326;
    wire [62:0] _9327;
    wire [63:0] _9329;
    wire _9330;
    wire _9331;
    wire _9319;
    wire [63:0] _9316;
    wire [63:0] _9317;
    wire [62:0] _9318;
    wire [63:0] _9320;
    wire _9321;
    wire _9322;
    wire _9310;
    wire [63:0] _9307;
    wire [63:0] _9308;
    wire [62:0] _9309;
    wire [63:0] _9311;
    wire _9312;
    wire _9313;
    wire _9301;
    wire [63:0] _9298;
    wire [63:0] _9299;
    wire [62:0] _9300;
    wire [63:0] _9302;
    wire _9303;
    wire _9304;
    wire _9292;
    wire [63:0] _9289;
    wire [63:0] _9290;
    wire [62:0] _9291;
    wire [63:0] _9293;
    wire _9294;
    wire _9295;
    wire _9283;
    wire [63:0] _9280;
    wire [63:0] _9281;
    wire [62:0] _9282;
    wire [63:0] _9284;
    wire _9285;
    wire _9286;
    wire _9274;
    wire [63:0] _9271;
    wire [63:0] _9272;
    wire [62:0] _9273;
    wire [63:0] _9275;
    wire _9276;
    wire _9277;
    wire _9265;
    wire [63:0] _9262;
    wire [63:0] _9263;
    wire [62:0] _9264;
    wire [63:0] _9266;
    wire _9267;
    wire _9268;
    wire _9256;
    wire [63:0] _9253;
    wire [63:0] _9254;
    wire [62:0] _9255;
    wire [63:0] _9257;
    wire _9258;
    wire _9259;
    wire _9247;
    wire [63:0] _9244;
    wire [63:0] _9245;
    wire [62:0] _9246;
    wire [63:0] _9248;
    wire _9249;
    wire _9250;
    wire _9238;
    wire [63:0] _9235;
    wire [63:0] _9236;
    wire [62:0] _9237;
    wire [63:0] _9239;
    wire _9240;
    wire _9241;
    wire _9229;
    wire [63:0] _9226;
    wire [63:0] _9227;
    wire [62:0] _9228;
    wire [63:0] _9230;
    wire _9231;
    wire _9232;
    wire _9220;
    wire [63:0] _9217;
    wire [63:0] _9218;
    wire [62:0] _9219;
    wire [63:0] _9221;
    wire _9222;
    wire _9223;
    wire _9211;
    wire [63:0] _9208;
    wire [63:0] _9209;
    wire [62:0] _9210;
    wire [63:0] _9212;
    wire _9213;
    wire _9214;
    wire _9202;
    wire [63:0] _9199;
    wire [63:0] _9200;
    wire [62:0] _9201;
    wire [63:0] _9203;
    wire _9204;
    wire _9205;
    wire _9193;
    wire [63:0] _9190;
    wire [63:0] _9191;
    wire [62:0] _9192;
    wire [63:0] _9194;
    wire _9195;
    wire _9196;
    wire _9184;
    wire [63:0] _9181;
    wire [63:0] _9182;
    wire [62:0] _9183;
    wire [63:0] _9185;
    wire _9186;
    wire _9187;
    wire _9175;
    wire [63:0] _9172;
    wire [63:0] _9173;
    wire [62:0] _9174;
    wire [63:0] _9176;
    wire _9177;
    wire _9178;
    wire _9166;
    wire [63:0] _9163;
    wire [63:0] _9164;
    wire [62:0] _9165;
    wire [63:0] _9167;
    wire _9168;
    wire _9169;
    wire _9157;
    wire [63:0] _9154;
    wire [63:0] _9155;
    wire [62:0] _9156;
    wire [63:0] _9158;
    wire _9159;
    wire _9160;
    wire _9148;
    wire [63:0] _9145;
    wire [63:0] _9146;
    wire [62:0] _9147;
    wire [63:0] _9149;
    wire _9150;
    wire _9151;
    wire _9139;
    wire [63:0] _9136;
    wire [63:0] _9137;
    wire [62:0] _9138;
    wire [63:0] _9140;
    wire _9141;
    wire _9142;
    wire _9130;
    wire [63:0] _9127;
    wire [63:0] _9128;
    wire [62:0] _9129;
    wire [63:0] _9131;
    wire _9132;
    wire _9133;
    wire _9121;
    wire [63:0] _9118;
    wire [63:0] _9119;
    wire [62:0] _9120;
    wire [63:0] _9122;
    wire _9123;
    wire _9124;
    wire _9112;
    wire [63:0] _9109;
    wire [63:0] _9110;
    wire [62:0] _9111;
    wire [63:0] _9113;
    wire _9114;
    wire _9115;
    wire _9103;
    wire [63:0] _9100;
    wire [63:0] _9101;
    wire [62:0] _9102;
    wire [63:0] _9104;
    wire _9105;
    wire _9106;
    wire _9094;
    wire [63:0] _9091;
    wire [63:0] _9092;
    wire [62:0] _9093;
    wire [63:0] _9095;
    wire _9096;
    wire _9097;
    wire _9085;
    wire [63:0] _9082;
    wire [63:0] _9083;
    wire [62:0] _9084;
    wire [63:0] _9086;
    wire _9087;
    wire _9088;
    wire _9076;
    wire [63:0] _9073;
    wire [63:0] _9074;
    wire [62:0] _9075;
    wire [63:0] _9077;
    wire _9078;
    wire _9079;
    wire _9067;
    wire [63:0] _9064;
    wire [63:0] _9065;
    wire [62:0] _9066;
    wire [63:0] _9068;
    wire _9069;
    wire _9070;
    wire _9058;
    wire [63:0] _9055;
    wire [63:0] _9056;
    wire [62:0] _9057;
    wire [63:0] _9059;
    wire _9060;
    wire _9061;
    wire _9049;
    wire [63:0] _9046;
    wire [63:0] _9047;
    wire [62:0] _9048;
    wire [63:0] _9050;
    wire _9051;
    wire _9052;
    wire _9040;
    wire [63:0] _9037;
    wire [63:0] _9038;
    wire [62:0] _9039;
    wire [63:0] _9041;
    wire _9042;
    wire _9043;
    wire _9031;
    wire [63:0] _9028;
    wire [63:0] _9029;
    wire [62:0] _9030;
    wire [63:0] _9032;
    wire _9033;
    wire _9034;
    wire _9022;
    wire [63:0] _9019;
    wire [63:0] _9020;
    wire [62:0] _9021;
    wire [63:0] _9023;
    wire _9024;
    wire _9025;
    wire _9013;
    wire [63:0] _9010;
    wire [63:0] _9011;
    wire [62:0] _9012;
    wire [63:0] _9014;
    wire _9015;
    wire _9016;
    wire _9004;
    wire [63:0] _9001;
    wire [63:0] _9002;
    wire [62:0] _9003;
    wire [63:0] _9005;
    wire _9006;
    wire _9007;
    wire _8995;
    wire [63:0] _8992;
    wire [63:0] _8993;
    wire [62:0] _8994;
    wire [63:0] _8996;
    wire _8997;
    wire _8998;
    wire _8986;
    wire [63:0] _8983;
    wire [63:0] _8984;
    wire [62:0] _8985;
    wire [63:0] _8987;
    wire _8988;
    wire _8989;
    wire _8977;
    wire [63:0] _8974;
    wire [63:0] _8975;
    wire [62:0] _8976;
    wire [63:0] _8978;
    wire _8979;
    wire _8980;
    wire _8968;
    wire [63:0] _8965;
    wire [63:0] _8966;
    wire [62:0] _8967;
    wire [63:0] _8969;
    wire _8970;
    wire _8971;
    wire _8959;
    wire [63:0] _8956;
    wire [63:0] _8957;
    wire [62:0] _8958;
    wire [63:0] _8960;
    wire _8961;
    wire _8962;
    wire _8950;
    wire [63:0] _8947;
    wire [63:0] _8948;
    wire [62:0] _8949;
    wire [63:0] _8951;
    wire _8952;
    wire _8953;
    wire _8941;
    wire [63:0] _8938;
    wire [63:0] _8939;
    wire [62:0] _8940;
    wire [63:0] _8942;
    wire _8943;
    wire _8944;
    wire _8932;
    wire [63:0] _8929;
    wire [63:0] _8930;
    wire [62:0] _8931;
    wire [63:0] _8933;
    wire _8934;
    wire _8935;
    wire _8923;
    wire [63:0] _8920;
    wire [63:0] _8921;
    wire [62:0] _8922;
    wire [63:0] _8924;
    wire _8925;
    wire _8926;
    wire _8914;
    wire [63:0] _8911;
    wire [63:0] _8912;
    wire [62:0] _8913;
    wire [63:0] _8915;
    wire _8916;
    wire _8917;
    wire _8905;
    wire [63:0] _8902;
    wire [63:0] _8903;
    wire [62:0] _8904;
    wire [63:0] _8906;
    wire _8907;
    wire _8908;
    wire _8896;
    wire [63:0] _8893;
    wire [63:0] _8894;
    wire [62:0] _8895;
    wire [63:0] _8897;
    wire _8898;
    wire _8899;
    wire _8887;
    wire [63:0] _8884;
    wire [63:0] _8885;
    wire [62:0] _8886;
    wire [63:0] _8888;
    wire _8889;
    wire _8890;
    wire _8878;
    wire [63:0] _8875;
    wire [63:0] _8876;
    wire [62:0] _8877;
    wire [63:0] _8879;
    wire _8880;
    wire _8881;
    wire _8869;
    wire [63:0] _8866;
    wire [63:0] _8867;
    wire [62:0] _8868;
    wire [63:0] _8870;
    wire _8871;
    wire _8872;
    wire _8860;
    wire [63:0] _8857;
    wire [63:0] _8858;
    wire [62:0] _8859;
    wire [63:0] _8861;
    wire _8862;
    wire _8863;
    wire _8851;
    wire [63:0] _8848;
    wire [63:0] _8849;
    wire [62:0] _8850;
    wire [63:0] _8852;
    wire _8853;
    wire _8854;
    wire _8842;
    wire [63:0] _8839;
    wire [63:0] _8840;
    wire [62:0] _8841;
    wire [63:0] _8843;
    wire _8844;
    wire _8845;
    wire _8833;
    wire [63:0] _8830;
    wire [63:0] _8831;
    wire [62:0] _8832;
    wire [63:0] _8834;
    wire _8835;
    wire _8836;
    wire _8824;
    wire [63:0] _8821;
    wire [63:0] _8822;
    wire [62:0] _8823;
    wire [63:0] _8825;
    wire _8826;
    wire _8827;
    wire _8815;
    wire [63:0] _8812;
    wire [63:0] _8813;
    wire [62:0] _8814;
    wire [63:0] _8816;
    wire _8817;
    wire _8818;
    wire _8806;
    wire [63:0] _8803;
    wire [63:0] _8804;
    wire [62:0] _8805;
    wire [63:0] _8807;
    wire _8808;
    wire _8809;
    wire _8797;
    wire [63:0] _8794;
    wire [63:0] _8795;
    wire [62:0] _8796;
    wire [63:0] _8798;
    wire _8799;
    wire _8800;
    wire _8788;
    wire [63:0] _8785;
    wire [63:0] _8786;
    wire [62:0] _8787;
    wire [63:0] _8789;
    wire _8790;
    wire _8791;
    wire _8779;
    wire [63:0] _8776;
    wire [63:0] _8777;
    wire [62:0] _8778;
    wire [63:0] _8780;
    wire _8781;
    wire _8782;
    wire [63:0] _8771;
    wire [63:0] _8767;
    wire [63:0] _8768;
    wire _8769;
    wire [63:0] _8770;
    wire _8772;
    wire _8773;
    wire [63:0] _8774;
    wire [62:0] _8775;
    wire [63:0] _8783;
    wire [62:0] _8784;
    wire [63:0] _8792;
    wire [62:0] _8793;
    wire [63:0] _8801;
    wire [62:0] _8802;
    wire [63:0] _8810;
    wire [62:0] _8811;
    wire [63:0] _8819;
    wire [62:0] _8820;
    wire [63:0] _8828;
    wire [62:0] _8829;
    wire [63:0] _8837;
    wire [62:0] _8838;
    wire [63:0] _8846;
    wire [62:0] _8847;
    wire [63:0] _8855;
    wire [62:0] _8856;
    wire [63:0] _8864;
    wire [62:0] _8865;
    wire [63:0] _8873;
    wire [62:0] _8874;
    wire [63:0] _8882;
    wire [62:0] _8883;
    wire [63:0] _8891;
    wire [62:0] _8892;
    wire [63:0] _8900;
    wire [62:0] _8901;
    wire [63:0] _8909;
    wire [62:0] _8910;
    wire [63:0] _8918;
    wire [62:0] _8919;
    wire [63:0] _8927;
    wire [62:0] _8928;
    wire [63:0] _8936;
    wire [62:0] _8937;
    wire [63:0] _8945;
    wire [62:0] _8946;
    wire [63:0] _8954;
    wire [62:0] _8955;
    wire [63:0] _8963;
    wire [62:0] _8964;
    wire [63:0] _8972;
    wire [62:0] _8973;
    wire [63:0] _8981;
    wire [62:0] _8982;
    wire [63:0] _8990;
    wire [62:0] _8991;
    wire [63:0] _8999;
    wire [62:0] _9000;
    wire [63:0] _9008;
    wire [62:0] _9009;
    wire [63:0] _9017;
    wire [62:0] _9018;
    wire [63:0] _9026;
    wire [62:0] _9027;
    wire [63:0] _9035;
    wire [62:0] _9036;
    wire [63:0] _9044;
    wire [62:0] _9045;
    wire [63:0] _9053;
    wire [62:0] _9054;
    wire [63:0] _9062;
    wire [62:0] _9063;
    wire [63:0] _9071;
    wire [62:0] _9072;
    wire [63:0] _9080;
    wire [62:0] _9081;
    wire [63:0] _9089;
    wire [62:0] _9090;
    wire [63:0] _9098;
    wire [62:0] _9099;
    wire [63:0] _9107;
    wire [62:0] _9108;
    wire [63:0] _9116;
    wire [62:0] _9117;
    wire [63:0] _9125;
    wire [62:0] _9126;
    wire [63:0] _9134;
    wire [62:0] _9135;
    wire [63:0] _9143;
    wire [62:0] _9144;
    wire [63:0] _9152;
    wire [62:0] _9153;
    wire [63:0] _9161;
    wire [62:0] _9162;
    wire [63:0] _9170;
    wire [62:0] _9171;
    wire [63:0] _9179;
    wire [62:0] _9180;
    wire [63:0] _9188;
    wire [62:0] _9189;
    wire [63:0] _9197;
    wire [62:0] _9198;
    wire [63:0] _9206;
    wire [62:0] _9207;
    wire [63:0] _9215;
    wire [62:0] _9216;
    wire [63:0] _9224;
    wire [62:0] _9225;
    wire [63:0] _9233;
    wire [62:0] _9234;
    wire [63:0] _9242;
    wire [62:0] _9243;
    wire [63:0] _9251;
    wire [62:0] _9252;
    wire [63:0] _9260;
    wire [62:0] _9261;
    wire [63:0] _9269;
    wire [62:0] _9270;
    wire [63:0] _9278;
    wire [62:0] _9279;
    wire [63:0] _9287;
    wire [62:0] _9288;
    wire [63:0] _9296;
    wire [62:0] _9297;
    wire [63:0] _9305;
    wire [62:0] _9306;
    wire [63:0] _9314;
    wire [62:0] _9315;
    wire [63:0] _9323;
    wire [62:0] _9324;
    wire [63:0] _9332;
    wire [62:0] _9333;
    wire [63:0] _9341;
    wire [127:0] _9342;
    wire [63:0] _9343;
    wire _9344;
    wire [63:0] _9345;
    wire [63:0] _8761;
    wire _8762;
    wire [63:0] _8763;
    wire _9346;
    wire _9347;
    wire [63:0] _10510;
    wire [63:0] _12261;
    wire [63:0] _14012;
    wire [63:0] _15763;
    wire [63:0] _17514;
    wire [63:0] _19265;
    wire [63:0] _19266;
    wire [63:0] _22768;
    wire _8751;
    wire [63:0] _8748;
    wire [63:0] _8749;
    wire [62:0] _8750;
    wire [63:0] _8752;
    wire _8753;
    wire _8754;
    wire _8742;
    wire [63:0] _8739;
    wire [63:0] _8740;
    wire [62:0] _8741;
    wire [63:0] _8743;
    wire _8744;
    wire _8745;
    wire _8733;
    wire [63:0] _8730;
    wire [63:0] _8731;
    wire [62:0] _8732;
    wire [63:0] _8734;
    wire _8735;
    wire _8736;
    wire _8724;
    wire [63:0] _8721;
    wire [63:0] _8722;
    wire [62:0] _8723;
    wire [63:0] _8725;
    wire _8726;
    wire _8727;
    wire _8715;
    wire [63:0] _8712;
    wire [63:0] _8713;
    wire [62:0] _8714;
    wire [63:0] _8716;
    wire _8717;
    wire _8718;
    wire _8706;
    wire [63:0] _8703;
    wire [63:0] _8704;
    wire [62:0] _8705;
    wire [63:0] _8707;
    wire _8708;
    wire _8709;
    wire _8697;
    wire [63:0] _8694;
    wire [63:0] _8695;
    wire [62:0] _8696;
    wire [63:0] _8698;
    wire _8699;
    wire _8700;
    wire _8688;
    wire [63:0] _8685;
    wire [63:0] _8686;
    wire [62:0] _8687;
    wire [63:0] _8689;
    wire _8690;
    wire _8691;
    wire _8679;
    wire [63:0] _8676;
    wire [63:0] _8677;
    wire [62:0] _8678;
    wire [63:0] _8680;
    wire _8681;
    wire _8682;
    wire _8670;
    wire [63:0] _8667;
    wire [63:0] _8668;
    wire [62:0] _8669;
    wire [63:0] _8671;
    wire _8672;
    wire _8673;
    wire _8661;
    wire [63:0] _8658;
    wire [63:0] _8659;
    wire [62:0] _8660;
    wire [63:0] _8662;
    wire _8663;
    wire _8664;
    wire _8652;
    wire [63:0] _8649;
    wire [63:0] _8650;
    wire [62:0] _8651;
    wire [63:0] _8653;
    wire _8654;
    wire _8655;
    wire _8643;
    wire [63:0] _8640;
    wire [63:0] _8641;
    wire [62:0] _8642;
    wire [63:0] _8644;
    wire _8645;
    wire _8646;
    wire _8634;
    wire [63:0] _8631;
    wire [63:0] _8632;
    wire [62:0] _8633;
    wire [63:0] _8635;
    wire _8636;
    wire _8637;
    wire _8625;
    wire [63:0] _8622;
    wire [63:0] _8623;
    wire [62:0] _8624;
    wire [63:0] _8626;
    wire _8627;
    wire _8628;
    wire _8616;
    wire [63:0] _8613;
    wire [63:0] _8614;
    wire [62:0] _8615;
    wire [63:0] _8617;
    wire _8618;
    wire _8619;
    wire _8607;
    wire [63:0] _8604;
    wire [63:0] _8605;
    wire [62:0] _8606;
    wire [63:0] _8608;
    wire _8609;
    wire _8610;
    wire _8598;
    wire [63:0] _8595;
    wire [63:0] _8596;
    wire [62:0] _8597;
    wire [63:0] _8599;
    wire _8600;
    wire _8601;
    wire _8589;
    wire [63:0] _8586;
    wire [63:0] _8587;
    wire [62:0] _8588;
    wire [63:0] _8590;
    wire _8591;
    wire _8592;
    wire _8580;
    wire [63:0] _8577;
    wire [63:0] _8578;
    wire [62:0] _8579;
    wire [63:0] _8581;
    wire _8582;
    wire _8583;
    wire _8571;
    wire [63:0] _8568;
    wire [63:0] _8569;
    wire [62:0] _8570;
    wire [63:0] _8572;
    wire _8573;
    wire _8574;
    wire _8562;
    wire [63:0] _8559;
    wire [63:0] _8560;
    wire [62:0] _8561;
    wire [63:0] _8563;
    wire _8564;
    wire _8565;
    wire _8553;
    wire [63:0] _8550;
    wire [63:0] _8551;
    wire [62:0] _8552;
    wire [63:0] _8554;
    wire _8555;
    wire _8556;
    wire _8544;
    wire [63:0] _8541;
    wire [63:0] _8542;
    wire [62:0] _8543;
    wire [63:0] _8545;
    wire _8546;
    wire _8547;
    wire _8535;
    wire [63:0] _8532;
    wire [63:0] _8533;
    wire [62:0] _8534;
    wire [63:0] _8536;
    wire _8537;
    wire _8538;
    wire _8526;
    wire [63:0] _8523;
    wire [63:0] _8524;
    wire [62:0] _8525;
    wire [63:0] _8527;
    wire _8528;
    wire _8529;
    wire _8517;
    wire [63:0] _8514;
    wire [63:0] _8515;
    wire [62:0] _8516;
    wire [63:0] _8518;
    wire _8519;
    wire _8520;
    wire _8508;
    wire [63:0] _8505;
    wire [63:0] _8506;
    wire [62:0] _8507;
    wire [63:0] _8509;
    wire _8510;
    wire _8511;
    wire _8499;
    wire [63:0] _8496;
    wire [63:0] _8497;
    wire [62:0] _8498;
    wire [63:0] _8500;
    wire _8501;
    wire _8502;
    wire _8490;
    wire [63:0] _8487;
    wire [63:0] _8488;
    wire [62:0] _8489;
    wire [63:0] _8491;
    wire _8492;
    wire _8493;
    wire _8481;
    wire [63:0] _8478;
    wire [63:0] _8479;
    wire [62:0] _8480;
    wire [63:0] _8482;
    wire _8483;
    wire _8484;
    wire _8472;
    wire [63:0] _8469;
    wire [63:0] _8470;
    wire [62:0] _8471;
    wire [63:0] _8473;
    wire _8474;
    wire _8475;
    wire _8463;
    wire [63:0] _8460;
    wire [63:0] _8461;
    wire [62:0] _8462;
    wire [63:0] _8464;
    wire _8465;
    wire _8466;
    wire _8454;
    wire [63:0] _8451;
    wire [63:0] _8452;
    wire [62:0] _8453;
    wire [63:0] _8455;
    wire _8456;
    wire _8457;
    wire _8445;
    wire [63:0] _8442;
    wire [63:0] _8443;
    wire [62:0] _8444;
    wire [63:0] _8446;
    wire _8447;
    wire _8448;
    wire _8436;
    wire [63:0] _8433;
    wire [63:0] _8434;
    wire [62:0] _8435;
    wire [63:0] _8437;
    wire _8438;
    wire _8439;
    wire _8427;
    wire [63:0] _8424;
    wire [63:0] _8425;
    wire [62:0] _8426;
    wire [63:0] _8428;
    wire _8429;
    wire _8430;
    wire _8418;
    wire [63:0] _8415;
    wire [63:0] _8416;
    wire [62:0] _8417;
    wire [63:0] _8419;
    wire _8420;
    wire _8421;
    wire _8409;
    wire [63:0] _8406;
    wire [63:0] _8407;
    wire [62:0] _8408;
    wire [63:0] _8410;
    wire _8411;
    wire _8412;
    wire _8400;
    wire [63:0] _8397;
    wire [63:0] _8398;
    wire [62:0] _8399;
    wire [63:0] _8401;
    wire _8402;
    wire _8403;
    wire _8391;
    wire [63:0] _8388;
    wire [63:0] _8389;
    wire [62:0] _8390;
    wire [63:0] _8392;
    wire _8393;
    wire _8394;
    wire _8382;
    wire [63:0] _8379;
    wire [63:0] _8380;
    wire [62:0] _8381;
    wire [63:0] _8383;
    wire _8384;
    wire _8385;
    wire _8373;
    wire [63:0] _8370;
    wire [63:0] _8371;
    wire [62:0] _8372;
    wire [63:0] _8374;
    wire _8375;
    wire _8376;
    wire _8364;
    wire [63:0] _8361;
    wire [63:0] _8362;
    wire [62:0] _8363;
    wire [63:0] _8365;
    wire _8366;
    wire _8367;
    wire _8355;
    wire [63:0] _8352;
    wire [63:0] _8353;
    wire [62:0] _8354;
    wire [63:0] _8356;
    wire _8357;
    wire _8358;
    wire _8346;
    wire [63:0] _8343;
    wire [63:0] _8344;
    wire [62:0] _8345;
    wire [63:0] _8347;
    wire _8348;
    wire _8349;
    wire _8337;
    wire [63:0] _8334;
    wire [63:0] _8335;
    wire [62:0] _8336;
    wire [63:0] _8338;
    wire _8339;
    wire _8340;
    wire _8328;
    wire [63:0] _8325;
    wire [63:0] _8326;
    wire [62:0] _8327;
    wire [63:0] _8329;
    wire _8330;
    wire _8331;
    wire _8319;
    wire [63:0] _8316;
    wire [63:0] _8317;
    wire [62:0] _8318;
    wire [63:0] _8320;
    wire _8321;
    wire _8322;
    wire _8310;
    wire [63:0] _8307;
    wire [63:0] _8308;
    wire [62:0] _8309;
    wire [63:0] _8311;
    wire _8312;
    wire _8313;
    wire _8301;
    wire [63:0] _8298;
    wire [63:0] _8299;
    wire [62:0] _8300;
    wire [63:0] _8302;
    wire _8303;
    wire _8304;
    wire _8292;
    wire [63:0] _8289;
    wire [63:0] _8290;
    wire [62:0] _8291;
    wire [63:0] _8293;
    wire _8294;
    wire _8295;
    wire _8283;
    wire [63:0] _8280;
    wire [63:0] _8281;
    wire [62:0] _8282;
    wire [63:0] _8284;
    wire _8285;
    wire _8286;
    wire _8274;
    wire [63:0] _8271;
    wire [63:0] _8272;
    wire [62:0] _8273;
    wire [63:0] _8275;
    wire _8276;
    wire _8277;
    wire _8265;
    wire [63:0] _8262;
    wire [63:0] _8263;
    wire [62:0] _8264;
    wire [63:0] _8266;
    wire _8267;
    wire _8268;
    wire _8256;
    wire [63:0] _8253;
    wire [63:0] _8254;
    wire [62:0] _8255;
    wire [63:0] _8257;
    wire _8258;
    wire _8259;
    wire _8247;
    wire [63:0] _8244;
    wire [63:0] _8245;
    wire [62:0] _8246;
    wire [63:0] _8248;
    wire _8249;
    wire _8250;
    wire _8238;
    wire [63:0] _8235;
    wire [63:0] _8236;
    wire [62:0] _8237;
    wire [63:0] _8239;
    wire _8240;
    wire _8241;
    wire _8229;
    wire [63:0] _8226;
    wire [63:0] _8227;
    wire [62:0] _8228;
    wire [63:0] _8230;
    wire _8231;
    wire _8232;
    wire _8220;
    wire [63:0] _8217;
    wire [63:0] _8218;
    wire [62:0] _8219;
    wire [63:0] _8221;
    wire _8222;
    wire _8223;
    wire _8211;
    wire [63:0] _8208;
    wire [63:0] _8209;
    wire [62:0] _8210;
    wire [63:0] _8212;
    wire _8213;
    wire _8214;
    wire _8202;
    wire [63:0] _8199;
    wire [63:0] _8200;
    wire [62:0] _8201;
    wire [63:0] _8203;
    wire _8204;
    wire _8205;
    wire _8193;
    wire [63:0] _8190;
    wire [63:0] _8191;
    wire [62:0] _8192;
    wire [63:0] _8194;
    wire _8195;
    wire _8196;
    wire [63:0] _8180;
    wire [127:0] _8181;
    wire [63:0] _8182;
    wire _8183;
    wire [63:0] _8184;
    wire _8186;
    wire _8187;
    wire [63:0] _8188;
    wire [62:0] _8189;
    wire [63:0] _8197;
    wire [62:0] _8198;
    wire [63:0] _8206;
    wire [62:0] _8207;
    wire [63:0] _8215;
    wire [62:0] _8216;
    wire [63:0] _8224;
    wire [62:0] _8225;
    wire [63:0] _8233;
    wire [62:0] _8234;
    wire [63:0] _8242;
    wire [62:0] _8243;
    wire [63:0] _8251;
    wire [62:0] _8252;
    wire [63:0] _8260;
    wire [62:0] _8261;
    wire [63:0] _8269;
    wire [62:0] _8270;
    wire [63:0] _8278;
    wire [62:0] _8279;
    wire [63:0] _8287;
    wire [62:0] _8288;
    wire [63:0] _8296;
    wire [62:0] _8297;
    wire [63:0] _8305;
    wire [62:0] _8306;
    wire [63:0] _8314;
    wire [62:0] _8315;
    wire [63:0] _8323;
    wire [62:0] _8324;
    wire [63:0] _8332;
    wire [62:0] _8333;
    wire [63:0] _8341;
    wire [62:0] _8342;
    wire [63:0] _8350;
    wire [62:0] _8351;
    wire [63:0] _8359;
    wire [62:0] _8360;
    wire [63:0] _8368;
    wire [62:0] _8369;
    wire [63:0] _8377;
    wire [62:0] _8378;
    wire [63:0] _8386;
    wire [62:0] _8387;
    wire [63:0] _8395;
    wire [62:0] _8396;
    wire [63:0] _8404;
    wire [62:0] _8405;
    wire [63:0] _8413;
    wire [62:0] _8414;
    wire [63:0] _8422;
    wire [62:0] _8423;
    wire [63:0] _8431;
    wire [62:0] _8432;
    wire [63:0] _8440;
    wire [62:0] _8441;
    wire [63:0] _8449;
    wire [62:0] _8450;
    wire [63:0] _8458;
    wire [62:0] _8459;
    wire [63:0] _8467;
    wire [62:0] _8468;
    wire [63:0] _8476;
    wire [62:0] _8477;
    wire [63:0] _8485;
    wire [62:0] _8486;
    wire [63:0] _8494;
    wire [62:0] _8495;
    wire [63:0] _8503;
    wire [62:0] _8504;
    wire [63:0] _8512;
    wire [62:0] _8513;
    wire [63:0] _8521;
    wire [62:0] _8522;
    wire [63:0] _8530;
    wire [62:0] _8531;
    wire [63:0] _8539;
    wire [62:0] _8540;
    wire [63:0] _8548;
    wire [62:0] _8549;
    wire [63:0] _8557;
    wire [62:0] _8558;
    wire [63:0] _8566;
    wire [62:0] _8567;
    wire [63:0] _8575;
    wire [62:0] _8576;
    wire [63:0] _8584;
    wire [62:0] _8585;
    wire [63:0] _8593;
    wire [62:0] _8594;
    wire [63:0] _8602;
    wire [62:0] _8603;
    wire [63:0] _8611;
    wire [62:0] _8612;
    wire [63:0] _8620;
    wire [62:0] _8621;
    wire [63:0] _8629;
    wire [62:0] _8630;
    wire [63:0] _8638;
    wire [62:0] _8639;
    wire [63:0] _8647;
    wire [62:0] _8648;
    wire [63:0] _8656;
    wire [62:0] _8657;
    wire [63:0] _8665;
    wire [62:0] _8666;
    wire [63:0] _8674;
    wire [62:0] _8675;
    wire [63:0] _8683;
    wire [62:0] _8684;
    wire [63:0] _8692;
    wire [62:0] _8693;
    wire [63:0] _8701;
    wire [62:0] _8702;
    wire [63:0] _8710;
    wire [62:0] _8711;
    wire [63:0] _8719;
    wire [62:0] _8720;
    wire [63:0] _8728;
    wire [62:0] _8729;
    wire [63:0] _8737;
    wire [62:0] _8738;
    wire [63:0] _8746;
    wire [62:0] _8747;
    wire [63:0] _8755;
    wire [127:0] _8756;
    wire [63:0] _8757;
    wire _8168;
    wire [63:0] _8165;
    wire [63:0] _8166;
    wire [62:0] _8167;
    wire [63:0] _8169;
    wire _8170;
    wire _8171;
    wire _8159;
    wire [63:0] _8156;
    wire [63:0] _8157;
    wire [62:0] _8158;
    wire [63:0] _8160;
    wire _8161;
    wire _8162;
    wire _8150;
    wire [63:0] _8147;
    wire [63:0] _8148;
    wire [62:0] _8149;
    wire [63:0] _8151;
    wire _8152;
    wire _8153;
    wire _8141;
    wire [63:0] _8138;
    wire [63:0] _8139;
    wire [62:0] _8140;
    wire [63:0] _8142;
    wire _8143;
    wire _8144;
    wire _8132;
    wire [63:0] _8129;
    wire [63:0] _8130;
    wire [62:0] _8131;
    wire [63:0] _8133;
    wire _8134;
    wire _8135;
    wire _8123;
    wire [63:0] _8120;
    wire [63:0] _8121;
    wire [62:0] _8122;
    wire [63:0] _8124;
    wire _8125;
    wire _8126;
    wire _8114;
    wire [63:0] _8111;
    wire [63:0] _8112;
    wire [62:0] _8113;
    wire [63:0] _8115;
    wire _8116;
    wire _8117;
    wire _8105;
    wire [63:0] _8102;
    wire [63:0] _8103;
    wire [62:0] _8104;
    wire [63:0] _8106;
    wire _8107;
    wire _8108;
    wire _8096;
    wire [63:0] _8093;
    wire [63:0] _8094;
    wire [62:0] _8095;
    wire [63:0] _8097;
    wire _8098;
    wire _8099;
    wire _8087;
    wire [63:0] _8084;
    wire [63:0] _8085;
    wire [62:0] _8086;
    wire [63:0] _8088;
    wire _8089;
    wire _8090;
    wire _8078;
    wire [63:0] _8075;
    wire [63:0] _8076;
    wire [62:0] _8077;
    wire [63:0] _8079;
    wire _8080;
    wire _8081;
    wire _8069;
    wire [63:0] _8066;
    wire [63:0] _8067;
    wire [62:0] _8068;
    wire [63:0] _8070;
    wire _8071;
    wire _8072;
    wire _8060;
    wire [63:0] _8057;
    wire [63:0] _8058;
    wire [62:0] _8059;
    wire [63:0] _8061;
    wire _8062;
    wire _8063;
    wire _8051;
    wire [63:0] _8048;
    wire [63:0] _8049;
    wire [62:0] _8050;
    wire [63:0] _8052;
    wire _8053;
    wire _8054;
    wire _8042;
    wire [63:0] _8039;
    wire [63:0] _8040;
    wire [62:0] _8041;
    wire [63:0] _8043;
    wire _8044;
    wire _8045;
    wire _8033;
    wire [63:0] _8030;
    wire [63:0] _8031;
    wire [62:0] _8032;
    wire [63:0] _8034;
    wire _8035;
    wire _8036;
    wire _8024;
    wire [63:0] _8021;
    wire [63:0] _8022;
    wire [62:0] _8023;
    wire [63:0] _8025;
    wire _8026;
    wire _8027;
    wire _8015;
    wire [63:0] _8012;
    wire [63:0] _8013;
    wire [62:0] _8014;
    wire [63:0] _8016;
    wire _8017;
    wire _8018;
    wire _8006;
    wire [63:0] _8003;
    wire [63:0] _8004;
    wire [62:0] _8005;
    wire [63:0] _8007;
    wire _8008;
    wire _8009;
    wire _7997;
    wire [63:0] _7994;
    wire [63:0] _7995;
    wire [62:0] _7996;
    wire [63:0] _7998;
    wire _7999;
    wire _8000;
    wire _7988;
    wire [63:0] _7985;
    wire [63:0] _7986;
    wire [62:0] _7987;
    wire [63:0] _7989;
    wire _7990;
    wire _7991;
    wire _7979;
    wire [63:0] _7976;
    wire [63:0] _7977;
    wire [62:0] _7978;
    wire [63:0] _7980;
    wire _7981;
    wire _7982;
    wire _7970;
    wire [63:0] _7967;
    wire [63:0] _7968;
    wire [62:0] _7969;
    wire [63:0] _7971;
    wire _7972;
    wire _7973;
    wire _7961;
    wire [63:0] _7958;
    wire [63:0] _7959;
    wire [62:0] _7960;
    wire [63:0] _7962;
    wire _7963;
    wire _7964;
    wire _7952;
    wire [63:0] _7949;
    wire [63:0] _7950;
    wire [62:0] _7951;
    wire [63:0] _7953;
    wire _7954;
    wire _7955;
    wire _7943;
    wire [63:0] _7940;
    wire [63:0] _7941;
    wire [62:0] _7942;
    wire [63:0] _7944;
    wire _7945;
    wire _7946;
    wire _7934;
    wire [63:0] _7931;
    wire [63:0] _7932;
    wire [62:0] _7933;
    wire [63:0] _7935;
    wire _7936;
    wire _7937;
    wire _7925;
    wire [63:0] _7922;
    wire [63:0] _7923;
    wire [62:0] _7924;
    wire [63:0] _7926;
    wire _7927;
    wire _7928;
    wire _7916;
    wire [63:0] _7913;
    wire [63:0] _7914;
    wire [62:0] _7915;
    wire [63:0] _7917;
    wire _7918;
    wire _7919;
    wire _7907;
    wire [63:0] _7904;
    wire [63:0] _7905;
    wire [62:0] _7906;
    wire [63:0] _7908;
    wire _7909;
    wire _7910;
    wire _7898;
    wire [63:0] _7895;
    wire [63:0] _7896;
    wire [62:0] _7897;
    wire [63:0] _7899;
    wire _7900;
    wire _7901;
    wire _7889;
    wire [63:0] _7886;
    wire [63:0] _7887;
    wire [62:0] _7888;
    wire [63:0] _7890;
    wire _7891;
    wire _7892;
    wire _7880;
    wire [63:0] _7877;
    wire [63:0] _7878;
    wire [62:0] _7879;
    wire [63:0] _7881;
    wire _7882;
    wire _7883;
    wire _7871;
    wire [63:0] _7868;
    wire [63:0] _7869;
    wire [62:0] _7870;
    wire [63:0] _7872;
    wire _7873;
    wire _7874;
    wire _7862;
    wire [63:0] _7859;
    wire [63:0] _7860;
    wire [62:0] _7861;
    wire [63:0] _7863;
    wire _7864;
    wire _7865;
    wire _7853;
    wire [63:0] _7850;
    wire [63:0] _7851;
    wire [62:0] _7852;
    wire [63:0] _7854;
    wire _7855;
    wire _7856;
    wire _7844;
    wire [63:0] _7841;
    wire [63:0] _7842;
    wire [62:0] _7843;
    wire [63:0] _7845;
    wire _7846;
    wire _7847;
    wire _7835;
    wire [63:0] _7832;
    wire [63:0] _7833;
    wire [62:0] _7834;
    wire [63:0] _7836;
    wire _7837;
    wire _7838;
    wire _7826;
    wire [63:0] _7823;
    wire [63:0] _7824;
    wire [62:0] _7825;
    wire [63:0] _7827;
    wire _7828;
    wire _7829;
    wire _7817;
    wire [63:0] _7814;
    wire [63:0] _7815;
    wire [62:0] _7816;
    wire [63:0] _7818;
    wire _7819;
    wire _7820;
    wire _7808;
    wire [63:0] _7805;
    wire [63:0] _7806;
    wire [62:0] _7807;
    wire [63:0] _7809;
    wire _7810;
    wire _7811;
    wire _7799;
    wire [63:0] _7796;
    wire [63:0] _7797;
    wire [62:0] _7798;
    wire [63:0] _7800;
    wire _7801;
    wire _7802;
    wire _7790;
    wire [63:0] _7787;
    wire [63:0] _7788;
    wire [62:0] _7789;
    wire [63:0] _7791;
    wire _7792;
    wire _7793;
    wire _7781;
    wire [63:0] _7778;
    wire [63:0] _7779;
    wire [62:0] _7780;
    wire [63:0] _7782;
    wire _7783;
    wire _7784;
    wire _7772;
    wire [63:0] _7769;
    wire [63:0] _7770;
    wire [62:0] _7771;
    wire [63:0] _7773;
    wire _7774;
    wire _7775;
    wire _7763;
    wire [63:0] _7760;
    wire [63:0] _7761;
    wire [62:0] _7762;
    wire [63:0] _7764;
    wire _7765;
    wire _7766;
    wire _7754;
    wire [63:0] _7751;
    wire [63:0] _7752;
    wire [62:0] _7753;
    wire [63:0] _7755;
    wire _7756;
    wire _7757;
    wire _7745;
    wire [63:0] _7742;
    wire [63:0] _7743;
    wire [62:0] _7744;
    wire [63:0] _7746;
    wire _7747;
    wire _7748;
    wire _7736;
    wire [63:0] _7733;
    wire [63:0] _7734;
    wire [62:0] _7735;
    wire [63:0] _7737;
    wire _7738;
    wire _7739;
    wire _7727;
    wire [63:0] _7724;
    wire [63:0] _7725;
    wire [62:0] _7726;
    wire [63:0] _7728;
    wire _7729;
    wire _7730;
    wire _7718;
    wire [63:0] _7715;
    wire [63:0] _7716;
    wire [62:0] _7717;
    wire [63:0] _7719;
    wire _7720;
    wire _7721;
    wire _7709;
    wire [63:0] _7706;
    wire [63:0] _7707;
    wire [62:0] _7708;
    wire [63:0] _7710;
    wire _7711;
    wire _7712;
    wire _7700;
    wire [63:0] _7697;
    wire [63:0] _7698;
    wire [62:0] _7699;
    wire [63:0] _7701;
    wire _7702;
    wire _7703;
    wire _7691;
    wire [63:0] _7688;
    wire [63:0] _7689;
    wire [62:0] _7690;
    wire [63:0] _7692;
    wire _7693;
    wire _7694;
    wire _7682;
    wire [63:0] _7679;
    wire [63:0] _7680;
    wire [62:0] _7681;
    wire [63:0] _7683;
    wire _7684;
    wire _7685;
    wire _7673;
    wire [63:0] _7670;
    wire [63:0] _7671;
    wire [62:0] _7672;
    wire [63:0] _7674;
    wire _7675;
    wire _7676;
    wire _7664;
    wire [63:0] _7661;
    wire [63:0] _7662;
    wire [62:0] _7663;
    wire [63:0] _7665;
    wire _7666;
    wire _7667;
    wire _7655;
    wire [63:0] _7652;
    wire [63:0] _7653;
    wire [62:0] _7654;
    wire [63:0] _7656;
    wire _7657;
    wire _7658;
    wire _7646;
    wire [63:0] _7643;
    wire [63:0] _7644;
    wire [62:0] _7645;
    wire [63:0] _7647;
    wire _7648;
    wire _7649;
    wire _7637;
    wire [63:0] _7634;
    wire [63:0] _7635;
    wire [62:0] _7636;
    wire [63:0] _7638;
    wire _7639;
    wire _7640;
    wire _7628;
    wire [63:0] _7625;
    wire [63:0] _7626;
    wire [62:0] _7627;
    wire [63:0] _7629;
    wire _7630;
    wire _7631;
    wire _7619;
    wire [63:0] _7616;
    wire [63:0] _7617;
    wire [62:0] _7618;
    wire [63:0] _7620;
    wire _7621;
    wire _7622;
    wire _7610;
    wire [63:0] _7607;
    wire [63:0] _7608;
    wire [62:0] _7609;
    wire [63:0] _7611;
    wire _7612;
    wire _7613;
    wire [63:0] _7600;
    wire _7601;
    wire [63:0] _7602;
    wire _7603;
    wire _7604;
    wire [63:0] _7605;
    wire [62:0] _7606;
    wire [63:0] _7614;
    wire [62:0] _7615;
    wire [63:0] _7623;
    wire [62:0] _7624;
    wire [63:0] _7632;
    wire [62:0] _7633;
    wire [63:0] _7641;
    wire [62:0] _7642;
    wire [63:0] _7650;
    wire [62:0] _7651;
    wire [63:0] _7659;
    wire [62:0] _7660;
    wire [63:0] _7668;
    wire [62:0] _7669;
    wire [63:0] _7677;
    wire [62:0] _7678;
    wire [63:0] _7686;
    wire [62:0] _7687;
    wire [63:0] _7695;
    wire [62:0] _7696;
    wire [63:0] _7704;
    wire [62:0] _7705;
    wire [63:0] _7713;
    wire [62:0] _7714;
    wire [63:0] _7722;
    wire [62:0] _7723;
    wire [63:0] _7731;
    wire [62:0] _7732;
    wire [63:0] _7740;
    wire [62:0] _7741;
    wire [63:0] _7749;
    wire [62:0] _7750;
    wire [63:0] _7758;
    wire [62:0] _7759;
    wire [63:0] _7767;
    wire [62:0] _7768;
    wire [63:0] _7776;
    wire [62:0] _7777;
    wire [63:0] _7785;
    wire [62:0] _7786;
    wire [63:0] _7794;
    wire [62:0] _7795;
    wire [63:0] _7803;
    wire [62:0] _7804;
    wire [63:0] _7812;
    wire [62:0] _7813;
    wire [63:0] _7821;
    wire [62:0] _7822;
    wire [63:0] _7830;
    wire [62:0] _7831;
    wire [63:0] _7839;
    wire [62:0] _7840;
    wire [63:0] _7848;
    wire [62:0] _7849;
    wire [63:0] _7857;
    wire [62:0] _7858;
    wire [63:0] _7866;
    wire [62:0] _7867;
    wire [63:0] _7875;
    wire [62:0] _7876;
    wire [63:0] _7884;
    wire [62:0] _7885;
    wire [63:0] _7893;
    wire [62:0] _7894;
    wire [63:0] _7902;
    wire [62:0] _7903;
    wire [63:0] _7911;
    wire [62:0] _7912;
    wire [63:0] _7920;
    wire [62:0] _7921;
    wire [63:0] _7929;
    wire [62:0] _7930;
    wire [63:0] _7938;
    wire [62:0] _7939;
    wire [63:0] _7947;
    wire [62:0] _7948;
    wire [63:0] _7956;
    wire [62:0] _7957;
    wire [63:0] _7965;
    wire [62:0] _7966;
    wire [63:0] _7974;
    wire [62:0] _7975;
    wire [63:0] _7983;
    wire [62:0] _7984;
    wire [63:0] _7992;
    wire [62:0] _7993;
    wire [63:0] _8001;
    wire [62:0] _8002;
    wire [63:0] _8010;
    wire [62:0] _8011;
    wire [63:0] _8019;
    wire [62:0] _8020;
    wire [63:0] _8028;
    wire [62:0] _8029;
    wire [63:0] _8037;
    wire [62:0] _8038;
    wire [63:0] _8046;
    wire [62:0] _8047;
    wire [63:0] _8055;
    wire [62:0] _8056;
    wire [63:0] _8064;
    wire [62:0] _8065;
    wire [63:0] _8073;
    wire [62:0] _8074;
    wire [63:0] _8082;
    wire [62:0] _8083;
    wire [63:0] _8091;
    wire [62:0] _8092;
    wire [63:0] _8100;
    wire [62:0] _8101;
    wire [63:0] _8109;
    wire [62:0] _8110;
    wire [63:0] _8118;
    wire [62:0] _8119;
    wire [63:0] _8127;
    wire [62:0] _8128;
    wire [63:0] _8136;
    wire [62:0] _8137;
    wire [63:0] _8145;
    wire [62:0] _8146;
    wire [63:0] _8154;
    wire [62:0] _8155;
    wire [63:0] _8163;
    wire [62:0] _8164;
    wire [63:0] _8172;
    wire [63:0] _8174;
    wire [127:0] _8175;
    wire [63:0] _8176;
    wire [63:0] _8758;
    wire _7586;
    wire [63:0] _7583;
    wire [63:0] _7584;
    wire [62:0] _7585;
    wire [63:0] _7587;
    wire _7588;
    wire _7589;
    wire _7577;
    wire [63:0] _7574;
    wire [63:0] _7575;
    wire [62:0] _7576;
    wire [63:0] _7578;
    wire _7579;
    wire _7580;
    wire _7568;
    wire [63:0] _7565;
    wire [63:0] _7566;
    wire [62:0] _7567;
    wire [63:0] _7569;
    wire _7570;
    wire _7571;
    wire _7559;
    wire [63:0] _7556;
    wire [63:0] _7557;
    wire [62:0] _7558;
    wire [63:0] _7560;
    wire _7561;
    wire _7562;
    wire _7550;
    wire [63:0] _7547;
    wire [63:0] _7548;
    wire [62:0] _7549;
    wire [63:0] _7551;
    wire _7552;
    wire _7553;
    wire _7541;
    wire [63:0] _7538;
    wire [63:0] _7539;
    wire [62:0] _7540;
    wire [63:0] _7542;
    wire _7543;
    wire _7544;
    wire _7532;
    wire [63:0] _7529;
    wire [63:0] _7530;
    wire [62:0] _7531;
    wire [63:0] _7533;
    wire _7534;
    wire _7535;
    wire _7523;
    wire [63:0] _7520;
    wire [63:0] _7521;
    wire [62:0] _7522;
    wire [63:0] _7524;
    wire _7525;
    wire _7526;
    wire _7514;
    wire [63:0] _7511;
    wire [63:0] _7512;
    wire [62:0] _7513;
    wire [63:0] _7515;
    wire _7516;
    wire _7517;
    wire _7505;
    wire [63:0] _7502;
    wire [63:0] _7503;
    wire [62:0] _7504;
    wire [63:0] _7506;
    wire _7507;
    wire _7508;
    wire _7496;
    wire [63:0] _7493;
    wire [63:0] _7494;
    wire [62:0] _7495;
    wire [63:0] _7497;
    wire _7498;
    wire _7499;
    wire _7487;
    wire [63:0] _7484;
    wire [63:0] _7485;
    wire [62:0] _7486;
    wire [63:0] _7488;
    wire _7489;
    wire _7490;
    wire _7478;
    wire [63:0] _7475;
    wire [63:0] _7476;
    wire [62:0] _7477;
    wire [63:0] _7479;
    wire _7480;
    wire _7481;
    wire _7469;
    wire [63:0] _7466;
    wire [63:0] _7467;
    wire [62:0] _7468;
    wire [63:0] _7470;
    wire _7471;
    wire _7472;
    wire _7460;
    wire [63:0] _7457;
    wire [63:0] _7458;
    wire [62:0] _7459;
    wire [63:0] _7461;
    wire _7462;
    wire _7463;
    wire _7451;
    wire [63:0] _7448;
    wire [63:0] _7449;
    wire [62:0] _7450;
    wire [63:0] _7452;
    wire _7453;
    wire _7454;
    wire _7442;
    wire [63:0] _7439;
    wire [63:0] _7440;
    wire [62:0] _7441;
    wire [63:0] _7443;
    wire _7444;
    wire _7445;
    wire _7433;
    wire [63:0] _7430;
    wire [63:0] _7431;
    wire [62:0] _7432;
    wire [63:0] _7434;
    wire _7435;
    wire _7436;
    wire _7424;
    wire [63:0] _7421;
    wire [63:0] _7422;
    wire [62:0] _7423;
    wire [63:0] _7425;
    wire _7426;
    wire _7427;
    wire _7415;
    wire [63:0] _7412;
    wire [63:0] _7413;
    wire [62:0] _7414;
    wire [63:0] _7416;
    wire _7417;
    wire _7418;
    wire _7406;
    wire [63:0] _7403;
    wire [63:0] _7404;
    wire [62:0] _7405;
    wire [63:0] _7407;
    wire _7408;
    wire _7409;
    wire _7397;
    wire [63:0] _7394;
    wire [63:0] _7395;
    wire [62:0] _7396;
    wire [63:0] _7398;
    wire _7399;
    wire _7400;
    wire _7388;
    wire [63:0] _7385;
    wire [63:0] _7386;
    wire [62:0] _7387;
    wire [63:0] _7389;
    wire _7390;
    wire _7391;
    wire _7379;
    wire [63:0] _7376;
    wire [63:0] _7377;
    wire [62:0] _7378;
    wire [63:0] _7380;
    wire _7381;
    wire _7382;
    wire _7370;
    wire [63:0] _7367;
    wire [63:0] _7368;
    wire [62:0] _7369;
    wire [63:0] _7371;
    wire _7372;
    wire _7373;
    wire _7361;
    wire [63:0] _7358;
    wire [63:0] _7359;
    wire [62:0] _7360;
    wire [63:0] _7362;
    wire _7363;
    wire _7364;
    wire _7352;
    wire [63:0] _7349;
    wire [63:0] _7350;
    wire [62:0] _7351;
    wire [63:0] _7353;
    wire _7354;
    wire _7355;
    wire _7343;
    wire [63:0] _7340;
    wire [63:0] _7341;
    wire [62:0] _7342;
    wire [63:0] _7344;
    wire _7345;
    wire _7346;
    wire _7334;
    wire [63:0] _7331;
    wire [63:0] _7332;
    wire [62:0] _7333;
    wire [63:0] _7335;
    wire _7336;
    wire _7337;
    wire _7325;
    wire [63:0] _7322;
    wire [63:0] _7323;
    wire [62:0] _7324;
    wire [63:0] _7326;
    wire _7327;
    wire _7328;
    wire _7316;
    wire [63:0] _7313;
    wire [63:0] _7314;
    wire [62:0] _7315;
    wire [63:0] _7317;
    wire _7318;
    wire _7319;
    wire _7307;
    wire [63:0] _7304;
    wire [63:0] _7305;
    wire [62:0] _7306;
    wire [63:0] _7308;
    wire _7309;
    wire _7310;
    wire _7298;
    wire [63:0] _7295;
    wire [63:0] _7296;
    wire [62:0] _7297;
    wire [63:0] _7299;
    wire _7300;
    wire _7301;
    wire _7289;
    wire [63:0] _7286;
    wire [63:0] _7287;
    wire [62:0] _7288;
    wire [63:0] _7290;
    wire _7291;
    wire _7292;
    wire _7280;
    wire [63:0] _7277;
    wire [63:0] _7278;
    wire [62:0] _7279;
    wire [63:0] _7281;
    wire _7282;
    wire _7283;
    wire _7271;
    wire [63:0] _7268;
    wire [63:0] _7269;
    wire [62:0] _7270;
    wire [63:0] _7272;
    wire _7273;
    wire _7274;
    wire _7262;
    wire [63:0] _7259;
    wire [63:0] _7260;
    wire [62:0] _7261;
    wire [63:0] _7263;
    wire _7264;
    wire _7265;
    wire _7253;
    wire [63:0] _7250;
    wire [63:0] _7251;
    wire [62:0] _7252;
    wire [63:0] _7254;
    wire _7255;
    wire _7256;
    wire _7244;
    wire [63:0] _7241;
    wire [63:0] _7242;
    wire [62:0] _7243;
    wire [63:0] _7245;
    wire _7246;
    wire _7247;
    wire _7235;
    wire [63:0] _7232;
    wire [63:0] _7233;
    wire [62:0] _7234;
    wire [63:0] _7236;
    wire _7237;
    wire _7238;
    wire _7226;
    wire [63:0] _7223;
    wire [63:0] _7224;
    wire [62:0] _7225;
    wire [63:0] _7227;
    wire _7228;
    wire _7229;
    wire _7217;
    wire [63:0] _7214;
    wire [63:0] _7215;
    wire [62:0] _7216;
    wire [63:0] _7218;
    wire _7219;
    wire _7220;
    wire _7208;
    wire [63:0] _7205;
    wire [63:0] _7206;
    wire [62:0] _7207;
    wire [63:0] _7209;
    wire _7210;
    wire _7211;
    wire _7199;
    wire [63:0] _7196;
    wire [63:0] _7197;
    wire [62:0] _7198;
    wire [63:0] _7200;
    wire _7201;
    wire _7202;
    wire _7190;
    wire [63:0] _7187;
    wire [63:0] _7188;
    wire [62:0] _7189;
    wire [63:0] _7191;
    wire _7192;
    wire _7193;
    wire _7181;
    wire [63:0] _7178;
    wire [63:0] _7179;
    wire [62:0] _7180;
    wire [63:0] _7182;
    wire _7183;
    wire _7184;
    wire _7172;
    wire [63:0] _7169;
    wire [63:0] _7170;
    wire [62:0] _7171;
    wire [63:0] _7173;
    wire _7174;
    wire _7175;
    wire _7163;
    wire [63:0] _7160;
    wire [63:0] _7161;
    wire [62:0] _7162;
    wire [63:0] _7164;
    wire _7165;
    wire _7166;
    wire _7154;
    wire [63:0] _7151;
    wire [63:0] _7152;
    wire [62:0] _7153;
    wire [63:0] _7155;
    wire _7156;
    wire _7157;
    wire _7145;
    wire [63:0] _7142;
    wire [63:0] _7143;
    wire [62:0] _7144;
    wire [63:0] _7146;
    wire _7147;
    wire _7148;
    wire _7136;
    wire [63:0] _7133;
    wire [63:0] _7134;
    wire [62:0] _7135;
    wire [63:0] _7137;
    wire _7138;
    wire _7139;
    wire _7127;
    wire [63:0] _7124;
    wire [63:0] _7125;
    wire [62:0] _7126;
    wire [63:0] _7128;
    wire _7129;
    wire _7130;
    wire _7118;
    wire [63:0] _7115;
    wire [63:0] _7116;
    wire [62:0] _7117;
    wire [63:0] _7119;
    wire _7120;
    wire _7121;
    wire _7109;
    wire [63:0] _7106;
    wire [63:0] _7107;
    wire [62:0] _7108;
    wire [63:0] _7110;
    wire _7111;
    wire _7112;
    wire _7100;
    wire [63:0] _7097;
    wire [63:0] _7098;
    wire [62:0] _7099;
    wire [63:0] _7101;
    wire _7102;
    wire _7103;
    wire _7091;
    wire [63:0] _7088;
    wire [63:0] _7089;
    wire [62:0] _7090;
    wire [63:0] _7092;
    wire _7093;
    wire _7094;
    wire _7082;
    wire [63:0] _7079;
    wire [63:0] _7080;
    wire [62:0] _7081;
    wire [63:0] _7083;
    wire _7084;
    wire _7085;
    wire _7073;
    wire [63:0] _7070;
    wire [63:0] _7071;
    wire [62:0] _7072;
    wire [63:0] _7074;
    wire _7075;
    wire _7076;
    wire _7064;
    wire [63:0] _7061;
    wire [63:0] _7062;
    wire [62:0] _7063;
    wire [63:0] _7065;
    wire _7066;
    wire _7067;
    wire _7055;
    wire [63:0] _7052;
    wire [63:0] _7053;
    wire [62:0] _7054;
    wire [63:0] _7056;
    wire _7057;
    wire _7058;
    wire _7046;
    wire [63:0] _7043;
    wire [63:0] _7044;
    wire [62:0] _7045;
    wire [63:0] _7047;
    wire _7048;
    wire _7049;
    wire _7037;
    wire [63:0] _7034;
    wire [63:0] _7035;
    wire [62:0] _7036;
    wire [63:0] _7038;
    wire _7039;
    wire _7040;
    wire _7028;
    wire [63:0] _7025;
    wire [63:0] _7026;
    wire [62:0] _7027;
    wire [63:0] _7029;
    wire _7030;
    wire _7031;
    wire [63:0] _7020;
    wire [63:0] _7016;
    wire [63:0] _7017;
    wire _7018;
    wire [63:0] _7019;
    wire _7021;
    wire _7022;
    wire [63:0] _7023;
    wire [62:0] _7024;
    wire [63:0] _7032;
    wire [62:0] _7033;
    wire [63:0] _7041;
    wire [62:0] _7042;
    wire [63:0] _7050;
    wire [62:0] _7051;
    wire [63:0] _7059;
    wire [62:0] _7060;
    wire [63:0] _7068;
    wire [62:0] _7069;
    wire [63:0] _7077;
    wire [62:0] _7078;
    wire [63:0] _7086;
    wire [62:0] _7087;
    wire [63:0] _7095;
    wire [62:0] _7096;
    wire [63:0] _7104;
    wire [62:0] _7105;
    wire [63:0] _7113;
    wire [62:0] _7114;
    wire [63:0] _7122;
    wire [62:0] _7123;
    wire [63:0] _7131;
    wire [62:0] _7132;
    wire [63:0] _7140;
    wire [62:0] _7141;
    wire [63:0] _7149;
    wire [62:0] _7150;
    wire [63:0] _7158;
    wire [62:0] _7159;
    wire [63:0] _7167;
    wire [62:0] _7168;
    wire [63:0] _7176;
    wire [62:0] _7177;
    wire [63:0] _7185;
    wire [62:0] _7186;
    wire [63:0] _7194;
    wire [62:0] _7195;
    wire [63:0] _7203;
    wire [62:0] _7204;
    wire [63:0] _7212;
    wire [62:0] _7213;
    wire [63:0] _7221;
    wire [62:0] _7222;
    wire [63:0] _7230;
    wire [62:0] _7231;
    wire [63:0] _7239;
    wire [62:0] _7240;
    wire [63:0] _7248;
    wire [62:0] _7249;
    wire [63:0] _7257;
    wire [62:0] _7258;
    wire [63:0] _7266;
    wire [62:0] _7267;
    wire [63:0] _7275;
    wire [62:0] _7276;
    wire [63:0] _7284;
    wire [62:0] _7285;
    wire [63:0] _7293;
    wire [62:0] _7294;
    wire [63:0] _7302;
    wire [62:0] _7303;
    wire [63:0] _7311;
    wire [62:0] _7312;
    wire [63:0] _7320;
    wire [62:0] _7321;
    wire [63:0] _7329;
    wire [62:0] _7330;
    wire [63:0] _7338;
    wire [62:0] _7339;
    wire [63:0] _7347;
    wire [62:0] _7348;
    wire [63:0] _7356;
    wire [62:0] _7357;
    wire [63:0] _7365;
    wire [62:0] _7366;
    wire [63:0] _7374;
    wire [62:0] _7375;
    wire [63:0] _7383;
    wire [62:0] _7384;
    wire [63:0] _7392;
    wire [62:0] _7393;
    wire [63:0] _7401;
    wire [62:0] _7402;
    wire [63:0] _7410;
    wire [62:0] _7411;
    wire [63:0] _7419;
    wire [62:0] _7420;
    wire [63:0] _7428;
    wire [62:0] _7429;
    wire [63:0] _7437;
    wire [62:0] _7438;
    wire [63:0] _7446;
    wire [62:0] _7447;
    wire [63:0] _7455;
    wire [62:0] _7456;
    wire [63:0] _7464;
    wire [62:0] _7465;
    wire [63:0] _7473;
    wire [62:0] _7474;
    wire [63:0] _7482;
    wire [62:0] _7483;
    wire [63:0] _7491;
    wire [62:0] _7492;
    wire [63:0] _7500;
    wire [62:0] _7501;
    wire [63:0] _7509;
    wire [62:0] _7510;
    wire [63:0] _7518;
    wire [62:0] _7519;
    wire [63:0] _7527;
    wire [62:0] _7528;
    wire [63:0] _7536;
    wire [62:0] _7537;
    wire [63:0] _7545;
    wire [62:0] _7546;
    wire [63:0] _7554;
    wire [62:0] _7555;
    wire [63:0] _7563;
    wire [62:0] _7564;
    wire [63:0] _7572;
    wire [62:0] _7573;
    wire [63:0] _7581;
    wire [62:0] _7582;
    wire [63:0] _7590;
    wire [127:0] _7591;
    wire [63:0] _7592;
    wire [63:0] _7013;
    wire _7593;
    wire [63:0] _7594;
    wire _7011;
    wire [63:0] _7012;
    wire _7595;
    wire _7596;
    wire [63:0] _8759;
    wire _7000;
    wire [63:0] _6997;
    wire [63:0] _6998;
    wire [62:0] _6999;
    wire [63:0] _7001;
    wire _7002;
    wire _7003;
    wire _6991;
    wire [63:0] _6988;
    wire [63:0] _6989;
    wire [62:0] _6990;
    wire [63:0] _6992;
    wire _6993;
    wire _6994;
    wire _6982;
    wire [63:0] _6979;
    wire [63:0] _6980;
    wire [62:0] _6981;
    wire [63:0] _6983;
    wire _6984;
    wire _6985;
    wire _6973;
    wire [63:0] _6970;
    wire [63:0] _6971;
    wire [62:0] _6972;
    wire [63:0] _6974;
    wire _6975;
    wire _6976;
    wire _6964;
    wire [63:0] _6961;
    wire [63:0] _6962;
    wire [62:0] _6963;
    wire [63:0] _6965;
    wire _6966;
    wire _6967;
    wire _6955;
    wire [63:0] _6952;
    wire [63:0] _6953;
    wire [62:0] _6954;
    wire [63:0] _6956;
    wire _6957;
    wire _6958;
    wire _6946;
    wire [63:0] _6943;
    wire [63:0] _6944;
    wire [62:0] _6945;
    wire [63:0] _6947;
    wire _6948;
    wire _6949;
    wire _6937;
    wire [63:0] _6934;
    wire [63:0] _6935;
    wire [62:0] _6936;
    wire [63:0] _6938;
    wire _6939;
    wire _6940;
    wire _6928;
    wire [63:0] _6925;
    wire [63:0] _6926;
    wire [62:0] _6927;
    wire [63:0] _6929;
    wire _6930;
    wire _6931;
    wire _6919;
    wire [63:0] _6916;
    wire [63:0] _6917;
    wire [62:0] _6918;
    wire [63:0] _6920;
    wire _6921;
    wire _6922;
    wire _6910;
    wire [63:0] _6907;
    wire [63:0] _6908;
    wire [62:0] _6909;
    wire [63:0] _6911;
    wire _6912;
    wire _6913;
    wire _6901;
    wire [63:0] _6898;
    wire [63:0] _6899;
    wire [62:0] _6900;
    wire [63:0] _6902;
    wire _6903;
    wire _6904;
    wire _6892;
    wire [63:0] _6889;
    wire [63:0] _6890;
    wire [62:0] _6891;
    wire [63:0] _6893;
    wire _6894;
    wire _6895;
    wire _6883;
    wire [63:0] _6880;
    wire [63:0] _6881;
    wire [62:0] _6882;
    wire [63:0] _6884;
    wire _6885;
    wire _6886;
    wire _6874;
    wire [63:0] _6871;
    wire [63:0] _6872;
    wire [62:0] _6873;
    wire [63:0] _6875;
    wire _6876;
    wire _6877;
    wire _6865;
    wire [63:0] _6862;
    wire [63:0] _6863;
    wire [62:0] _6864;
    wire [63:0] _6866;
    wire _6867;
    wire _6868;
    wire _6856;
    wire [63:0] _6853;
    wire [63:0] _6854;
    wire [62:0] _6855;
    wire [63:0] _6857;
    wire _6858;
    wire _6859;
    wire _6847;
    wire [63:0] _6844;
    wire [63:0] _6845;
    wire [62:0] _6846;
    wire [63:0] _6848;
    wire _6849;
    wire _6850;
    wire _6838;
    wire [63:0] _6835;
    wire [63:0] _6836;
    wire [62:0] _6837;
    wire [63:0] _6839;
    wire _6840;
    wire _6841;
    wire _6829;
    wire [63:0] _6826;
    wire [63:0] _6827;
    wire [62:0] _6828;
    wire [63:0] _6830;
    wire _6831;
    wire _6832;
    wire _6820;
    wire [63:0] _6817;
    wire [63:0] _6818;
    wire [62:0] _6819;
    wire [63:0] _6821;
    wire _6822;
    wire _6823;
    wire _6811;
    wire [63:0] _6808;
    wire [63:0] _6809;
    wire [62:0] _6810;
    wire [63:0] _6812;
    wire _6813;
    wire _6814;
    wire _6802;
    wire [63:0] _6799;
    wire [63:0] _6800;
    wire [62:0] _6801;
    wire [63:0] _6803;
    wire _6804;
    wire _6805;
    wire _6793;
    wire [63:0] _6790;
    wire [63:0] _6791;
    wire [62:0] _6792;
    wire [63:0] _6794;
    wire _6795;
    wire _6796;
    wire _6784;
    wire [63:0] _6781;
    wire [63:0] _6782;
    wire [62:0] _6783;
    wire [63:0] _6785;
    wire _6786;
    wire _6787;
    wire _6775;
    wire [63:0] _6772;
    wire [63:0] _6773;
    wire [62:0] _6774;
    wire [63:0] _6776;
    wire _6777;
    wire _6778;
    wire _6766;
    wire [63:0] _6763;
    wire [63:0] _6764;
    wire [62:0] _6765;
    wire [63:0] _6767;
    wire _6768;
    wire _6769;
    wire _6757;
    wire [63:0] _6754;
    wire [63:0] _6755;
    wire [62:0] _6756;
    wire [63:0] _6758;
    wire _6759;
    wire _6760;
    wire _6748;
    wire [63:0] _6745;
    wire [63:0] _6746;
    wire [62:0] _6747;
    wire [63:0] _6749;
    wire _6750;
    wire _6751;
    wire _6739;
    wire [63:0] _6736;
    wire [63:0] _6737;
    wire [62:0] _6738;
    wire [63:0] _6740;
    wire _6741;
    wire _6742;
    wire _6730;
    wire [63:0] _6727;
    wire [63:0] _6728;
    wire [62:0] _6729;
    wire [63:0] _6731;
    wire _6732;
    wire _6733;
    wire _6721;
    wire [63:0] _6718;
    wire [63:0] _6719;
    wire [62:0] _6720;
    wire [63:0] _6722;
    wire _6723;
    wire _6724;
    wire _6712;
    wire [63:0] _6709;
    wire [63:0] _6710;
    wire [62:0] _6711;
    wire [63:0] _6713;
    wire _6714;
    wire _6715;
    wire _6703;
    wire [63:0] _6700;
    wire [63:0] _6701;
    wire [62:0] _6702;
    wire [63:0] _6704;
    wire _6705;
    wire _6706;
    wire _6694;
    wire [63:0] _6691;
    wire [63:0] _6692;
    wire [62:0] _6693;
    wire [63:0] _6695;
    wire _6696;
    wire _6697;
    wire _6685;
    wire [63:0] _6682;
    wire [63:0] _6683;
    wire [62:0] _6684;
    wire [63:0] _6686;
    wire _6687;
    wire _6688;
    wire _6676;
    wire [63:0] _6673;
    wire [63:0] _6674;
    wire [62:0] _6675;
    wire [63:0] _6677;
    wire _6678;
    wire _6679;
    wire _6667;
    wire [63:0] _6664;
    wire [63:0] _6665;
    wire [62:0] _6666;
    wire [63:0] _6668;
    wire _6669;
    wire _6670;
    wire _6658;
    wire [63:0] _6655;
    wire [63:0] _6656;
    wire [62:0] _6657;
    wire [63:0] _6659;
    wire _6660;
    wire _6661;
    wire _6649;
    wire [63:0] _6646;
    wire [63:0] _6647;
    wire [62:0] _6648;
    wire [63:0] _6650;
    wire _6651;
    wire _6652;
    wire _6640;
    wire [63:0] _6637;
    wire [63:0] _6638;
    wire [62:0] _6639;
    wire [63:0] _6641;
    wire _6642;
    wire _6643;
    wire _6631;
    wire [63:0] _6628;
    wire [63:0] _6629;
    wire [62:0] _6630;
    wire [63:0] _6632;
    wire _6633;
    wire _6634;
    wire _6622;
    wire [63:0] _6619;
    wire [63:0] _6620;
    wire [62:0] _6621;
    wire [63:0] _6623;
    wire _6624;
    wire _6625;
    wire _6613;
    wire [63:0] _6610;
    wire [63:0] _6611;
    wire [62:0] _6612;
    wire [63:0] _6614;
    wire _6615;
    wire _6616;
    wire _6604;
    wire [63:0] _6601;
    wire [63:0] _6602;
    wire [62:0] _6603;
    wire [63:0] _6605;
    wire _6606;
    wire _6607;
    wire _6595;
    wire [63:0] _6592;
    wire [63:0] _6593;
    wire [62:0] _6594;
    wire [63:0] _6596;
    wire _6597;
    wire _6598;
    wire _6586;
    wire [63:0] _6583;
    wire [63:0] _6584;
    wire [62:0] _6585;
    wire [63:0] _6587;
    wire _6588;
    wire _6589;
    wire _6577;
    wire [63:0] _6574;
    wire [63:0] _6575;
    wire [62:0] _6576;
    wire [63:0] _6578;
    wire _6579;
    wire _6580;
    wire _6568;
    wire [63:0] _6565;
    wire [63:0] _6566;
    wire [62:0] _6567;
    wire [63:0] _6569;
    wire _6570;
    wire _6571;
    wire _6559;
    wire [63:0] _6556;
    wire [63:0] _6557;
    wire [62:0] _6558;
    wire [63:0] _6560;
    wire _6561;
    wire _6562;
    wire _6550;
    wire [63:0] _6547;
    wire [63:0] _6548;
    wire [62:0] _6549;
    wire [63:0] _6551;
    wire _6552;
    wire _6553;
    wire _6541;
    wire [63:0] _6538;
    wire [63:0] _6539;
    wire [62:0] _6540;
    wire [63:0] _6542;
    wire _6543;
    wire _6544;
    wire _6532;
    wire [63:0] _6529;
    wire [63:0] _6530;
    wire [62:0] _6531;
    wire [63:0] _6533;
    wire _6534;
    wire _6535;
    wire _6523;
    wire [63:0] _6520;
    wire [63:0] _6521;
    wire [62:0] _6522;
    wire [63:0] _6524;
    wire _6525;
    wire _6526;
    wire _6514;
    wire [63:0] _6511;
    wire [63:0] _6512;
    wire [62:0] _6513;
    wire [63:0] _6515;
    wire _6516;
    wire _6517;
    wire _6505;
    wire [63:0] _6502;
    wire [63:0] _6503;
    wire [62:0] _6504;
    wire [63:0] _6506;
    wire _6507;
    wire _6508;
    wire _6496;
    wire [63:0] _6493;
    wire [63:0] _6494;
    wire [62:0] _6495;
    wire [63:0] _6497;
    wire _6498;
    wire _6499;
    wire _6487;
    wire [63:0] _6484;
    wire [63:0] _6485;
    wire [62:0] _6486;
    wire [63:0] _6488;
    wire _6489;
    wire _6490;
    wire _6478;
    wire [63:0] _6475;
    wire [63:0] _6476;
    wire [62:0] _6477;
    wire [63:0] _6479;
    wire _6480;
    wire _6481;
    wire _6469;
    wire [63:0] _6466;
    wire [63:0] _6467;
    wire [62:0] _6468;
    wire [63:0] _6470;
    wire _6471;
    wire _6472;
    wire _6460;
    wire [63:0] _6457;
    wire [63:0] _6458;
    wire [62:0] _6459;
    wire [63:0] _6461;
    wire _6462;
    wire _6463;
    wire _6451;
    wire [63:0] _6448;
    wire [63:0] _6449;
    wire [62:0] _6450;
    wire [63:0] _6452;
    wire _6453;
    wire _6454;
    wire _6442;
    wire [63:0] _6439;
    wire [63:0] _6440;
    wire [62:0] _6441;
    wire [63:0] _6443;
    wire _6444;
    wire _6445;
    wire [63:0] _6429;
    wire [127:0] _6430;
    wire [63:0] _6431;
    wire _6432;
    wire [63:0] _6433;
    wire _6435;
    wire _6436;
    wire [63:0] _6437;
    wire [62:0] _6438;
    wire [63:0] _6446;
    wire [62:0] _6447;
    wire [63:0] _6455;
    wire [62:0] _6456;
    wire [63:0] _6464;
    wire [62:0] _6465;
    wire [63:0] _6473;
    wire [62:0] _6474;
    wire [63:0] _6482;
    wire [62:0] _6483;
    wire [63:0] _6491;
    wire [62:0] _6492;
    wire [63:0] _6500;
    wire [62:0] _6501;
    wire [63:0] _6509;
    wire [62:0] _6510;
    wire [63:0] _6518;
    wire [62:0] _6519;
    wire [63:0] _6527;
    wire [62:0] _6528;
    wire [63:0] _6536;
    wire [62:0] _6537;
    wire [63:0] _6545;
    wire [62:0] _6546;
    wire [63:0] _6554;
    wire [62:0] _6555;
    wire [63:0] _6563;
    wire [62:0] _6564;
    wire [63:0] _6572;
    wire [62:0] _6573;
    wire [63:0] _6581;
    wire [62:0] _6582;
    wire [63:0] _6590;
    wire [62:0] _6591;
    wire [63:0] _6599;
    wire [62:0] _6600;
    wire [63:0] _6608;
    wire [62:0] _6609;
    wire [63:0] _6617;
    wire [62:0] _6618;
    wire [63:0] _6626;
    wire [62:0] _6627;
    wire [63:0] _6635;
    wire [62:0] _6636;
    wire [63:0] _6644;
    wire [62:0] _6645;
    wire [63:0] _6653;
    wire [62:0] _6654;
    wire [63:0] _6662;
    wire [62:0] _6663;
    wire [63:0] _6671;
    wire [62:0] _6672;
    wire [63:0] _6680;
    wire [62:0] _6681;
    wire [63:0] _6689;
    wire [62:0] _6690;
    wire [63:0] _6698;
    wire [62:0] _6699;
    wire [63:0] _6707;
    wire [62:0] _6708;
    wire [63:0] _6716;
    wire [62:0] _6717;
    wire [63:0] _6725;
    wire [62:0] _6726;
    wire [63:0] _6734;
    wire [62:0] _6735;
    wire [63:0] _6743;
    wire [62:0] _6744;
    wire [63:0] _6752;
    wire [62:0] _6753;
    wire [63:0] _6761;
    wire [62:0] _6762;
    wire [63:0] _6770;
    wire [62:0] _6771;
    wire [63:0] _6779;
    wire [62:0] _6780;
    wire [63:0] _6788;
    wire [62:0] _6789;
    wire [63:0] _6797;
    wire [62:0] _6798;
    wire [63:0] _6806;
    wire [62:0] _6807;
    wire [63:0] _6815;
    wire [62:0] _6816;
    wire [63:0] _6824;
    wire [62:0] _6825;
    wire [63:0] _6833;
    wire [62:0] _6834;
    wire [63:0] _6842;
    wire [62:0] _6843;
    wire [63:0] _6851;
    wire [62:0] _6852;
    wire [63:0] _6860;
    wire [62:0] _6861;
    wire [63:0] _6869;
    wire [62:0] _6870;
    wire [63:0] _6878;
    wire [62:0] _6879;
    wire [63:0] _6887;
    wire [62:0] _6888;
    wire [63:0] _6896;
    wire [62:0] _6897;
    wire [63:0] _6905;
    wire [62:0] _6906;
    wire [63:0] _6914;
    wire [62:0] _6915;
    wire [63:0] _6923;
    wire [62:0] _6924;
    wire [63:0] _6932;
    wire [62:0] _6933;
    wire [63:0] _6941;
    wire [62:0] _6942;
    wire [63:0] _6950;
    wire [62:0] _6951;
    wire [63:0] _6959;
    wire [62:0] _6960;
    wire [63:0] _6968;
    wire [62:0] _6969;
    wire [63:0] _6977;
    wire [62:0] _6978;
    wire [63:0] _6986;
    wire [62:0] _6987;
    wire [63:0] _6995;
    wire [62:0] _6996;
    wire [63:0] _7004;
    wire [127:0] _7005;
    wire [63:0] _7006;
    wire _6417;
    wire [63:0] _6414;
    wire [63:0] _6415;
    wire [62:0] _6416;
    wire [63:0] _6418;
    wire _6419;
    wire _6420;
    wire _6408;
    wire [63:0] _6405;
    wire [63:0] _6406;
    wire [62:0] _6407;
    wire [63:0] _6409;
    wire _6410;
    wire _6411;
    wire _6399;
    wire [63:0] _6396;
    wire [63:0] _6397;
    wire [62:0] _6398;
    wire [63:0] _6400;
    wire _6401;
    wire _6402;
    wire _6390;
    wire [63:0] _6387;
    wire [63:0] _6388;
    wire [62:0] _6389;
    wire [63:0] _6391;
    wire _6392;
    wire _6393;
    wire _6381;
    wire [63:0] _6378;
    wire [63:0] _6379;
    wire [62:0] _6380;
    wire [63:0] _6382;
    wire _6383;
    wire _6384;
    wire _6372;
    wire [63:0] _6369;
    wire [63:0] _6370;
    wire [62:0] _6371;
    wire [63:0] _6373;
    wire _6374;
    wire _6375;
    wire _6363;
    wire [63:0] _6360;
    wire [63:0] _6361;
    wire [62:0] _6362;
    wire [63:0] _6364;
    wire _6365;
    wire _6366;
    wire _6354;
    wire [63:0] _6351;
    wire [63:0] _6352;
    wire [62:0] _6353;
    wire [63:0] _6355;
    wire _6356;
    wire _6357;
    wire _6345;
    wire [63:0] _6342;
    wire [63:0] _6343;
    wire [62:0] _6344;
    wire [63:0] _6346;
    wire _6347;
    wire _6348;
    wire _6336;
    wire [63:0] _6333;
    wire [63:0] _6334;
    wire [62:0] _6335;
    wire [63:0] _6337;
    wire _6338;
    wire _6339;
    wire _6327;
    wire [63:0] _6324;
    wire [63:0] _6325;
    wire [62:0] _6326;
    wire [63:0] _6328;
    wire _6329;
    wire _6330;
    wire _6318;
    wire [63:0] _6315;
    wire [63:0] _6316;
    wire [62:0] _6317;
    wire [63:0] _6319;
    wire _6320;
    wire _6321;
    wire _6309;
    wire [63:0] _6306;
    wire [63:0] _6307;
    wire [62:0] _6308;
    wire [63:0] _6310;
    wire _6311;
    wire _6312;
    wire _6300;
    wire [63:0] _6297;
    wire [63:0] _6298;
    wire [62:0] _6299;
    wire [63:0] _6301;
    wire _6302;
    wire _6303;
    wire _6291;
    wire [63:0] _6288;
    wire [63:0] _6289;
    wire [62:0] _6290;
    wire [63:0] _6292;
    wire _6293;
    wire _6294;
    wire _6282;
    wire [63:0] _6279;
    wire [63:0] _6280;
    wire [62:0] _6281;
    wire [63:0] _6283;
    wire _6284;
    wire _6285;
    wire _6273;
    wire [63:0] _6270;
    wire [63:0] _6271;
    wire [62:0] _6272;
    wire [63:0] _6274;
    wire _6275;
    wire _6276;
    wire _6264;
    wire [63:0] _6261;
    wire [63:0] _6262;
    wire [62:0] _6263;
    wire [63:0] _6265;
    wire _6266;
    wire _6267;
    wire _6255;
    wire [63:0] _6252;
    wire [63:0] _6253;
    wire [62:0] _6254;
    wire [63:0] _6256;
    wire _6257;
    wire _6258;
    wire _6246;
    wire [63:0] _6243;
    wire [63:0] _6244;
    wire [62:0] _6245;
    wire [63:0] _6247;
    wire _6248;
    wire _6249;
    wire _6237;
    wire [63:0] _6234;
    wire [63:0] _6235;
    wire [62:0] _6236;
    wire [63:0] _6238;
    wire _6239;
    wire _6240;
    wire _6228;
    wire [63:0] _6225;
    wire [63:0] _6226;
    wire [62:0] _6227;
    wire [63:0] _6229;
    wire _6230;
    wire _6231;
    wire _6219;
    wire [63:0] _6216;
    wire [63:0] _6217;
    wire [62:0] _6218;
    wire [63:0] _6220;
    wire _6221;
    wire _6222;
    wire _6210;
    wire [63:0] _6207;
    wire [63:0] _6208;
    wire [62:0] _6209;
    wire [63:0] _6211;
    wire _6212;
    wire _6213;
    wire _6201;
    wire [63:0] _6198;
    wire [63:0] _6199;
    wire [62:0] _6200;
    wire [63:0] _6202;
    wire _6203;
    wire _6204;
    wire _6192;
    wire [63:0] _6189;
    wire [63:0] _6190;
    wire [62:0] _6191;
    wire [63:0] _6193;
    wire _6194;
    wire _6195;
    wire _6183;
    wire [63:0] _6180;
    wire [63:0] _6181;
    wire [62:0] _6182;
    wire [63:0] _6184;
    wire _6185;
    wire _6186;
    wire _6174;
    wire [63:0] _6171;
    wire [63:0] _6172;
    wire [62:0] _6173;
    wire [63:0] _6175;
    wire _6176;
    wire _6177;
    wire _6165;
    wire [63:0] _6162;
    wire [63:0] _6163;
    wire [62:0] _6164;
    wire [63:0] _6166;
    wire _6167;
    wire _6168;
    wire _6156;
    wire [63:0] _6153;
    wire [63:0] _6154;
    wire [62:0] _6155;
    wire [63:0] _6157;
    wire _6158;
    wire _6159;
    wire _6147;
    wire [63:0] _6144;
    wire [63:0] _6145;
    wire [62:0] _6146;
    wire [63:0] _6148;
    wire _6149;
    wire _6150;
    wire _6138;
    wire [63:0] _6135;
    wire [63:0] _6136;
    wire [62:0] _6137;
    wire [63:0] _6139;
    wire _6140;
    wire _6141;
    wire _6129;
    wire [63:0] _6126;
    wire [63:0] _6127;
    wire [62:0] _6128;
    wire [63:0] _6130;
    wire _6131;
    wire _6132;
    wire _6120;
    wire [63:0] _6117;
    wire [63:0] _6118;
    wire [62:0] _6119;
    wire [63:0] _6121;
    wire _6122;
    wire _6123;
    wire _6111;
    wire [63:0] _6108;
    wire [63:0] _6109;
    wire [62:0] _6110;
    wire [63:0] _6112;
    wire _6113;
    wire _6114;
    wire _6102;
    wire [63:0] _6099;
    wire [63:0] _6100;
    wire [62:0] _6101;
    wire [63:0] _6103;
    wire _6104;
    wire _6105;
    wire _6093;
    wire [63:0] _6090;
    wire [63:0] _6091;
    wire [62:0] _6092;
    wire [63:0] _6094;
    wire _6095;
    wire _6096;
    wire _6084;
    wire [63:0] _6081;
    wire [63:0] _6082;
    wire [62:0] _6083;
    wire [63:0] _6085;
    wire _6086;
    wire _6087;
    wire _6075;
    wire [63:0] _6072;
    wire [63:0] _6073;
    wire [62:0] _6074;
    wire [63:0] _6076;
    wire _6077;
    wire _6078;
    wire _6066;
    wire [63:0] _6063;
    wire [63:0] _6064;
    wire [62:0] _6065;
    wire [63:0] _6067;
    wire _6068;
    wire _6069;
    wire _6057;
    wire [63:0] _6054;
    wire [63:0] _6055;
    wire [62:0] _6056;
    wire [63:0] _6058;
    wire _6059;
    wire _6060;
    wire _6048;
    wire [63:0] _6045;
    wire [63:0] _6046;
    wire [62:0] _6047;
    wire [63:0] _6049;
    wire _6050;
    wire _6051;
    wire _6039;
    wire [63:0] _6036;
    wire [63:0] _6037;
    wire [62:0] _6038;
    wire [63:0] _6040;
    wire _6041;
    wire _6042;
    wire _6030;
    wire [63:0] _6027;
    wire [63:0] _6028;
    wire [62:0] _6029;
    wire [63:0] _6031;
    wire _6032;
    wire _6033;
    wire _6021;
    wire [63:0] _6018;
    wire [63:0] _6019;
    wire [62:0] _6020;
    wire [63:0] _6022;
    wire _6023;
    wire _6024;
    wire _6012;
    wire [63:0] _6009;
    wire [63:0] _6010;
    wire [62:0] _6011;
    wire [63:0] _6013;
    wire _6014;
    wire _6015;
    wire _6003;
    wire [63:0] _6000;
    wire [63:0] _6001;
    wire [62:0] _6002;
    wire [63:0] _6004;
    wire _6005;
    wire _6006;
    wire _5994;
    wire [63:0] _5991;
    wire [63:0] _5992;
    wire [62:0] _5993;
    wire [63:0] _5995;
    wire _5996;
    wire _5997;
    wire _5985;
    wire [63:0] _5982;
    wire [63:0] _5983;
    wire [62:0] _5984;
    wire [63:0] _5986;
    wire _5987;
    wire _5988;
    wire _5976;
    wire [63:0] _5973;
    wire [63:0] _5974;
    wire [62:0] _5975;
    wire [63:0] _5977;
    wire _5978;
    wire _5979;
    wire _5967;
    wire [63:0] _5964;
    wire [63:0] _5965;
    wire [62:0] _5966;
    wire [63:0] _5968;
    wire _5969;
    wire _5970;
    wire _5958;
    wire [63:0] _5955;
    wire [63:0] _5956;
    wire [62:0] _5957;
    wire [63:0] _5959;
    wire _5960;
    wire _5961;
    wire _5949;
    wire [63:0] _5946;
    wire [63:0] _5947;
    wire [62:0] _5948;
    wire [63:0] _5950;
    wire _5951;
    wire _5952;
    wire _5940;
    wire [63:0] _5937;
    wire [63:0] _5938;
    wire [62:0] _5939;
    wire [63:0] _5941;
    wire _5942;
    wire _5943;
    wire _5931;
    wire [63:0] _5928;
    wire [63:0] _5929;
    wire [62:0] _5930;
    wire [63:0] _5932;
    wire _5933;
    wire _5934;
    wire _5922;
    wire [63:0] _5919;
    wire [63:0] _5920;
    wire [62:0] _5921;
    wire [63:0] _5923;
    wire _5924;
    wire _5925;
    wire _5913;
    wire [63:0] _5910;
    wire [63:0] _5911;
    wire [62:0] _5912;
    wire [63:0] _5914;
    wire _5915;
    wire _5916;
    wire _5904;
    wire [63:0] _5901;
    wire [63:0] _5902;
    wire [62:0] _5903;
    wire [63:0] _5905;
    wire _5906;
    wire _5907;
    wire _5895;
    wire [63:0] _5892;
    wire [63:0] _5893;
    wire [62:0] _5894;
    wire [63:0] _5896;
    wire _5897;
    wire _5898;
    wire _5886;
    wire [63:0] _5883;
    wire [63:0] _5884;
    wire [62:0] _5885;
    wire [63:0] _5887;
    wire _5888;
    wire _5889;
    wire _5877;
    wire [63:0] _5874;
    wire [63:0] _5875;
    wire [62:0] _5876;
    wire [63:0] _5878;
    wire _5879;
    wire _5880;
    wire _5868;
    wire [63:0] _5865;
    wire [63:0] _5866;
    wire [62:0] _5867;
    wire [63:0] _5869;
    wire _5870;
    wire _5871;
    wire _5859;
    wire [63:0] _5856;
    wire [63:0] _5857;
    wire [62:0] _5858;
    wire [63:0] _5860;
    wire _5861;
    wire _5862;
    wire [63:0] _5849;
    wire _5850;
    wire [63:0] _5851;
    wire _5852;
    wire _5853;
    wire [63:0] _5854;
    wire [62:0] _5855;
    wire [63:0] _5863;
    wire [62:0] _5864;
    wire [63:0] _5872;
    wire [62:0] _5873;
    wire [63:0] _5881;
    wire [62:0] _5882;
    wire [63:0] _5890;
    wire [62:0] _5891;
    wire [63:0] _5899;
    wire [62:0] _5900;
    wire [63:0] _5908;
    wire [62:0] _5909;
    wire [63:0] _5917;
    wire [62:0] _5918;
    wire [63:0] _5926;
    wire [62:0] _5927;
    wire [63:0] _5935;
    wire [62:0] _5936;
    wire [63:0] _5944;
    wire [62:0] _5945;
    wire [63:0] _5953;
    wire [62:0] _5954;
    wire [63:0] _5962;
    wire [62:0] _5963;
    wire [63:0] _5971;
    wire [62:0] _5972;
    wire [63:0] _5980;
    wire [62:0] _5981;
    wire [63:0] _5989;
    wire [62:0] _5990;
    wire [63:0] _5998;
    wire [62:0] _5999;
    wire [63:0] _6007;
    wire [62:0] _6008;
    wire [63:0] _6016;
    wire [62:0] _6017;
    wire [63:0] _6025;
    wire [62:0] _6026;
    wire [63:0] _6034;
    wire [62:0] _6035;
    wire [63:0] _6043;
    wire [62:0] _6044;
    wire [63:0] _6052;
    wire [62:0] _6053;
    wire [63:0] _6061;
    wire [62:0] _6062;
    wire [63:0] _6070;
    wire [62:0] _6071;
    wire [63:0] _6079;
    wire [62:0] _6080;
    wire [63:0] _6088;
    wire [62:0] _6089;
    wire [63:0] _6097;
    wire [62:0] _6098;
    wire [63:0] _6106;
    wire [62:0] _6107;
    wire [63:0] _6115;
    wire [62:0] _6116;
    wire [63:0] _6124;
    wire [62:0] _6125;
    wire [63:0] _6133;
    wire [62:0] _6134;
    wire [63:0] _6142;
    wire [62:0] _6143;
    wire [63:0] _6151;
    wire [62:0] _6152;
    wire [63:0] _6160;
    wire [62:0] _6161;
    wire [63:0] _6169;
    wire [62:0] _6170;
    wire [63:0] _6178;
    wire [62:0] _6179;
    wire [63:0] _6187;
    wire [62:0] _6188;
    wire [63:0] _6196;
    wire [62:0] _6197;
    wire [63:0] _6205;
    wire [62:0] _6206;
    wire [63:0] _6214;
    wire [62:0] _6215;
    wire [63:0] _6223;
    wire [62:0] _6224;
    wire [63:0] _6232;
    wire [62:0] _6233;
    wire [63:0] _6241;
    wire [62:0] _6242;
    wire [63:0] _6250;
    wire [62:0] _6251;
    wire [63:0] _6259;
    wire [62:0] _6260;
    wire [63:0] _6268;
    wire [62:0] _6269;
    wire [63:0] _6277;
    wire [62:0] _6278;
    wire [63:0] _6286;
    wire [62:0] _6287;
    wire [63:0] _6295;
    wire [62:0] _6296;
    wire [63:0] _6304;
    wire [62:0] _6305;
    wire [63:0] _6313;
    wire [62:0] _6314;
    wire [63:0] _6322;
    wire [62:0] _6323;
    wire [63:0] _6331;
    wire [62:0] _6332;
    wire [63:0] _6340;
    wire [62:0] _6341;
    wire [63:0] _6349;
    wire [62:0] _6350;
    wire [63:0] _6358;
    wire [62:0] _6359;
    wire [63:0] _6367;
    wire [62:0] _6368;
    wire [63:0] _6376;
    wire [62:0] _6377;
    wire [63:0] _6385;
    wire [62:0] _6386;
    wire [63:0] _6394;
    wire [62:0] _6395;
    wire [63:0] _6403;
    wire [62:0] _6404;
    wire [63:0] _6412;
    wire [62:0] _6413;
    wire [63:0] _6421;
    wire [63:0] _6423;
    wire [127:0] _6424;
    wire [63:0] _6425;
    wire [63:0] _7007;
    wire _5835;
    wire [63:0] _5832;
    wire [63:0] _5833;
    wire [62:0] _5834;
    wire [63:0] _5836;
    wire _5837;
    wire _5838;
    wire _5826;
    wire [63:0] _5823;
    wire [63:0] _5824;
    wire [62:0] _5825;
    wire [63:0] _5827;
    wire _5828;
    wire _5829;
    wire _5817;
    wire [63:0] _5814;
    wire [63:0] _5815;
    wire [62:0] _5816;
    wire [63:0] _5818;
    wire _5819;
    wire _5820;
    wire _5808;
    wire [63:0] _5805;
    wire [63:0] _5806;
    wire [62:0] _5807;
    wire [63:0] _5809;
    wire _5810;
    wire _5811;
    wire _5799;
    wire [63:0] _5796;
    wire [63:0] _5797;
    wire [62:0] _5798;
    wire [63:0] _5800;
    wire _5801;
    wire _5802;
    wire _5790;
    wire [63:0] _5787;
    wire [63:0] _5788;
    wire [62:0] _5789;
    wire [63:0] _5791;
    wire _5792;
    wire _5793;
    wire _5781;
    wire [63:0] _5778;
    wire [63:0] _5779;
    wire [62:0] _5780;
    wire [63:0] _5782;
    wire _5783;
    wire _5784;
    wire _5772;
    wire [63:0] _5769;
    wire [63:0] _5770;
    wire [62:0] _5771;
    wire [63:0] _5773;
    wire _5774;
    wire _5775;
    wire _5763;
    wire [63:0] _5760;
    wire [63:0] _5761;
    wire [62:0] _5762;
    wire [63:0] _5764;
    wire _5765;
    wire _5766;
    wire _5754;
    wire [63:0] _5751;
    wire [63:0] _5752;
    wire [62:0] _5753;
    wire [63:0] _5755;
    wire _5756;
    wire _5757;
    wire _5745;
    wire [63:0] _5742;
    wire [63:0] _5743;
    wire [62:0] _5744;
    wire [63:0] _5746;
    wire _5747;
    wire _5748;
    wire _5736;
    wire [63:0] _5733;
    wire [63:0] _5734;
    wire [62:0] _5735;
    wire [63:0] _5737;
    wire _5738;
    wire _5739;
    wire _5727;
    wire [63:0] _5724;
    wire [63:0] _5725;
    wire [62:0] _5726;
    wire [63:0] _5728;
    wire _5729;
    wire _5730;
    wire _5718;
    wire [63:0] _5715;
    wire [63:0] _5716;
    wire [62:0] _5717;
    wire [63:0] _5719;
    wire _5720;
    wire _5721;
    wire _5709;
    wire [63:0] _5706;
    wire [63:0] _5707;
    wire [62:0] _5708;
    wire [63:0] _5710;
    wire _5711;
    wire _5712;
    wire _5700;
    wire [63:0] _5697;
    wire [63:0] _5698;
    wire [62:0] _5699;
    wire [63:0] _5701;
    wire _5702;
    wire _5703;
    wire _5691;
    wire [63:0] _5688;
    wire [63:0] _5689;
    wire [62:0] _5690;
    wire [63:0] _5692;
    wire _5693;
    wire _5694;
    wire _5682;
    wire [63:0] _5679;
    wire [63:0] _5680;
    wire [62:0] _5681;
    wire [63:0] _5683;
    wire _5684;
    wire _5685;
    wire _5673;
    wire [63:0] _5670;
    wire [63:0] _5671;
    wire [62:0] _5672;
    wire [63:0] _5674;
    wire _5675;
    wire _5676;
    wire _5664;
    wire [63:0] _5661;
    wire [63:0] _5662;
    wire [62:0] _5663;
    wire [63:0] _5665;
    wire _5666;
    wire _5667;
    wire _5655;
    wire [63:0] _5652;
    wire [63:0] _5653;
    wire [62:0] _5654;
    wire [63:0] _5656;
    wire _5657;
    wire _5658;
    wire _5646;
    wire [63:0] _5643;
    wire [63:0] _5644;
    wire [62:0] _5645;
    wire [63:0] _5647;
    wire _5648;
    wire _5649;
    wire _5637;
    wire [63:0] _5634;
    wire [63:0] _5635;
    wire [62:0] _5636;
    wire [63:0] _5638;
    wire _5639;
    wire _5640;
    wire _5628;
    wire [63:0] _5625;
    wire [63:0] _5626;
    wire [62:0] _5627;
    wire [63:0] _5629;
    wire _5630;
    wire _5631;
    wire _5619;
    wire [63:0] _5616;
    wire [63:0] _5617;
    wire [62:0] _5618;
    wire [63:0] _5620;
    wire _5621;
    wire _5622;
    wire _5610;
    wire [63:0] _5607;
    wire [63:0] _5608;
    wire [62:0] _5609;
    wire [63:0] _5611;
    wire _5612;
    wire _5613;
    wire _5601;
    wire [63:0] _5598;
    wire [63:0] _5599;
    wire [62:0] _5600;
    wire [63:0] _5602;
    wire _5603;
    wire _5604;
    wire _5592;
    wire [63:0] _5589;
    wire [63:0] _5590;
    wire [62:0] _5591;
    wire [63:0] _5593;
    wire _5594;
    wire _5595;
    wire _5583;
    wire [63:0] _5580;
    wire [63:0] _5581;
    wire [62:0] _5582;
    wire [63:0] _5584;
    wire _5585;
    wire _5586;
    wire _5574;
    wire [63:0] _5571;
    wire [63:0] _5572;
    wire [62:0] _5573;
    wire [63:0] _5575;
    wire _5576;
    wire _5577;
    wire _5565;
    wire [63:0] _5562;
    wire [63:0] _5563;
    wire [62:0] _5564;
    wire [63:0] _5566;
    wire _5567;
    wire _5568;
    wire _5556;
    wire [63:0] _5553;
    wire [63:0] _5554;
    wire [62:0] _5555;
    wire [63:0] _5557;
    wire _5558;
    wire _5559;
    wire _5547;
    wire [63:0] _5544;
    wire [63:0] _5545;
    wire [62:0] _5546;
    wire [63:0] _5548;
    wire _5549;
    wire _5550;
    wire _5538;
    wire [63:0] _5535;
    wire [63:0] _5536;
    wire [62:0] _5537;
    wire [63:0] _5539;
    wire _5540;
    wire _5541;
    wire _5529;
    wire [63:0] _5526;
    wire [63:0] _5527;
    wire [62:0] _5528;
    wire [63:0] _5530;
    wire _5531;
    wire _5532;
    wire _5520;
    wire [63:0] _5517;
    wire [63:0] _5518;
    wire [62:0] _5519;
    wire [63:0] _5521;
    wire _5522;
    wire _5523;
    wire _5511;
    wire [63:0] _5508;
    wire [63:0] _5509;
    wire [62:0] _5510;
    wire [63:0] _5512;
    wire _5513;
    wire _5514;
    wire _5502;
    wire [63:0] _5499;
    wire [63:0] _5500;
    wire [62:0] _5501;
    wire [63:0] _5503;
    wire _5504;
    wire _5505;
    wire _5493;
    wire [63:0] _5490;
    wire [63:0] _5491;
    wire [62:0] _5492;
    wire [63:0] _5494;
    wire _5495;
    wire _5496;
    wire _5484;
    wire [63:0] _5481;
    wire [63:0] _5482;
    wire [62:0] _5483;
    wire [63:0] _5485;
    wire _5486;
    wire _5487;
    wire _5475;
    wire [63:0] _5472;
    wire [63:0] _5473;
    wire [62:0] _5474;
    wire [63:0] _5476;
    wire _5477;
    wire _5478;
    wire _5466;
    wire [63:0] _5463;
    wire [63:0] _5464;
    wire [62:0] _5465;
    wire [63:0] _5467;
    wire _5468;
    wire _5469;
    wire _5457;
    wire [63:0] _5454;
    wire [63:0] _5455;
    wire [62:0] _5456;
    wire [63:0] _5458;
    wire _5459;
    wire _5460;
    wire _5448;
    wire [63:0] _5445;
    wire [63:0] _5446;
    wire [62:0] _5447;
    wire [63:0] _5449;
    wire _5450;
    wire _5451;
    wire _5439;
    wire [63:0] _5436;
    wire [63:0] _5437;
    wire [62:0] _5438;
    wire [63:0] _5440;
    wire _5441;
    wire _5442;
    wire _5430;
    wire [63:0] _5427;
    wire [63:0] _5428;
    wire [62:0] _5429;
    wire [63:0] _5431;
    wire _5432;
    wire _5433;
    wire _5421;
    wire [63:0] _5418;
    wire [63:0] _5419;
    wire [62:0] _5420;
    wire [63:0] _5422;
    wire _5423;
    wire _5424;
    wire _5412;
    wire [63:0] _5409;
    wire [63:0] _5410;
    wire [62:0] _5411;
    wire [63:0] _5413;
    wire _5414;
    wire _5415;
    wire _5403;
    wire [63:0] _5400;
    wire [63:0] _5401;
    wire [62:0] _5402;
    wire [63:0] _5404;
    wire _5405;
    wire _5406;
    wire _5394;
    wire [63:0] _5391;
    wire [63:0] _5392;
    wire [62:0] _5393;
    wire [63:0] _5395;
    wire _5396;
    wire _5397;
    wire _5385;
    wire [63:0] _5382;
    wire [63:0] _5383;
    wire [62:0] _5384;
    wire [63:0] _5386;
    wire _5387;
    wire _5388;
    wire _5376;
    wire [63:0] _5373;
    wire [63:0] _5374;
    wire [62:0] _5375;
    wire [63:0] _5377;
    wire _5378;
    wire _5379;
    wire _5367;
    wire [63:0] _5364;
    wire [63:0] _5365;
    wire [62:0] _5366;
    wire [63:0] _5368;
    wire _5369;
    wire _5370;
    wire _5358;
    wire [63:0] _5355;
    wire [63:0] _5356;
    wire [62:0] _5357;
    wire [63:0] _5359;
    wire _5360;
    wire _5361;
    wire _5349;
    wire [63:0] _5346;
    wire [63:0] _5347;
    wire [62:0] _5348;
    wire [63:0] _5350;
    wire _5351;
    wire _5352;
    wire _5340;
    wire [63:0] _5337;
    wire [63:0] _5338;
    wire [62:0] _5339;
    wire [63:0] _5341;
    wire _5342;
    wire _5343;
    wire _5331;
    wire [63:0] _5328;
    wire [63:0] _5329;
    wire [62:0] _5330;
    wire [63:0] _5332;
    wire _5333;
    wire _5334;
    wire _5322;
    wire [63:0] _5319;
    wire [63:0] _5320;
    wire [62:0] _5321;
    wire [63:0] _5323;
    wire _5324;
    wire _5325;
    wire _5313;
    wire [63:0] _5310;
    wire [63:0] _5311;
    wire [62:0] _5312;
    wire [63:0] _5314;
    wire _5315;
    wire _5316;
    wire _5304;
    wire [63:0] _5301;
    wire [63:0] _5302;
    wire [62:0] _5303;
    wire [63:0] _5305;
    wire _5306;
    wire _5307;
    wire _5295;
    wire [63:0] _5292;
    wire [63:0] _5293;
    wire [62:0] _5294;
    wire [63:0] _5296;
    wire _5297;
    wire _5298;
    wire _5286;
    wire [63:0] _5283;
    wire [63:0] _5284;
    wire [62:0] _5285;
    wire [63:0] _5287;
    wire _5288;
    wire _5289;
    wire _5277;
    wire [63:0] _5274;
    wire [63:0] _5275;
    wire [62:0] _5276;
    wire [63:0] _5278;
    wire _5279;
    wire _5280;
    wire [63:0] _5269;
    wire [63:0] _5265;
    wire [63:0] _5266;
    wire _5267;
    wire [63:0] _5268;
    wire _5270;
    wire _5271;
    wire [63:0] _5272;
    wire [62:0] _5273;
    wire [63:0] _5281;
    wire [62:0] _5282;
    wire [63:0] _5290;
    wire [62:0] _5291;
    wire [63:0] _5299;
    wire [62:0] _5300;
    wire [63:0] _5308;
    wire [62:0] _5309;
    wire [63:0] _5317;
    wire [62:0] _5318;
    wire [63:0] _5326;
    wire [62:0] _5327;
    wire [63:0] _5335;
    wire [62:0] _5336;
    wire [63:0] _5344;
    wire [62:0] _5345;
    wire [63:0] _5353;
    wire [62:0] _5354;
    wire [63:0] _5362;
    wire [62:0] _5363;
    wire [63:0] _5371;
    wire [62:0] _5372;
    wire [63:0] _5380;
    wire [62:0] _5381;
    wire [63:0] _5389;
    wire [62:0] _5390;
    wire [63:0] _5398;
    wire [62:0] _5399;
    wire [63:0] _5407;
    wire [62:0] _5408;
    wire [63:0] _5416;
    wire [62:0] _5417;
    wire [63:0] _5425;
    wire [62:0] _5426;
    wire [63:0] _5434;
    wire [62:0] _5435;
    wire [63:0] _5443;
    wire [62:0] _5444;
    wire [63:0] _5452;
    wire [62:0] _5453;
    wire [63:0] _5461;
    wire [62:0] _5462;
    wire [63:0] _5470;
    wire [62:0] _5471;
    wire [63:0] _5479;
    wire [62:0] _5480;
    wire [63:0] _5488;
    wire [62:0] _5489;
    wire [63:0] _5497;
    wire [62:0] _5498;
    wire [63:0] _5506;
    wire [62:0] _5507;
    wire [63:0] _5515;
    wire [62:0] _5516;
    wire [63:0] _5524;
    wire [62:0] _5525;
    wire [63:0] _5533;
    wire [62:0] _5534;
    wire [63:0] _5542;
    wire [62:0] _5543;
    wire [63:0] _5551;
    wire [62:0] _5552;
    wire [63:0] _5560;
    wire [62:0] _5561;
    wire [63:0] _5569;
    wire [62:0] _5570;
    wire [63:0] _5578;
    wire [62:0] _5579;
    wire [63:0] _5587;
    wire [62:0] _5588;
    wire [63:0] _5596;
    wire [62:0] _5597;
    wire [63:0] _5605;
    wire [62:0] _5606;
    wire [63:0] _5614;
    wire [62:0] _5615;
    wire [63:0] _5623;
    wire [62:0] _5624;
    wire [63:0] _5632;
    wire [62:0] _5633;
    wire [63:0] _5641;
    wire [62:0] _5642;
    wire [63:0] _5650;
    wire [62:0] _5651;
    wire [63:0] _5659;
    wire [62:0] _5660;
    wire [63:0] _5668;
    wire [62:0] _5669;
    wire [63:0] _5677;
    wire [62:0] _5678;
    wire [63:0] _5686;
    wire [62:0] _5687;
    wire [63:0] _5695;
    wire [62:0] _5696;
    wire [63:0] _5704;
    wire [62:0] _5705;
    wire [63:0] _5713;
    wire [62:0] _5714;
    wire [63:0] _5722;
    wire [62:0] _5723;
    wire [63:0] _5731;
    wire [62:0] _5732;
    wire [63:0] _5740;
    wire [62:0] _5741;
    wire [63:0] _5749;
    wire [62:0] _5750;
    wire [63:0] _5758;
    wire [62:0] _5759;
    wire [63:0] _5767;
    wire [62:0] _5768;
    wire [63:0] _5776;
    wire [62:0] _5777;
    wire [63:0] _5785;
    wire [62:0] _5786;
    wire [63:0] _5794;
    wire [62:0] _5795;
    wire [63:0] _5803;
    wire [62:0] _5804;
    wire [63:0] _5812;
    wire [62:0] _5813;
    wire [63:0] _5821;
    wire [62:0] _5822;
    wire [63:0] _5830;
    wire [62:0] _5831;
    wire [63:0] _5839;
    wire [127:0] _5840;
    wire [63:0] _5841;
    wire [63:0] _5262;
    wire _5842;
    wire [63:0] _5843;
    wire [63:0] _5259;
    wire _5260;
    wire [63:0] _5261;
    wire _5844;
    wire _5845;
    wire [63:0] _7008;
    wire _5249;
    wire [63:0] _5246;
    wire [63:0] _5247;
    wire [62:0] _5248;
    wire [63:0] _5250;
    wire _5251;
    wire _5252;
    wire _5240;
    wire [63:0] _5237;
    wire [63:0] _5238;
    wire [62:0] _5239;
    wire [63:0] _5241;
    wire _5242;
    wire _5243;
    wire _5231;
    wire [63:0] _5228;
    wire [63:0] _5229;
    wire [62:0] _5230;
    wire [63:0] _5232;
    wire _5233;
    wire _5234;
    wire _5222;
    wire [63:0] _5219;
    wire [63:0] _5220;
    wire [62:0] _5221;
    wire [63:0] _5223;
    wire _5224;
    wire _5225;
    wire _5213;
    wire [63:0] _5210;
    wire [63:0] _5211;
    wire [62:0] _5212;
    wire [63:0] _5214;
    wire _5215;
    wire _5216;
    wire _5204;
    wire [63:0] _5201;
    wire [63:0] _5202;
    wire [62:0] _5203;
    wire [63:0] _5205;
    wire _5206;
    wire _5207;
    wire _5195;
    wire [63:0] _5192;
    wire [63:0] _5193;
    wire [62:0] _5194;
    wire [63:0] _5196;
    wire _5197;
    wire _5198;
    wire _5186;
    wire [63:0] _5183;
    wire [63:0] _5184;
    wire [62:0] _5185;
    wire [63:0] _5187;
    wire _5188;
    wire _5189;
    wire _5177;
    wire [63:0] _5174;
    wire [63:0] _5175;
    wire [62:0] _5176;
    wire [63:0] _5178;
    wire _5179;
    wire _5180;
    wire _5168;
    wire [63:0] _5165;
    wire [63:0] _5166;
    wire [62:0] _5167;
    wire [63:0] _5169;
    wire _5170;
    wire _5171;
    wire _5159;
    wire [63:0] _5156;
    wire [63:0] _5157;
    wire [62:0] _5158;
    wire [63:0] _5160;
    wire _5161;
    wire _5162;
    wire _5150;
    wire [63:0] _5147;
    wire [63:0] _5148;
    wire [62:0] _5149;
    wire [63:0] _5151;
    wire _5152;
    wire _5153;
    wire _5141;
    wire [63:0] _5138;
    wire [63:0] _5139;
    wire [62:0] _5140;
    wire [63:0] _5142;
    wire _5143;
    wire _5144;
    wire _5132;
    wire [63:0] _5129;
    wire [63:0] _5130;
    wire [62:0] _5131;
    wire [63:0] _5133;
    wire _5134;
    wire _5135;
    wire _5123;
    wire [63:0] _5120;
    wire [63:0] _5121;
    wire [62:0] _5122;
    wire [63:0] _5124;
    wire _5125;
    wire _5126;
    wire _5114;
    wire [63:0] _5111;
    wire [63:0] _5112;
    wire [62:0] _5113;
    wire [63:0] _5115;
    wire _5116;
    wire _5117;
    wire _5105;
    wire [63:0] _5102;
    wire [63:0] _5103;
    wire [62:0] _5104;
    wire [63:0] _5106;
    wire _5107;
    wire _5108;
    wire _5096;
    wire [63:0] _5093;
    wire [63:0] _5094;
    wire [62:0] _5095;
    wire [63:0] _5097;
    wire _5098;
    wire _5099;
    wire _5087;
    wire [63:0] _5084;
    wire [63:0] _5085;
    wire [62:0] _5086;
    wire [63:0] _5088;
    wire _5089;
    wire _5090;
    wire _5078;
    wire [63:0] _5075;
    wire [63:0] _5076;
    wire [62:0] _5077;
    wire [63:0] _5079;
    wire _5080;
    wire _5081;
    wire _5069;
    wire [63:0] _5066;
    wire [63:0] _5067;
    wire [62:0] _5068;
    wire [63:0] _5070;
    wire _5071;
    wire _5072;
    wire _5060;
    wire [63:0] _5057;
    wire [63:0] _5058;
    wire [62:0] _5059;
    wire [63:0] _5061;
    wire _5062;
    wire _5063;
    wire _5051;
    wire [63:0] _5048;
    wire [63:0] _5049;
    wire [62:0] _5050;
    wire [63:0] _5052;
    wire _5053;
    wire _5054;
    wire _5042;
    wire [63:0] _5039;
    wire [63:0] _5040;
    wire [62:0] _5041;
    wire [63:0] _5043;
    wire _5044;
    wire _5045;
    wire _5033;
    wire [63:0] _5030;
    wire [63:0] _5031;
    wire [62:0] _5032;
    wire [63:0] _5034;
    wire _5035;
    wire _5036;
    wire _5024;
    wire [63:0] _5021;
    wire [63:0] _5022;
    wire [62:0] _5023;
    wire [63:0] _5025;
    wire _5026;
    wire _5027;
    wire _5015;
    wire [63:0] _5012;
    wire [63:0] _5013;
    wire [62:0] _5014;
    wire [63:0] _5016;
    wire _5017;
    wire _5018;
    wire _5006;
    wire [63:0] _5003;
    wire [63:0] _5004;
    wire [62:0] _5005;
    wire [63:0] _5007;
    wire _5008;
    wire _5009;
    wire _4997;
    wire [63:0] _4994;
    wire [63:0] _4995;
    wire [62:0] _4996;
    wire [63:0] _4998;
    wire _4999;
    wire _5000;
    wire _4988;
    wire [63:0] _4985;
    wire [63:0] _4986;
    wire [62:0] _4987;
    wire [63:0] _4989;
    wire _4990;
    wire _4991;
    wire _4979;
    wire [63:0] _4976;
    wire [63:0] _4977;
    wire [62:0] _4978;
    wire [63:0] _4980;
    wire _4981;
    wire _4982;
    wire _4970;
    wire [63:0] _4967;
    wire [63:0] _4968;
    wire [62:0] _4969;
    wire [63:0] _4971;
    wire _4972;
    wire _4973;
    wire _4961;
    wire [63:0] _4958;
    wire [63:0] _4959;
    wire [62:0] _4960;
    wire [63:0] _4962;
    wire _4963;
    wire _4964;
    wire _4952;
    wire [63:0] _4949;
    wire [63:0] _4950;
    wire [62:0] _4951;
    wire [63:0] _4953;
    wire _4954;
    wire _4955;
    wire _4943;
    wire [63:0] _4940;
    wire [63:0] _4941;
    wire [62:0] _4942;
    wire [63:0] _4944;
    wire _4945;
    wire _4946;
    wire _4934;
    wire [63:0] _4931;
    wire [63:0] _4932;
    wire [62:0] _4933;
    wire [63:0] _4935;
    wire _4936;
    wire _4937;
    wire _4925;
    wire [63:0] _4922;
    wire [63:0] _4923;
    wire [62:0] _4924;
    wire [63:0] _4926;
    wire _4927;
    wire _4928;
    wire _4916;
    wire [63:0] _4913;
    wire [63:0] _4914;
    wire [62:0] _4915;
    wire [63:0] _4917;
    wire _4918;
    wire _4919;
    wire _4907;
    wire [63:0] _4904;
    wire [63:0] _4905;
    wire [62:0] _4906;
    wire [63:0] _4908;
    wire _4909;
    wire _4910;
    wire _4898;
    wire [63:0] _4895;
    wire [63:0] _4896;
    wire [62:0] _4897;
    wire [63:0] _4899;
    wire _4900;
    wire _4901;
    wire _4889;
    wire [63:0] _4886;
    wire [63:0] _4887;
    wire [62:0] _4888;
    wire [63:0] _4890;
    wire _4891;
    wire _4892;
    wire _4880;
    wire [63:0] _4877;
    wire [63:0] _4878;
    wire [62:0] _4879;
    wire [63:0] _4881;
    wire _4882;
    wire _4883;
    wire _4871;
    wire [63:0] _4868;
    wire [63:0] _4869;
    wire [62:0] _4870;
    wire [63:0] _4872;
    wire _4873;
    wire _4874;
    wire _4862;
    wire [63:0] _4859;
    wire [63:0] _4860;
    wire [62:0] _4861;
    wire [63:0] _4863;
    wire _4864;
    wire _4865;
    wire _4853;
    wire [63:0] _4850;
    wire [63:0] _4851;
    wire [62:0] _4852;
    wire [63:0] _4854;
    wire _4855;
    wire _4856;
    wire _4844;
    wire [63:0] _4841;
    wire [63:0] _4842;
    wire [62:0] _4843;
    wire [63:0] _4845;
    wire _4846;
    wire _4847;
    wire _4835;
    wire [63:0] _4832;
    wire [63:0] _4833;
    wire [62:0] _4834;
    wire [63:0] _4836;
    wire _4837;
    wire _4838;
    wire _4826;
    wire [63:0] _4823;
    wire [63:0] _4824;
    wire [62:0] _4825;
    wire [63:0] _4827;
    wire _4828;
    wire _4829;
    wire _4817;
    wire [63:0] _4814;
    wire [63:0] _4815;
    wire [62:0] _4816;
    wire [63:0] _4818;
    wire _4819;
    wire _4820;
    wire _4808;
    wire [63:0] _4805;
    wire [63:0] _4806;
    wire [62:0] _4807;
    wire [63:0] _4809;
    wire _4810;
    wire _4811;
    wire _4799;
    wire [63:0] _4796;
    wire [63:0] _4797;
    wire [62:0] _4798;
    wire [63:0] _4800;
    wire _4801;
    wire _4802;
    wire _4790;
    wire [63:0] _4787;
    wire [63:0] _4788;
    wire [62:0] _4789;
    wire [63:0] _4791;
    wire _4792;
    wire _4793;
    wire _4781;
    wire [63:0] _4778;
    wire [63:0] _4779;
    wire [62:0] _4780;
    wire [63:0] _4782;
    wire _4783;
    wire _4784;
    wire _4772;
    wire [63:0] _4769;
    wire [63:0] _4770;
    wire [62:0] _4771;
    wire [63:0] _4773;
    wire _4774;
    wire _4775;
    wire _4763;
    wire [63:0] _4760;
    wire [63:0] _4761;
    wire [62:0] _4762;
    wire [63:0] _4764;
    wire _4765;
    wire _4766;
    wire _4754;
    wire [63:0] _4751;
    wire [63:0] _4752;
    wire [62:0] _4753;
    wire [63:0] _4755;
    wire _4756;
    wire _4757;
    wire _4745;
    wire [63:0] _4742;
    wire [63:0] _4743;
    wire [62:0] _4744;
    wire [63:0] _4746;
    wire _4747;
    wire _4748;
    wire _4736;
    wire [63:0] _4733;
    wire [63:0] _4734;
    wire [62:0] _4735;
    wire [63:0] _4737;
    wire _4738;
    wire _4739;
    wire _4727;
    wire [63:0] _4724;
    wire [63:0] _4725;
    wire [62:0] _4726;
    wire [63:0] _4728;
    wire _4729;
    wire _4730;
    wire _4718;
    wire [63:0] _4715;
    wire [63:0] _4716;
    wire [62:0] _4717;
    wire [63:0] _4719;
    wire _4720;
    wire _4721;
    wire _4709;
    wire [63:0] _4706;
    wire [63:0] _4707;
    wire [62:0] _4708;
    wire [63:0] _4710;
    wire _4711;
    wire _4712;
    wire _4700;
    wire [63:0] _4697;
    wire [63:0] _4698;
    wire [62:0] _4699;
    wire [63:0] _4701;
    wire _4702;
    wire _4703;
    wire _4691;
    wire [63:0] _4688;
    wire [63:0] _4689;
    wire [62:0] _4690;
    wire [63:0] _4692;
    wire _4693;
    wire _4694;
    wire [63:0] _4678;
    wire [127:0] _4679;
    wire [63:0] _4680;
    wire _4681;
    wire [63:0] _4682;
    wire _4684;
    wire _4685;
    wire [63:0] _4686;
    wire [62:0] _4687;
    wire [63:0] _4695;
    wire [62:0] _4696;
    wire [63:0] _4704;
    wire [62:0] _4705;
    wire [63:0] _4713;
    wire [62:0] _4714;
    wire [63:0] _4722;
    wire [62:0] _4723;
    wire [63:0] _4731;
    wire [62:0] _4732;
    wire [63:0] _4740;
    wire [62:0] _4741;
    wire [63:0] _4749;
    wire [62:0] _4750;
    wire [63:0] _4758;
    wire [62:0] _4759;
    wire [63:0] _4767;
    wire [62:0] _4768;
    wire [63:0] _4776;
    wire [62:0] _4777;
    wire [63:0] _4785;
    wire [62:0] _4786;
    wire [63:0] _4794;
    wire [62:0] _4795;
    wire [63:0] _4803;
    wire [62:0] _4804;
    wire [63:0] _4812;
    wire [62:0] _4813;
    wire [63:0] _4821;
    wire [62:0] _4822;
    wire [63:0] _4830;
    wire [62:0] _4831;
    wire [63:0] _4839;
    wire [62:0] _4840;
    wire [63:0] _4848;
    wire [62:0] _4849;
    wire [63:0] _4857;
    wire [62:0] _4858;
    wire [63:0] _4866;
    wire [62:0] _4867;
    wire [63:0] _4875;
    wire [62:0] _4876;
    wire [63:0] _4884;
    wire [62:0] _4885;
    wire [63:0] _4893;
    wire [62:0] _4894;
    wire [63:0] _4902;
    wire [62:0] _4903;
    wire [63:0] _4911;
    wire [62:0] _4912;
    wire [63:0] _4920;
    wire [62:0] _4921;
    wire [63:0] _4929;
    wire [62:0] _4930;
    wire [63:0] _4938;
    wire [62:0] _4939;
    wire [63:0] _4947;
    wire [62:0] _4948;
    wire [63:0] _4956;
    wire [62:0] _4957;
    wire [63:0] _4965;
    wire [62:0] _4966;
    wire [63:0] _4974;
    wire [62:0] _4975;
    wire [63:0] _4983;
    wire [62:0] _4984;
    wire [63:0] _4992;
    wire [62:0] _4993;
    wire [63:0] _5001;
    wire [62:0] _5002;
    wire [63:0] _5010;
    wire [62:0] _5011;
    wire [63:0] _5019;
    wire [62:0] _5020;
    wire [63:0] _5028;
    wire [62:0] _5029;
    wire [63:0] _5037;
    wire [62:0] _5038;
    wire [63:0] _5046;
    wire [62:0] _5047;
    wire [63:0] _5055;
    wire [62:0] _5056;
    wire [63:0] _5064;
    wire [62:0] _5065;
    wire [63:0] _5073;
    wire [62:0] _5074;
    wire [63:0] _5082;
    wire [62:0] _5083;
    wire [63:0] _5091;
    wire [62:0] _5092;
    wire [63:0] _5100;
    wire [62:0] _5101;
    wire [63:0] _5109;
    wire [62:0] _5110;
    wire [63:0] _5118;
    wire [62:0] _5119;
    wire [63:0] _5127;
    wire [62:0] _5128;
    wire [63:0] _5136;
    wire [62:0] _5137;
    wire [63:0] _5145;
    wire [62:0] _5146;
    wire [63:0] _5154;
    wire [62:0] _5155;
    wire [63:0] _5163;
    wire [62:0] _5164;
    wire [63:0] _5172;
    wire [62:0] _5173;
    wire [63:0] _5181;
    wire [62:0] _5182;
    wire [63:0] _5190;
    wire [62:0] _5191;
    wire [63:0] _5199;
    wire [62:0] _5200;
    wire [63:0] _5208;
    wire [62:0] _5209;
    wire [63:0] _5217;
    wire [62:0] _5218;
    wire [63:0] _5226;
    wire [62:0] _5227;
    wire [63:0] _5235;
    wire [62:0] _5236;
    wire [63:0] _5244;
    wire [62:0] _5245;
    wire [63:0] _5253;
    wire [127:0] _5254;
    wire [63:0] _5255;
    wire _4666;
    wire [63:0] _4663;
    wire [63:0] _4664;
    wire [62:0] _4665;
    wire [63:0] _4667;
    wire _4668;
    wire _4669;
    wire _4657;
    wire [63:0] _4654;
    wire [63:0] _4655;
    wire [62:0] _4656;
    wire [63:0] _4658;
    wire _4659;
    wire _4660;
    wire _4648;
    wire [63:0] _4645;
    wire [63:0] _4646;
    wire [62:0] _4647;
    wire [63:0] _4649;
    wire _4650;
    wire _4651;
    wire _4639;
    wire [63:0] _4636;
    wire [63:0] _4637;
    wire [62:0] _4638;
    wire [63:0] _4640;
    wire _4641;
    wire _4642;
    wire _4630;
    wire [63:0] _4627;
    wire [63:0] _4628;
    wire [62:0] _4629;
    wire [63:0] _4631;
    wire _4632;
    wire _4633;
    wire _4621;
    wire [63:0] _4618;
    wire [63:0] _4619;
    wire [62:0] _4620;
    wire [63:0] _4622;
    wire _4623;
    wire _4624;
    wire _4612;
    wire [63:0] _4609;
    wire [63:0] _4610;
    wire [62:0] _4611;
    wire [63:0] _4613;
    wire _4614;
    wire _4615;
    wire _4603;
    wire [63:0] _4600;
    wire [63:0] _4601;
    wire [62:0] _4602;
    wire [63:0] _4604;
    wire _4605;
    wire _4606;
    wire _4594;
    wire [63:0] _4591;
    wire [63:0] _4592;
    wire [62:0] _4593;
    wire [63:0] _4595;
    wire _4596;
    wire _4597;
    wire _4585;
    wire [63:0] _4582;
    wire [63:0] _4583;
    wire [62:0] _4584;
    wire [63:0] _4586;
    wire _4587;
    wire _4588;
    wire _4576;
    wire [63:0] _4573;
    wire [63:0] _4574;
    wire [62:0] _4575;
    wire [63:0] _4577;
    wire _4578;
    wire _4579;
    wire _4567;
    wire [63:0] _4564;
    wire [63:0] _4565;
    wire [62:0] _4566;
    wire [63:0] _4568;
    wire _4569;
    wire _4570;
    wire _4558;
    wire [63:0] _4555;
    wire [63:0] _4556;
    wire [62:0] _4557;
    wire [63:0] _4559;
    wire _4560;
    wire _4561;
    wire _4549;
    wire [63:0] _4546;
    wire [63:0] _4547;
    wire [62:0] _4548;
    wire [63:0] _4550;
    wire _4551;
    wire _4552;
    wire _4540;
    wire [63:0] _4537;
    wire [63:0] _4538;
    wire [62:0] _4539;
    wire [63:0] _4541;
    wire _4542;
    wire _4543;
    wire _4531;
    wire [63:0] _4528;
    wire [63:0] _4529;
    wire [62:0] _4530;
    wire [63:0] _4532;
    wire _4533;
    wire _4534;
    wire _4522;
    wire [63:0] _4519;
    wire [63:0] _4520;
    wire [62:0] _4521;
    wire [63:0] _4523;
    wire _4524;
    wire _4525;
    wire _4513;
    wire [63:0] _4510;
    wire [63:0] _4511;
    wire [62:0] _4512;
    wire [63:0] _4514;
    wire _4515;
    wire _4516;
    wire _4504;
    wire [63:0] _4501;
    wire [63:0] _4502;
    wire [62:0] _4503;
    wire [63:0] _4505;
    wire _4506;
    wire _4507;
    wire _4495;
    wire [63:0] _4492;
    wire [63:0] _4493;
    wire [62:0] _4494;
    wire [63:0] _4496;
    wire _4497;
    wire _4498;
    wire _4486;
    wire [63:0] _4483;
    wire [63:0] _4484;
    wire [62:0] _4485;
    wire [63:0] _4487;
    wire _4488;
    wire _4489;
    wire _4477;
    wire [63:0] _4474;
    wire [63:0] _4475;
    wire [62:0] _4476;
    wire [63:0] _4478;
    wire _4479;
    wire _4480;
    wire _4468;
    wire [63:0] _4465;
    wire [63:0] _4466;
    wire [62:0] _4467;
    wire [63:0] _4469;
    wire _4470;
    wire _4471;
    wire _4459;
    wire [63:0] _4456;
    wire [63:0] _4457;
    wire [62:0] _4458;
    wire [63:0] _4460;
    wire _4461;
    wire _4462;
    wire _4450;
    wire [63:0] _4447;
    wire [63:0] _4448;
    wire [62:0] _4449;
    wire [63:0] _4451;
    wire _4452;
    wire _4453;
    wire _4441;
    wire [63:0] _4438;
    wire [63:0] _4439;
    wire [62:0] _4440;
    wire [63:0] _4442;
    wire _4443;
    wire _4444;
    wire _4432;
    wire [63:0] _4429;
    wire [63:0] _4430;
    wire [62:0] _4431;
    wire [63:0] _4433;
    wire _4434;
    wire _4435;
    wire _4423;
    wire [63:0] _4420;
    wire [63:0] _4421;
    wire [62:0] _4422;
    wire [63:0] _4424;
    wire _4425;
    wire _4426;
    wire _4414;
    wire [63:0] _4411;
    wire [63:0] _4412;
    wire [62:0] _4413;
    wire [63:0] _4415;
    wire _4416;
    wire _4417;
    wire _4405;
    wire [63:0] _4402;
    wire [63:0] _4403;
    wire [62:0] _4404;
    wire [63:0] _4406;
    wire _4407;
    wire _4408;
    wire _4396;
    wire [63:0] _4393;
    wire [63:0] _4394;
    wire [62:0] _4395;
    wire [63:0] _4397;
    wire _4398;
    wire _4399;
    wire _4387;
    wire [63:0] _4384;
    wire [63:0] _4385;
    wire [62:0] _4386;
    wire [63:0] _4388;
    wire _4389;
    wire _4390;
    wire _4378;
    wire [63:0] _4375;
    wire [63:0] _4376;
    wire [62:0] _4377;
    wire [63:0] _4379;
    wire _4380;
    wire _4381;
    wire _4369;
    wire [63:0] _4366;
    wire [63:0] _4367;
    wire [62:0] _4368;
    wire [63:0] _4370;
    wire _4371;
    wire _4372;
    wire _4360;
    wire [63:0] _4357;
    wire [63:0] _4358;
    wire [62:0] _4359;
    wire [63:0] _4361;
    wire _4362;
    wire _4363;
    wire _4351;
    wire [63:0] _4348;
    wire [63:0] _4349;
    wire [62:0] _4350;
    wire [63:0] _4352;
    wire _4353;
    wire _4354;
    wire _4342;
    wire [63:0] _4339;
    wire [63:0] _4340;
    wire [62:0] _4341;
    wire [63:0] _4343;
    wire _4344;
    wire _4345;
    wire _4333;
    wire [63:0] _4330;
    wire [63:0] _4331;
    wire [62:0] _4332;
    wire [63:0] _4334;
    wire _4335;
    wire _4336;
    wire _4324;
    wire [63:0] _4321;
    wire [63:0] _4322;
    wire [62:0] _4323;
    wire [63:0] _4325;
    wire _4326;
    wire _4327;
    wire _4315;
    wire [63:0] _4312;
    wire [63:0] _4313;
    wire [62:0] _4314;
    wire [63:0] _4316;
    wire _4317;
    wire _4318;
    wire _4306;
    wire [63:0] _4303;
    wire [63:0] _4304;
    wire [62:0] _4305;
    wire [63:0] _4307;
    wire _4308;
    wire _4309;
    wire _4297;
    wire [63:0] _4294;
    wire [63:0] _4295;
    wire [62:0] _4296;
    wire [63:0] _4298;
    wire _4299;
    wire _4300;
    wire _4288;
    wire [63:0] _4285;
    wire [63:0] _4286;
    wire [62:0] _4287;
    wire [63:0] _4289;
    wire _4290;
    wire _4291;
    wire _4279;
    wire [63:0] _4276;
    wire [63:0] _4277;
    wire [62:0] _4278;
    wire [63:0] _4280;
    wire _4281;
    wire _4282;
    wire _4270;
    wire [63:0] _4267;
    wire [63:0] _4268;
    wire [62:0] _4269;
    wire [63:0] _4271;
    wire _4272;
    wire _4273;
    wire _4261;
    wire [63:0] _4258;
    wire [63:0] _4259;
    wire [62:0] _4260;
    wire [63:0] _4262;
    wire _4263;
    wire _4264;
    wire _4252;
    wire [63:0] _4249;
    wire [63:0] _4250;
    wire [62:0] _4251;
    wire [63:0] _4253;
    wire _4254;
    wire _4255;
    wire _4243;
    wire [63:0] _4240;
    wire [63:0] _4241;
    wire [62:0] _4242;
    wire [63:0] _4244;
    wire _4245;
    wire _4246;
    wire _4234;
    wire [63:0] _4231;
    wire [63:0] _4232;
    wire [62:0] _4233;
    wire [63:0] _4235;
    wire _4236;
    wire _4237;
    wire _4225;
    wire [63:0] _4222;
    wire [63:0] _4223;
    wire [62:0] _4224;
    wire [63:0] _4226;
    wire _4227;
    wire _4228;
    wire _4216;
    wire [63:0] _4213;
    wire [63:0] _4214;
    wire [62:0] _4215;
    wire [63:0] _4217;
    wire _4218;
    wire _4219;
    wire _4207;
    wire [63:0] _4204;
    wire [63:0] _4205;
    wire [62:0] _4206;
    wire [63:0] _4208;
    wire _4209;
    wire _4210;
    wire _4198;
    wire [63:0] _4195;
    wire [63:0] _4196;
    wire [62:0] _4197;
    wire [63:0] _4199;
    wire _4200;
    wire _4201;
    wire _4189;
    wire [63:0] _4186;
    wire [63:0] _4187;
    wire [62:0] _4188;
    wire [63:0] _4190;
    wire _4191;
    wire _4192;
    wire _4180;
    wire [63:0] _4177;
    wire [63:0] _4178;
    wire [62:0] _4179;
    wire [63:0] _4181;
    wire _4182;
    wire _4183;
    wire _4171;
    wire [63:0] _4168;
    wire [63:0] _4169;
    wire [62:0] _4170;
    wire [63:0] _4172;
    wire _4173;
    wire _4174;
    wire _4162;
    wire [63:0] _4159;
    wire [63:0] _4160;
    wire [62:0] _4161;
    wire [63:0] _4163;
    wire _4164;
    wire _4165;
    wire _4153;
    wire [63:0] _4150;
    wire [63:0] _4151;
    wire [62:0] _4152;
    wire [63:0] _4154;
    wire _4155;
    wire _4156;
    wire _4144;
    wire [63:0] _4141;
    wire [63:0] _4142;
    wire [62:0] _4143;
    wire [63:0] _4145;
    wire _4146;
    wire _4147;
    wire _4135;
    wire [63:0] _4132;
    wire [63:0] _4133;
    wire [62:0] _4134;
    wire [63:0] _4136;
    wire _4137;
    wire _4138;
    wire _4126;
    wire [63:0] _4123;
    wire [63:0] _4124;
    wire [62:0] _4125;
    wire [63:0] _4127;
    wire _4128;
    wire _4129;
    wire _4117;
    wire [63:0] _4114;
    wire [63:0] _4115;
    wire [62:0] _4116;
    wire [63:0] _4118;
    wire _4119;
    wire _4120;
    wire _4108;
    wire [63:0] _4105;
    wire [63:0] _4106;
    wire [62:0] _4107;
    wire [63:0] _4109;
    wire _4110;
    wire _4111;
    wire [63:0] _4098;
    wire _4099;
    wire [63:0] _4100;
    wire _4101;
    wire _4102;
    wire [63:0] _4103;
    wire [62:0] _4104;
    wire [63:0] _4112;
    wire [62:0] _4113;
    wire [63:0] _4121;
    wire [62:0] _4122;
    wire [63:0] _4130;
    wire [62:0] _4131;
    wire [63:0] _4139;
    wire [62:0] _4140;
    wire [63:0] _4148;
    wire [62:0] _4149;
    wire [63:0] _4157;
    wire [62:0] _4158;
    wire [63:0] _4166;
    wire [62:0] _4167;
    wire [63:0] _4175;
    wire [62:0] _4176;
    wire [63:0] _4184;
    wire [62:0] _4185;
    wire [63:0] _4193;
    wire [62:0] _4194;
    wire [63:0] _4202;
    wire [62:0] _4203;
    wire [63:0] _4211;
    wire [62:0] _4212;
    wire [63:0] _4220;
    wire [62:0] _4221;
    wire [63:0] _4229;
    wire [62:0] _4230;
    wire [63:0] _4238;
    wire [62:0] _4239;
    wire [63:0] _4247;
    wire [62:0] _4248;
    wire [63:0] _4256;
    wire [62:0] _4257;
    wire [63:0] _4265;
    wire [62:0] _4266;
    wire [63:0] _4274;
    wire [62:0] _4275;
    wire [63:0] _4283;
    wire [62:0] _4284;
    wire [63:0] _4292;
    wire [62:0] _4293;
    wire [63:0] _4301;
    wire [62:0] _4302;
    wire [63:0] _4310;
    wire [62:0] _4311;
    wire [63:0] _4319;
    wire [62:0] _4320;
    wire [63:0] _4328;
    wire [62:0] _4329;
    wire [63:0] _4337;
    wire [62:0] _4338;
    wire [63:0] _4346;
    wire [62:0] _4347;
    wire [63:0] _4355;
    wire [62:0] _4356;
    wire [63:0] _4364;
    wire [62:0] _4365;
    wire [63:0] _4373;
    wire [62:0] _4374;
    wire [63:0] _4382;
    wire [62:0] _4383;
    wire [63:0] _4391;
    wire [62:0] _4392;
    wire [63:0] _4400;
    wire [62:0] _4401;
    wire [63:0] _4409;
    wire [62:0] _4410;
    wire [63:0] _4418;
    wire [62:0] _4419;
    wire [63:0] _4427;
    wire [62:0] _4428;
    wire [63:0] _4436;
    wire [62:0] _4437;
    wire [63:0] _4445;
    wire [62:0] _4446;
    wire [63:0] _4454;
    wire [62:0] _4455;
    wire [63:0] _4463;
    wire [62:0] _4464;
    wire [63:0] _4472;
    wire [62:0] _4473;
    wire [63:0] _4481;
    wire [62:0] _4482;
    wire [63:0] _4490;
    wire [62:0] _4491;
    wire [63:0] _4499;
    wire [62:0] _4500;
    wire [63:0] _4508;
    wire [62:0] _4509;
    wire [63:0] _4517;
    wire [62:0] _4518;
    wire [63:0] _4526;
    wire [62:0] _4527;
    wire [63:0] _4535;
    wire [62:0] _4536;
    wire [63:0] _4544;
    wire [62:0] _4545;
    wire [63:0] _4553;
    wire [62:0] _4554;
    wire [63:0] _4562;
    wire [62:0] _4563;
    wire [63:0] _4571;
    wire [62:0] _4572;
    wire [63:0] _4580;
    wire [62:0] _4581;
    wire [63:0] _4589;
    wire [62:0] _4590;
    wire [63:0] _4598;
    wire [62:0] _4599;
    wire [63:0] _4607;
    wire [62:0] _4608;
    wire [63:0] _4616;
    wire [62:0] _4617;
    wire [63:0] _4625;
    wire [62:0] _4626;
    wire [63:0] _4634;
    wire [62:0] _4635;
    wire [63:0] _4643;
    wire [62:0] _4644;
    wire [63:0] _4652;
    wire [62:0] _4653;
    wire [63:0] _4661;
    wire [62:0] _4662;
    wire [63:0] _4670;
    wire [63:0] _4672;
    wire [127:0] _4673;
    wire [63:0] _4674;
    wire [63:0] _5256;
    wire _4084;
    wire [63:0] _4081;
    wire [63:0] _4082;
    wire [62:0] _4083;
    wire [63:0] _4085;
    wire _4086;
    wire _4087;
    wire _4075;
    wire [63:0] _4072;
    wire [63:0] _4073;
    wire [62:0] _4074;
    wire [63:0] _4076;
    wire _4077;
    wire _4078;
    wire _4066;
    wire [63:0] _4063;
    wire [63:0] _4064;
    wire [62:0] _4065;
    wire [63:0] _4067;
    wire _4068;
    wire _4069;
    wire _4057;
    wire [63:0] _4054;
    wire [63:0] _4055;
    wire [62:0] _4056;
    wire [63:0] _4058;
    wire _4059;
    wire _4060;
    wire _4048;
    wire [63:0] _4045;
    wire [63:0] _4046;
    wire [62:0] _4047;
    wire [63:0] _4049;
    wire _4050;
    wire _4051;
    wire _4039;
    wire [63:0] _4036;
    wire [63:0] _4037;
    wire [62:0] _4038;
    wire [63:0] _4040;
    wire _4041;
    wire _4042;
    wire _4030;
    wire [63:0] _4027;
    wire [63:0] _4028;
    wire [62:0] _4029;
    wire [63:0] _4031;
    wire _4032;
    wire _4033;
    wire _4021;
    wire [63:0] _4018;
    wire [63:0] _4019;
    wire [62:0] _4020;
    wire [63:0] _4022;
    wire _4023;
    wire _4024;
    wire _4012;
    wire [63:0] _4009;
    wire [63:0] _4010;
    wire [62:0] _4011;
    wire [63:0] _4013;
    wire _4014;
    wire _4015;
    wire _4003;
    wire [63:0] _4000;
    wire [63:0] _4001;
    wire [62:0] _4002;
    wire [63:0] _4004;
    wire _4005;
    wire _4006;
    wire _3994;
    wire [63:0] _3991;
    wire [63:0] _3992;
    wire [62:0] _3993;
    wire [63:0] _3995;
    wire _3996;
    wire _3997;
    wire _3985;
    wire [63:0] _3982;
    wire [63:0] _3983;
    wire [62:0] _3984;
    wire [63:0] _3986;
    wire _3987;
    wire _3988;
    wire _3976;
    wire [63:0] _3973;
    wire [63:0] _3974;
    wire [62:0] _3975;
    wire [63:0] _3977;
    wire _3978;
    wire _3979;
    wire _3967;
    wire [63:0] _3964;
    wire [63:0] _3965;
    wire [62:0] _3966;
    wire [63:0] _3968;
    wire _3969;
    wire _3970;
    wire _3958;
    wire [63:0] _3955;
    wire [63:0] _3956;
    wire [62:0] _3957;
    wire [63:0] _3959;
    wire _3960;
    wire _3961;
    wire _3949;
    wire [63:0] _3946;
    wire [63:0] _3947;
    wire [62:0] _3948;
    wire [63:0] _3950;
    wire _3951;
    wire _3952;
    wire _3940;
    wire [63:0] _3937;
    wire [63:0] _3938;
    wire [62:0] _3939;
    wire [63:0] _3941;
    wire _3942;
    wire _3943;
    wire _3931;
    wire [63:0] _3928;
    wire [63:0] _3929;
    wire [62:0] _3930;
    wire [63:0] _3932;
    wire _3933;
    wire _3934;
    wire _3922;
    wire [63:0] _3919;
    wire [63:0] _3920;
    wire [62:0] _3921;
    wire [63:0] _3923;
    wire _3924;
    wire _3925;
    wire _3913;
    wire [63:0] _3910;
    wire [63:0] _3911;
    wire [62:0] _3912;
    wire [63:0] _3914;
    wire _3915;
    wire _3916;
    wire _3904;
    wire [63:0] _3901;
    wire [63:0] _3902;
    wire [62:0] _3903;
    wire [63:0] _3905;
    wire _3906;
    wire _3907;
    wire _3895;
    wire [63:0] _3892;
    wire [63:0] _3893;
    wire [62:0] _3894;
    wire [63:0] _3896;
    wire _3897;
    wire _3898;
    wire _3886;
    wire [63:0] _3883;
    wire [63:0] _3884;
    wire [62:0] _3885;
    wire [63:0] _3887;
    wire _3888;
    wire _3889;
    wire _3877;
    wire [63:0] _3874;
    wire [63:0] _3875;
    wire [62:0] _3876;
    wire [63:0] _3878;
    wire _3879;
    wire _3880;
    wire _3868;
    wire [63:0] _3865;
    wire [63:0] _3866;
    wire [62:0] _3867;
    wire [63:0] _3869;
    wire _3870;
    wire _3871;
    wire _3859;
    wire [63:0] _3856;
    wire [63:0] _3857;
    wire [62:0] _3858;
    wire [63:0] _3860;
    wire _3861;
    wire _3862;
    wire _3850;
    wire [63:0] _3847;
    wire [63:0] _3848;
    wire [62:0] _3849;
    wire [63:0] _3851;
    wire _3852;
    wire _3853;
    wire _3841;
    wire [63:0] _3838;
    wire [63:0] _3839;
    wire [62:0] _3840;
    wire [63:0] _3842;
    wire _3843;
    wire _3844;
    wire _3832;
    wire [63:0] _3829;
    wire [63:0] _3830;
    wire [62:0] _3831;
    wire [63:0] _3833;
    wire _3834;
    wire _3835;
    wire _3823;
    wire [63:0] _3820;
    wire [63:0] _3821;
    wire [62:0] _3822;
    wire [63:0] _3824;
    wire _3825;
    wire _3826;
    wire _3814;
    wire [63:0] _3811;
    wire [63:0] _3812;
    wire [62:0] _3813;
    wire [63:0] _3815;
    wire _3816;
    wire _3817;
    wire _3805;
    wire [63:0] _3802;
    wire [63:0] _3803;
    wire [62:0] _3804;
    wire [63:0] _3806;
    wire _3807;
    wire _3808;
    wire _3796;
    wire [63:0] _3793;
    wire [63:0] _3794;
    wire [62:0] _3795;
    wire [63:0] _3797;
    wire _3798;
    wire _3799;
    wire _3787;
    wire [63:0] _3784;
    wire [63:0] _3785;
    wire [62:0] _3786;
    wire [63:0] _3788;
    wire _3789;
    wire _3790;
    wire _3778;
    wire [63:0] _3775;
    wire [63:0] _3776;
    wire [62:0] _3777;
    wire [63:0] _3779;
    wire _3780;
    wire _3781;
    wire _3769;
    wire [63:0] _3766;
    wire [63:0] _3767;
    wire [62:0] _3768;
    wire [63:0] _3770;
    wire _3771;
    wire _3772;
    wire _3760;
    wire [63:0] _3757;
    wire [63:0] _3758;
    wire [62:0] _3759;
    wire [63:0] _3761;
    wire _3762;
    wire _3763;
    wire _3751;
    wire [63:0] _3748;
    wire [63:0] _3749;
    wire [62:0] _3750;
    wire [63:0] _3752;
    wire _3753;
    wire _3754;
    wire _3742;
    wire [63:0] _3739;
    wire [63:0] _3740;
    wire [62:0] _3741;
    wire [63:0] _3743;
    wire _3744;
    wire _3745;
    wire _3733;
    wire [63:0] _3730;
    wire [63:0] _3731;
    wire [62:0] _3732;
    wire [63:0] _3734;
    wire _3735;
    wire _3736;
    wire _3724;
    wire [63:0] _3721;
    wire [63:0] _3722;
    wire [62:0] _3723;
    wire [63:0] _3725;
    wire _3726;
    wire _3727;
    wire _3715;
    wire [63:0] _3712;
    wire [63:0] _3713;
    wire [62:0] _3714;
    wire [63:0] _3716;
    wire _3717;
    wire _3718;
    wire _3706;
    wire [63:0] _3703;
    wire [63:0] _3704;
    wire [62:0] _3705;
    wire [63:0] _3707;
    wire _3708;
    wire _3709;
    wire _3697;
    wire [63:0] _3694;
    wire [63:0] _3695;
    wire [62:0] _3696;
    wire [63:0] _3698;
    wire _3699;
    wire _3700;
    wire _3688;
    wire [63:0] _3685;
    wire [63:0] _3686;
    wire [62:0] _3687;
    wire [63:0] _3689;
    wire _3690;
    wire _3691;
    wire _3679;
    wire [63:0] _3676;
    wire [63:0] _3677;
    wire [62:0] _3678;
    wire [63:0] _3680;
    wire _3681;
    wire _3682;
    wire _3670;
    wire [63:0] _3667;
    wire [63:0] _3668;
    wire [62:0] _3669;
    wire [63:0] _3671;
    wire _3672;
    wire _3673;
    wire _3661;
    wire [63:0] _3658;
    wire [63:0] _3659;
    wire [62:0] _3660;
    wire [63:0] _3662;
    wire _3663;
    wire _3664;
    wire _3652;
    wire [63:0] _3649;
    wire [63:0] _3650;
    wire [62:0] _3651;
    wire [63:0] _3653;
    wire _3654;
    wire _3655;
    wire _3643;
    wire [63:0] _3640;
    wire [63:0] _3641;
    wire [62:0] _3642;
    wire [63:0] _3644;
    wire _3645;
    wire _3646;
    wire _3634;
    wire [63:0] _3631;
    wire [63:0] _3632;
    wire [62:0] _3633;
    wire [63:0] _3635;
    wire _3636;
    wire _3637;
    wire _3625;
    wire [63:0] _3622;
    wire [63:0] _3623;
    wire [62:0] _3624;
    wire [63:0] _3626;
    wire _3627;
    wire _3628;
    wire _3616;
    wire [63:0] _3613;
    wire [63:0] _3614;
    wire [62:0] _3615;
    wire [63:0] _3617;
    wire _3618;
    wire _3619;
    wire _3607;
    wire [63:0] _3604;
    wire [63:0] _3605;
    wire [62:0] _3606;
    wire [63:0] _3608;
    wire _3609;
    wire _3610;
    wire _3598;
    wire [63:0] _3595;
    wire [63:0] _3596;
    wire [62:0] _3597;
    wire [63:0] _3599;
    wire _3600;
    wire _3601;
    wire _3589;
    wire [63:0] _3586;
    wire [63:0] _3587;
    wire [62:0] _3588;
    wire [63:0] _3590;
    wire _3591;
    wire _3592;
    wire _3580;
    wire [63:0] _3577;
    wire [63:0] _3578;
    wire [62:0] _3579;
    wire [63:0] _3581;
    wire _3582;
    wire _3583;
    wire _3571;
    wire [63:0] _3568;
    wire [63:0] _3569;
    wire [62:0] _3570;
    wire [63:0] _3572;
    wire _3573;
    wire _3574;
    wire _3562;
    wire [63:0] _3559;
    wire [63:0] _3560;
    wire [62:0] _3561;
    wire [63:0] _3563;
    wire _3564;
    wire _3565;
    wire _3553;
    wire [63:0] _3550;
    wire [63:0] _3551;
    wire [62:0] _3552;
    wire [63:0] _3554;
    wire _3555;
    wire _3556;
    wire _3544;
    wire [63:0] _3541;
    wire [63:0] _3542;
    wire [62:0] _3543;
    wire [63:0] _3545;
    wire _3546;
    wire _3547;
    wire _3535;
    wire [63:0] _3532;
    wire [63:0] _3533;
    wire [62:0] _3534;
    wire [63:0] _3536;
    wire _3537;
    wire _3538;
    wire _3526;
    wire [63:0] _3523;
    wire [63:0] _3524;
    wire [62:0] _3525;
    wire [63:0] _3527;
    wire _3528;
    wire _3529;
    wire [63:0] _3518;
    wire [63:0] _3514;
    wire [63:0] _3515;
    wire _3516;
    wire [63:0] _3517;
    wire _3519;
    wire _3520;
    wire [63:0] _3521;
    wire [62:0] _3522;
    wire [63:0] _3530;
    wire [62:0] _3531;
    wire [63:0] _3539;
    wire [62:0] _3540;
    wire [63:0] _3548;
    wire [62:0] _3549;
    wire [63:0] _3557;
    wire [62:0] _3558;
    wire [63:0] _3566;
    wire [62:0] _3567;
    wire [63:0] _3575;
    wire [62:0] _3576;
    wire [63:0] _3584;
    wire [62:0] _3585;
    wire [63:0] _3593;
    wire [62:0] _3594;
    wire [63:0] _3602;
    wire [62:0] _3603;
    wire [63:0] _3611;
    wire [62:0] _3612;
    wire [63:0] _3620;
    wire [62:0] _3621;
    wire [63:0] _3629;
    wire [62:0] _3630;
    wire [63:0] _3638;
    wire [62:0] _3639;
    wire [63:0] _3647;
    wire [62:0] _3648;
    wire [63:0] _3656;
    wire [62:0] _3657;
    wire [63:0] _3665;
    wire [62:0] _3666;
    wire [63:0] _3674;
    wire [62:0] _3675;
    wire [63:0] _3683;
    wire [62:0] _3684;
    wire [63:0] _3692;
    wire [62:0] _3693;
    wire [63:0] _3701;
    wire [62:0] _3702;
    wire [63:0] _3710;
    wire [62:0] _3711;
    wire [63:0] _3719;
    wire [62:0] _3720;
    wire [63:0] _3728;
    wire [62:0] _3729;
    wire [63:0] _3737;
    wire [62:0] _3738;
    wire [63:0] _3746;
    wire [62:0] _3747;
    wire [63:0] _3755;
    wire [62:0] _3756;
    wire [63:0] _3764;
    wire [62:0] _3765;
    wire [63:0] _3773;
    wire [62:0] _3774;
    wire [63:0] _3782;
    wire [62:0] _3783;
    wire [63:0] _3791;
    wire [62:0] _3792;
    wire [63:0] _3800;
    wire [62:0] _3801;
    wire [63:0] _3809;
    wire [62:0] _3810;
    wire [63:0] _3818;
    wire [62:0] _3819;
    wire [63:0] _3827;
    wire [62:0] _3828;
    wire [63:0] _3836;
    wire [62:0] _3837;
    wire [63:0] _3845;
    wire [62:0] _3846;
    wire [63:0] _3854;
    wire [62:0] _3855;
    wire [63:0] _3863;
    wire [62:0] _3864;
    wire [63:0] _3872;
    wire [62:0] _3873;
    wire [63:0] _3881;
    wire [62:0] _3882;
    wire [63:0] _3890;
    wire [62:0] _3891;
    wire [63:0] _3899;
    wire [62:0] _3900;
    wire [63:0] _3908;
    wire [62:0] _3909;
    wire [63:0] _3917;
    wire [62:0] _3918;
    wire [63:0] _3926;
    wire [62:0] _3927;
    wire [63:0] _3935;
    wire [62:0] _3936;
    wire [63:0] _3944;
    wire [62:0] _3945;
    wire [63:0] _3953;
    wire [62:0] _3954;
    wire [63:0] _3962;
    wire [62:0] _3963;
    wire [63:0] _3971;
    wire [62:0] _3972;
    wire [63:0] _3980;
    wire [62:0] _3981;
    wire [63:0] _3989;
    wire [62:0] _3990;
    wire [63:0] _3998;
    wire [62:0] _3999;
    wire [63:0] _4007;
    wire [62:0] _4008;
    wire [63:0] _4016;
    wire [62:0] _4017;
    wire [63:0] _4025;
    wire [62:0] _4026;
    wire [63:0] _4034;
    wire [62:0] _4035;
    wire [63:0] _4043;
    wire [62:0] _4044;
    wire [63:0] _4052;
    wire [62:0] _4053;
    wire [63:0] _4061;
    wire [62:0] _4062;
    wire [63:0] _4070;
    wire [62:0] _4071;
    wire [63:0] _4079;
    wire [62:0] _4080;
    wire [63:0] _4088;
    wire [127:0] _4089;
    wire [63:0] _4090;
    wire [63:0] _3511;
    wire _4091;
    wire [63:0] _4092;
    wire _3509;
    wire [63:0] _3510;
    wire _4093;
    wire _4094;
    wire [63:0] _5257;
    wire _3498;
    wire [63:0] _3495;
    wire [63:0] _3496;
    wire [62:0] _3497;
    wire [63:0] _3499;
    wire _3500;
    wire _3501;
    wire _3489;
    wire [63:0] _3486;
    wire [63:0] _3487;
    wire [62:0] _3488;
    wire [63:0] _3490;
    wire _3491;
    wire _3492;
    wire _3480;
    wire [63:0] _3477;
    wire [63:0] _3478;
    wire [62:0] _3479;
    wire [63:0] _3481;
    wire _3482;
    wire _3483;
    wire _3471;
    wire [63:0] _3468;
    wire [63:0] _3469;
    wire [62:0] _3470;
    wire [63:0] _3472;
    wire _3473;
    wire _3474;
    wire _3462;
    wire [63:0] _3459;
    wire [63:0] _3460;
    wire [62:0] _3461;
    wire [63:0] _3463;
    wire _3464;
    wire _3465;
    wire _3453;
    wire [63:0] _3450;
    wire [63:0] _3451;
    wire [62:0] _3452;
    wire [63:0] _3454;
    wire _3455;
    wire _3456;
    wire _3444;
    wire [63:0] _3441;
    wire [63:0] _3442;
    wire [62:0] _3443;
    wire [63:0] _3445;
    wire _3446;
    wire _3447;
    wire _3435;
    wire [63:0] _3432;
    wire [63:0] _3433;
    wire [62:0] _3434;
    wire [63:0] _3436;
    wire _3437;
    wire _3438;
    wire _3426;
    wire [63:0] _3423;
    wire [63:0] _3424;
    wire [62:0] _3425;
    wire [63:0] _3427;
    wire _3428;
    wire _3429;
    wire _3417;
    wire [63:0] _3414;
    wire [63:0] _3415;
    wire [62:0] _3416;
    wire [63:0] _3418;
    wire _3419;
    wire _3420;
    wire _3408;
    wire [63:0] _3405;
    wire [63:0] _3406;
    wire [62:0] _3407;
    wire [63:0] _3409;
    wire _3410;
    wire _3411;
    wire _3399;
    wire [63:0] _3396;
    wire [63:0] _3397;
    wire [62:0] _3398;
    wire [63:0] _3400;
    wire _3401;
    wire _3402;
    wire _3390;
    wire [63:0] _3387;
    wire [63:0] _3388;
    wire [62:0] _3389;
    wire [63:0] _3391;
    wire _3392;
    wire _3393;
    wire _3381;
    wire [63:0] _3378;
    wire [63:0] _3379;
    wire [62:0] _3380;
    wire [63:0] _3382;
    wire _3383;
    wire _3384;
    wire _3372;
    wire [63:0] _3369;
    wire [63:0] _3370;
    wire [62:0] _3371;
    wire [63:0] _3373;
    wire _3374;
    wire _3375;
    wire _3363;
    wire [63:0] _3360;
    wire [63:0] _3361;
    wire [62:0] _3362;
    wire [63:0] _3364;
    wire _3365;
    wire _3366;
    wire _3354;
    wire [63:0] _3351;
    wire [63:0] _3352;
    wire [62:0] _3353;
    wire [63:0] _3355;
    wire _3356;
    wire _3357;
    wire _3345;
    wire [63:0] _3342;
    wire [63:0] _3343;
    wire [62:0] _3344;
    wire [63:0] _3346;
    wire _3347;
    wire _3348;
    wire _3336;
    wire [63:0] _3333;
    wire [63:0] _3334;
    wire [62:0] _3335;
    wire [63:0] _3337;
    wire _3338;
    wire _3339;
    wire _3327;
    wire [63:0] _3324;
    wire [63:0] _3325;
    wire [62:0] _3326;
    wire [63:0] _3328;
    wire _3329;
    wire _3330;
    wire _3318;
    wire [63:0] _3315;
    wire [63:0] _3316;
    wire [62:0] _3317;
    wire [63:0] _3319;
    wire _3320;
    wire _3321;
    wire _3309;
    wire [63:0] _3306;
    wire [63:0] _3307;
    wire [62:0] _3308;
    wire [63:0] _3310;
    wire _3311;
    wire _3312;
    wire _3300;
    wire [63:0] _3297;
    wire [63:0] _3298;
    wire [62:0] _3299;
    wire [63:0] _3301;
    wire _3302;
    wire _3303;
    wire _3291;
    wire [63:0] _3288;
    wire [63:0] _3289;
    wire [62:0] _3290;
    wire [63:0] _3292;
    wire _3293;
    wire _3294;
    wire _3282;
    wire [63:0] _3279;
    wire [63:0] _3280;
    wire [62:0] _3281;
    wire [63:0] _3283;
    wire _3284;
    wire _3285;
    wire _3273;
    wire [63:0] _3270;
    wire [63:0] _3271;
    wire [62:0] _3272;
    wire [63:0] _3274;
    wire _3275;
    wire _3276;
    wire _3264;
    wire [63:0] _3261;
    wire [63:0] _3262;
    wire [62:0] _3263;
    wire [63:0] _3265;
    wire _3266;
    wire _3267;
    wire _3255;
    wire [63:0] _3252;
    wire [63:0] _3253;
    wire [62:0] _3254;
    wire [63:0] _3256;
    wire _3257;
    wire _3258;
    wire _3246;
    wire [63:0] _3243;
    wire [63:0] _3244;
    wire [62:0] _3245;
    wire [63:0] _3247;
    wire _3248;
    wire _3249;
    wire _3237;
    wire [63:0] _3234;
    wire [63:0] _3235;
    wire [62:0] _3236;
    wire [63:0] _3238;
    wire _3239;
    wire _3240;
    wire _3228;
    wire [63:0] _3225;
    wire [63:0] _3226;
    wire [62:0] _3227;
    wire [63:0] _3229;
    wire _3230;
    wire _3231;
    wire _3219;
    wire [63:0] _3216;
    wire [63:0] _3217;
    wire [62:0] _3218;
    wire [63:0] _3220;
    wire _3221;
    wire _3222;
    wire _3210;
    wire [63:0] _3207;
    wire [63:0] _3208;
    wire [62:0] _3209;
    wire [63:0] _3211;
    wire _3212;
    wire _3213;
    wire _3201;
    wire [63:0] _3198;
    wire [63:0] _3199;
    wire [62:0] _3200;
    wire [63:0] _3202;
    wire _3203;
    wire _3204;
    wire _3192;
    wire [63:0] _3189;
    wire [63:0] _3190;
    wire [62:0] _3191;
    wire [63:0] _3193;
    wire _3194;
    wire _3195;
    wire _3183;
    wire [63:0] _3180;
    wire [63:0] _3181;
    wire [62:0] _3182;
    wire [63:0] _3184;
    wire _3185;
    wire _3186;
    wire _3174;
    wire [63:0] _3171;
    wire [63:0] _3172;
    wire [62:0] _3173;
    wire [63:0] _3175;
    wire _3176;
    wire _3177;
    wire _3165;
    wire [63:0] _3162;
    wire [63:0] _3163;
    wire [62:0] _3164;
    wire [63:0] _3166;
    wire _3167;
    wire _3168;
    wire _3156;
    wire [63:0] _3153;
    wire [63:0] _3154;
    wire [62:0] _3155;
    wire [63:0] _3157;
    wire _3158;
    wire _3159;
    wire _3147;
    wire [63:0] _3144;
    wire [63:0] _3145;
    wire [62:0] _3146;
    wire [63:0] _3148;
    wire _3149;
    wire _3150;
    wire _3138;
    wire [63:0] _3135;
    wire [63:0] _3136;
    wire [62:0] _3137;
    wire [63:0] _3139;
    wire _3140;
    wire _3141;
    wire _3129;
    wire [63:0] _3126;
    wire [63:0] _3127;
    wire [62:0] _3128;
    wire [63:0] _3130;
    wire _3131;
    wire _3132;
    wire _3120;
    wire [63:0] _3117;
    wire [63:0] _3118;
    wire [62:0] _3119;
    wire [63:0] _3121;
    wire _3122;
    wire _3123;
    wire _3111;
    wire [63:0] _3108;
    wire [63:0] _3109;
    wire [62:0] _3110;
    wire [63:0] _3112;
    wire _3113;
    wire _3114;
    wire _3102;
    wire [63:0] _3099;
    wire [63:0] _3100;
    wire [62:0] _3101;
    wire [63:0] _3103;
    wire _3104;
    wire _3105;
    wire _3093;
    wire [63:0] _3090;
    wire [63:0] _3091;
    wire [62:0] _3092;
    wire [63:0] _3094;
    wire _3095;
    wire _3096;
    wire _3084;
    wire [63:0] _3081;
    wire [63:0] _3082;
    wire [62:0] _3083;
    wire [63:0] _3085;
    wire _3086;
    wire _3087;
    wire _3075;
    wire [63:0] _3072;
    wire [63:0] _3073;
    wire [62:0] _3074;
    wire [63:0] _3076;
    wire _3077;
    wire _3078;
    wire _3066;
    wire [63:0] _3063;
    wire [63:0] _3064;
    wire [62:0] _3065;
    wire [63:0] _3067;
    wire _3068;
    wire _3069;
    wire _3057;
    wire [63:0] _3054;
    wire [63:0] _3055;
    wire [62:0] _3056;
    wire [63:0] _3058;
    wire _3059;
    wire _3060;
    wire _3048;
    wire [63:0] _3045;
    wire [63:0] _3046;
    wire [62:0] _3047;
    wire [63:0] _3049;
    wire _3050;
    wire _3051;
    wire _3039;
    wire [63:0] _3036;
    wire [63:0] _3037;
    wire [62:0] _3038;
    wire [63:0] _3040;
    wire _3041;
    wire _3042;
    wire _3030;
    wire [63:0] _3027;
    wire [63:0] _3028;
    wire [62:0] _3029;
    wire [63:0] _3031;
    wire _3032;
    wire _3033;
    wire _3021;
    wire [63:0] _3018;
    wire [63:0] _3019;
    wire [62:0] _3020;
    wire [63:0] _3022;
    wire _3023;
    wire _3024;
    wire _3012;
    wire [63:0] _3009;
    wire [63:0] _3010;
    wire [62:0] _3011;
    wire [63:0] _3013;
    wire _3014;
    wire _3015;
    wire _3003;
    wire [63:0] _3000;
    wire [63:0] _3001;
    wire [62:0] _3002;
    wire [63:0] _3004;
    wire _3005;
    wire _3006;
    wire _2994;
    wire [63:0] _2991;
    wire [63:0] _2992;
    wire [62:0] _2993;
    wire [63:0] _2995;
    wire _2996;
    wire _2997;
    wire _2985;
    wire [63:0] _2982;
    wire [63:0] _2983;
    wire [62:0] _2984;
    wire [63:0] _2986;
    wire _2987;
    wire _2988;
    wire _2976;
    wire [63:0] _2973;
    wire [63:0] _2974;
    wire [62:0] _2975;
    wire [63:0] _2977;
    wire _2978;
    wire _2979;
    wire _2967;
    wire [63:0] _2964;
    wire [63:0] _2965;
    wire [62:0] _2966;
    wire [63:0] _2968;
    wire _2969;
    wire _2970;
    wire _2958;
    wire [63:0] _2955;
    wire [63:0] _2956;
    wire [62:0] _2957;
    wire [63:0] _2959;
    wire _2960;
    wire _2961;
    wire _2949;
    wire [63:0] _2946;
    wire [63:0] _2947;
    wire [62:0] _2948;
    wire [63:0] _2950;
    wire _2951;
    wire _2952;
    wire _2940;
    wire [63:0] _2937;
    wire [63:0] _2938;
    wire [62:0] _2939;
    wire [63:0] _2941;
    wire _2942;
    wire _2943;
    wire [63:0] _2927;
    wire [127:0] _2928;
    wire [63:0] _2929;
    wire _2930;
    wire [63:0] _2931;
    wire _2933;
    wire _2934;
    wire [63:0] _2935;
    wire [62:0] _2936;
    wire [63:0] _2944;
    wire [62:0] _2945;
    wire [63:0] _2953;
    wire [62:0] _2954;
    wire [63:0] _2962;
    wire [62:0] _2963;
    wire [63:0] _2971;
    wire [62:0] _2972;
    wire [63:0] _2980;
    wire [62:0] _2981;
    wire [63:0] _2989;
    wire [62:0] _2990;
    wire [63:0] _2998;
    wire [62:0] _2999;
    wire [63:0] _3007;
    wire [62:0] _3008;
    wire [63:0] _3016;
    wire [62:0] _3017;
    wire [63:0] _3025;
    wire [62:0] _3026;
    wire [63:0] _3034;
    wire [62:0] _3035;
    wire [63:0] _3043;
    wire [62:0] _3044;
    wire [63:0] _3052;
    wire [62:0] _3053;
    wire [63:0] _3061;
    wire [62:0] _3062;
    wire [63:0] _3070;
    wire [62:0] _3071;
    wire [63:0] _3079;
    wire [62:0] _3080;
    wire [63:0] _3088;
    wire [62:0] _3089;
    wire [63:0] _3097;
    wire [62:0] _3098;
    wire [63:0] _3106;
    wire [62:0] _3107;
    wire [63:0] _3115;
    wire [62:0] _3116;
    wire [63:0] _3124;
    wire [62:0] _3125;
    wire [63:0] _3133;
    wire [62:0] _3134;
    wire [63:0] _3142;
    wire [62:0] _3143;
    wire [63:0] _3151;
    wire [62:0] _3152;
    wire [63:0] _3160;
    wire [62:0] _3161;
    wire [63:0] _3169;
    wire [62:0] _3170;
    wire [63:0] _3178;
    wire [62:0] _3179;
    wire [63:0] _3187;
    wire [62:0] _3188;
    wire [63:0] _3196;
    wire [62:0] _3197;
    wire [63:0] _3205;
    wire [62:0] _3206;
    wire [63:0] _3214;
    wire [62:0] _3215;
    wire [63:0] _3223;
    wire [62:0] _3224;
    wire [63:0] _3232;
    wire [62:0] _3233;
    wire [63:0] _3241;
    wire [62:0] _3242;
    wire [63:0] _3250;
    wire [62:0] _3251;
    wire [63:0] _3259;
    wire [62:0] _3260;
    wire [63:0] _3268;
    wire [62:0] _3269;
    wire [63:0] _3277;
    wire [62:0] _3278;
    wire [63:0] _3286;
    wire [62:0] _3287;
    wire [63:0] _3295;
    wire [62:0] _3296;
    wire [63:0] _3304;
    wire [62:0] _3305;
    wire [63:0] _3313;
    wire [62:0] _3314;
    wire [63:0] _3322;
    wire [62:0] _3323;
    wire [63:0] _3331;
    wire [62:0] _3332;
    wire [63:0] _3340;
    wire [62:0] _3341;
    wire [63:0] _3349;
    wire [62:0] _3350;
    wire [63:0] _3358;
    wire [62:0] _3359;
    wire [63:0] _3367;
    wire [62:0] _3368;
    wire [63:0] _3376;
    wire [62:0] _3377;
    wire [63:0] _3385;
    wire [62:0] _3386;
    wire [63:0] _3394;
    wire [62:0] _3395;
    wire [63:0] _3403;
    wire [62:0] _3404;
    wire [63:0] _3412;
    wire [62:0] _3413;
    wire [63:0] _3421;
    wire [62:0] _3422;
    wire [63:0] _3430;
    wire [62:0] _3431;
    wire [63:0] _3439;
    wire [62:0] _3440;
    wire [63:0] _3448;
    wire [62:0] _3449;
    wire [63:0] _3457;
    wire [62:0] _3458;
    wire [63:0] _3466;
    wire [62:0] _3467;
    wire [63:0] _3475;
    wire [62:0] _3476;
    wire [63:0] _3484;
    wire [62:0] _3485;
    wire [63:0] _3493;
    wire [62:0] _3494;
    wire [63:0] _3502;
    wire [127:0] _3503;
    wire [63:0] _3504;
    wire _2915;
    wire [63:0] _2912;
    wire [63:0] _2913;
    wire [62:0] _2914;
    wire [63:0] _2916;
    wire _2917;
    wire _2918;
    wire _2906;
    wire [63:0] _2903;
    wire [63:0] _2904;
    wire [62:0] _2905;
    wire [63:0] _2907;
    wire _2908;
    wire _2909;
    wire _2897;
    wire [63:0] _2894;
    wire [63:0] _2895;
    wire [62:0] _2896;
    wire [63:0] _2898;
    wire _2899;
    wire _2900;
    wire _2888;
    wire [63:0] _2885;
    wire [63:0] _2886;
    wire [62:0] _2887;
    wire [63:0] _2889;
    wire _2890;
    wire _2891;
    wire _2879;
    wire [63:0] _2876;
    wire [63:0] _2877;
    wire [62:0] _2878;
    wire [63:0] _2880;
    wire _2881;
    wire _2882;
    wire _2870;
    wire [63:0] _2867;
    wire [63:0] _2868;
    wire [62:0] _2869;
    wire [63:0] _2871;
    wire _2872;
    wire _2873;
    wire _2861;
    wire [63:0] _2858;
    wire [63:0] _2859;
    wire [62:0] _2860;
    wire [63:0] _2862;
    wire _2863;
    wire _2864;
    wire _2852;
    wire [63:0] _2849;
    wire [63:0] _2850;
    wire [62:0] _2851;
    wire [63:0] _2853;
    wire _2854;
    wire _2855;
    wire _2843;
    wire [63:0] _2840;
    wire [63:0] _2841;
    wire [62:0] _2842;
    wire [63:0] _2844;
    wire _2845;
    wire _2846;
    wire _2834;
    wire [63:0] _2831;
    wire [63:0] _2832;
    wire [62:0] _2833;
    wire [63:0] _2835;
    wire _2836;
    wire _2837;
    wire _2825;
    wire [63:0] _2822;
    wire [63:0] _2823;
    wire [62:0] _2824;
    wire [63:0] _2826;
    wire _2827;
    wire _2828;
    wire _2816;
    wire [63:0] _2813;
    wire [63:0] _2814;
    wire [62:0] _2815;
    wire [63:0] _2817;
    wire _2818;
    wire _2819;
    wire _2807;
    wire [63:0] _2804;
    wire [63:0] _2805;
    wire [62:0] _2806;
    wire [63:0] _2808;
    wire _2809;
    wire _2810;
    wire _2798;
    wire [63:0] _2795;
    wire [63:0] _2796;
    wire [62:0] _2797;
    wire [63:0] _2799;
    wire _2800;
    wire _2801;
    wire _2789;
    wire [63:0] _2786;
    wire [63:0] _2787;
    wire [62:0] _2788;
    wire [63:0] _2790;
    wire _2791;
    wire _2792;
    wire _2780;
    wire [63:0] _2777;
    wire [63:0] _2778;
    wire [62:0] _2779;
    wire [63:0] _2781;
    wire _2782;
    wire _2783;
    wire _2771;
    wire [63:0] _2768;
    wire [63:0] _2769;
    wire [62:0] _2770;
    wire [63:0] _2772;
    wire _2773;
    wire _2774;
    wire _2762;
    wire [63:0] _2759;
    wire [63:0] _2760;
    wire [62:0] _2761;
    wire [63:0] _2763;
    wire _2764;
    wire _2765;
    wire _2753;
    wire [63:0] _2750;
    wire [63:0] _2751;
    wire [62:0] _2752;
    wire [63:0] _2754;
    wire _2755;
    wire _2756;
    wire _2744;
    wire [63:0] _2741;
    wire [63:0] _2742;
    wire [62:0] _2743;
    wire [63:0] _2745;
    wire _2746;
    wire _2747;
    wire _2735;
    wire [63:0] _2732;
    wire [63:0] _2733;
    wire [62:0] _2734;
    wire [63:0] _2736;
    wire _2737;
    wire _2738;
    wire _2726;
    wire [63:0] _2723;
    wire [63:0] _2724;
    wire [62:0] _2725;
    wire [63:0] _2727;
    wire _2728;
    wire _2729;
    wire _2717;
    wire [63:0] _2714;
    wire [63:0] _2715;
    wire [62:0] _2716;
    wire [63:0] _2718;
    wire _2719;
    wire _2720;
    wire _2708;
    wire [63:0] _2705;
    wire [63:0] _2706;
    wire [62:0] _2707;
    wire [63:0] _2709;
    wire _2710;
    wire _2711;
    wire _2699;
    wire [63:0] _2696;
    wire [63:0] _2697;
    wire [62:0] _2698;
    wire [63:0] _2700;
    wire _2701;
    wire _2702;
    wire _2690;
    wire [63:0] _2687;
    wire [63:0] _2688;
    wire [62:0] _2689;
    wire [63:0] _2691;
    wire _2692;
    wire _2693;
    wire _2681;
    wire [63:0] _2678;
    wire [63:0] _2679;
    wire [62:0] _2680;
    wire [63:0] _2682;
    wire _2683;
    wire _2684;
    wire _2672;
    wire [63:0] _2669;
    wire [63:0] _2670;
    wire [62:0] _2671;
    wire [63:0] _2673;
    wire _2674;
    wire _2675;
    wire _2663;
    wire [63:0] _2660;
    wire [63:0] _2661;
    wire [62:0] _2662;
    wire [63:0] _2664;
    wire _2665;
    wire _2666;
    wire _2654;
    wire [63:0] _2651;
    wire [63:0] _2652;
    wire [62:0] _2653;
    wire [63:0] _2655;
    wire _2656;
    wire _2657;
    wire _2645;
    wire [63:0] _2642;
    wire [63:0] _2643;
    wire [62:0] _2644;
    wire [63:0] _2646;
    wire _2647;
    wire _2648;
    wire _2636;
    wire [63:0] _2633;
    wire [63:0] _2634;
    wire [62:0] _2635;
    wire [63:0] _2637;
    wire _2638;
    wire _2639;
    wire _2627;
    wire [63:0] _2624;
    wire [63:0] _2625;
    wire [62:0] _2626;
    wire [63:0] _2628;
    wire _2629;
    wire _2630;
    wire _2618;
    wire [63:0] _2615;
    wire [63:0] _2616;
    wire [62:0] _2617;
    wire [63:0] _2619;
    wire _2620;
    wire _2621;
    wire _2609;
    wire [63:0] _2606;
    wire [63:0] _2607;
    wire [62:0] _2608;
    wire [63:0] _2610;
    wire _2611;
    wire _2612;
    wire _2600;
    wire [63:0] _2597;
    wire [63:0] _2598;
    wire [62:0] _2599;
    wire [63:0] _2601;
    wire _2602;
    wire _2603;
    wire _2591;
    wire [63:0] _2588;
    wire [63:0] _2589;
    wire [62:0] _2590;
    wire [63:0] _2592;
    wire _2593;
    wire _2594;
    wire _2582;
    wire [63:0] _2579;
    wire [63:0] _2580;
    wire [62:0] _2581;
    wire [63:0] _2583;
    wire _2584;
    wire _2585;
    wire _2573;
    wire [63:0] _2570;
    wire [63:0] _2571;
    wire [62:0] _2572;
    wire [63:0] _2574;
    wire _2575;
    wire _2576;
    wire _2564;
    wire [63:0] _2561;
    wire [63:0] _2562;
    wire [62:0] _2563;
    wire [63:0] _2565;
    wire _2566;
    wire _2567;
    wire _2555;
    wire [63:0] _2552;
    wire [63:0] _2553;
    wire [62:0] _2554;
    wire [63:0] _2556;
    wire _2557;
    wire _2558;
    wire _2546;
    wire [63:0] _2543;
    wire [63:0] _2544;
    wire [62:0] _2545;
    wire [63:0] _2547;
    wire _2548;
    wire _2549;
    wire _2537;
    wire [63:0] _2534;
    wire [63:0] _2535;
    wire [62:0] _2536;
    wire [63:0] _2538;
    wire _2539;
    wire _2540;
    wire _2528;
    wire [63:0] _2525;
    wire [63:0] _2526;
    wire [62:0] _2527;
    wire [63:0] _2529;
    wire _2530;
    wire _2531;
    wire _2519;
    wire [63:0] _2516;
    wire [63:0] _2517;
    wire [62:0] _2518;
    wire [63:0] _2520;
    wire _2521;
    wire _2522;
    wire _2510;
    wire [63:0] _2507;
    wire [63:0] _2508;
    wire [62:0] _2509;
    wire [63:0] _2511;
    wire _2512;
    wire _2513;
    wire _2501;
    wire [63:0] _2498;
    wire [63:0] _2499;
    wire [62:0] _2500;
    wire [63:0] _2502;
    wire _2503;
    wire _2504;
    wire _2492;
    wire [63:0] _2489;
    wire [63:0] _2490;
    wire [62:0] _2491;
    wire [63:0] _2493;
    wire _2494;
    wire _2495;
    wire _2483;
    wire [63:0] _2480;
    wire [63:0] _2481;
    wire [62:0] _2482;
    wire [63:0] _2484;
    wire _2485;
    wire _2486;
    wire _2474;
    wire [63:0] _2471;
    wire [63:0] _2472;
    wire [62:0] _2473;
    wire [63:0] _2475;
    wire _2476;
    wire _2477;
    wire _2465;
    wire [63:0] _2462;
    wire [63:0] _2463;
    wire [62:0] _2464;
    wire [63:0] _2466;
    wire _2467;
    wire _2468;
    wire _2456;
    wire [63:0] _2453;
    wire [63:0] _2454;
    wire [62:0] _2455;
    wire [63:0] _2457;
    wire _2458;
    wire _2459;
    wire _2447;
    wire [63:0] _2444;
    wire [63:0] _2445;
    wire [62:0] _2446;
    wire [63:0] _2448;
    wire _2449;
    wire _2450;
    wire _2438;
    wire [63:0] _2435;
    wire [63:0] _2436;
    wire [62:0] _2437;
    wire [63:0] _2439;
    wire _2440;
    wire _2441;
    wire _2429;
    wire [63:0] _2426;
    wire [63:0] _2427;
    wire [62:0] _2428;
    wire [63:0] _2430;
    wire _2431;
    wire _2432;
    wire _2420;
    wire [63:0] _2417;
    wire [63:0] _2418;
    wire [62:0] _2419;
    wire [63:0] _2421;
    wire _2422;
    wire _2423;
    wire _2411;
    wire [63:0] _2408;
    wire [63:0] _2409;
    wire [62:0] _2410;
    wire [63:0] _2412;
    wire _2413;
    wire _2414;
    wire _2402;
    wire [63:0] _2399;
    wire [63:0] _2400;
    wire [62:0] _2401;
    wire [63:0] _2403;
    wire _2404;
    wire _2405;
    wire _2393;
    wire [63:0] _2390;
    wire [63:0] _2391;
    wire [62:0] _2392;
    wire [63:0] _2394;
    wire _2395;
    wire _2396;
    wire _2384;
    wire [63:0] _2381;
    wire [63:0] _2382;
    wire [62:0] _2383;
    wire [63:0] _2385;
    wire _2386;
    wire _2387;
    wire _2375;
    wire [63:0] _2372;
    wire [63:0] _2373;
    wire [62:0] _2374;
    wire [63:0] _2376;
    wire _2377;
    wire _2378;
    wire _2366;
    wire [63:0] _2363;
    wire [63:0] _2364;
    wire [62:0] _2365;
    wire [63:0] _2367;
    wire _2368;
    wire _2369;
    wire _2357;
    wire [63:0] _2354;
    wire [63:0] _2355;
    wire [62:0] _2356;
    wire [63:0] _2358;
    wire _2359;
    wire _2360;
    wire [63:0] _2347;
    wire _2348;
    wire [63:0] _2349;
    wire _2350;
    wire _2351;
    wire [63:0] _2352;
    wire [62:0] _2353;
    wire [63:0] _2361;
    wire [62:0] _2362;
    wire [63:0] _2370;
    wire [62:0] _2371;
    wire [63:0] _2379;
    wire [62:0] _2380;
    wire [63:0] _2388;
    wire [62:0] _2389;
    wire [63:0] _2397;
    wire [62:0] _2398;
    wire [63:0] _2406;
    wire [62:0] _2407;
    wire [63:0] _2415;
    wire [62:0] _2416;
    wire [63:0] _2424;
    wire [62:0] _2425;
    wire [63:0] _2433;
    wire [62:0] _2434;
    wire [63:0] _2442;
    wire [62:0] _2443;
    wire [63:0] _2451;
    wire [62:0] _2452;
    wire [63:0] _2460;
    wire [62:0] _2461;
    wire [63:0] _2469;
    wire [62:0] _2470;
    wire [63:0] _2478;
    wire [62:0] _2479;
    wire [63:0] _2487;
    wire [62:0] _2488;
    wire [63:0] _2496;
    wire [62:0] _2497;
    wire [63:0] _2505;
    wire [62:0] _2506;
    wire [63:0] _2514;
    wire [62:0] _2515;
    wire [63:0] _2523;
    wire [62:0] _2524;
    wire [63:0] _2532;
    wire [62:0] _2533;
    wire [63:0] _2541;
    wire [62:0] _2542;
    wire [63:0] _2550;
    wire [62:0] _2551;
    wire [63:0] _2559;
    wire [62:0] _2560;
    wire [63:0] _2568;
    wire [62:0] _2569;
    wire [63:0] _2577;
    wire [62:0] _2578;
    wire [63:0] _2586;
    wire [62:0] _2587;
    wire [63:0] _2595;
    wire [62:0] _2596;
    wire [63:0] _2604;
    wire [62:0] _2605;
    wire [63:0] _2613;
    wire [62:0] _2614;
    wire [63:0] _2622;
    wire [62:0] _2623;
    wire [63:0] _2631;
    wire [62:0] _2632;
    wire [63:0] _2640;
    wire [62:0] _2641;
    wire [63:0] _2649;
    wire [62:0] _2650;
    wire [63:0] _2658;
    wire [62:0] _2659;
    wire [63:0] _2667;
    wire [62:0] _2668;
    wire [63:0] _2676;
    wire [62:0] _2677;
    wire [63:0] _2685;
    wire [62:0] _2686;
    wire [63:0] _2694;
    wire [62:0] _2695;
    wire [63:0] _2703;
    wire [62:0] _2704;
    wire [63:0] _2712;
    wire [62:0] _2713;
    wire [63:0] _2721;
    wire [62:0] _2722;
    wire [63:0] _2730;
    wire [62:0] _2731;
    wire [63:0] _2739;
    wire [62:0] _2740;
    wire [63:0] _2748;
    wire [62:0] _2749;
    wire [63:0] _2757;
    wire [62:0] _2758;
    wire [63:0] _2766;
    wire [62:0] _2767;
    wire [63:0] _2775;
    wire [62:0] _2776;
    wire [63:0] _2784;
    wire [62:0] _2785;
    wire [63:0] _2793;
    wire [62:0] _2794;
    wire [63:0] _2802;
    wire [62:0] _2803;
    wire [63:0] _2811;
    wire [62:0] _2812;
    wire [63:0] _2820;
    wire [62:0] _2821;
    wire [63:0] _2829;
    wire [62:0] _2830;
    wire [63:0] _2838;
    wire [62:0] _2839;
    wire [63:0] _2847;
    wire [62:0] _2848;
    wire [63:0] _2856;
    wire [62:0] _2857;
    wire [63:0] _2865;
    wire [62:0] _2866;
    wire [63:0] _2874;
    wire [62:0] _2875;
    wire [63:0] _2883;
    wire [62:0] _2884;
    wire [63:0] _2892;
    wire [62:0] _2893;
    wire [63:0] _2901;
    wire [62:0] _2902;
    wire [63:0] _2910;
    wire [62:0] _2911;
    wire [63:0] _2919;
    wire [63:0] _2921;
    wire [127:0] _2922;
    wire [63:0] _2923;
    wire [63:0] _3505;
    wire _2333;
    wire [63:0] _2330;
    wire [63:0] _2331;
    wire [62:0] _2332;
    wire [63:0] _2334;
    wire _2335;
    wire _2336;
    wire _2324;
    wire [63:0] _2321;
    wire [63:0] _2322;
    wire [62:0] _2323;
    wire [63:0] _2325;
    wire _2326;
    wire _2327;
    wire _2315;
    wire [63:0] _2312;
    wire [63:0] _2313;
    wire [62:0] _2314;
    wire [63:0] _2316;
    wire _2317;
    wire _2318;
    wire _2306;
    wire [63:0] _2303;
    wire [63:0] _2304;
    wire [62:0] _2305;
    wire [63:0] _2307;
    wire _2308;
    wire _2309;
    wire _2297;
    wire [63:0] _2294;
    wire [63:0] _2295;
    wire [62:0] _2296;
    wire [63:0] _2298;
    wire _2299;
    wire _2300;
    wire _2288;
    wire [63:0] _2285;
    wire [63:0] _2286;
    wire [62:0] _2287;
    wire [63:0] _2289;
    wire _2290;
    wire _2291;
    wire _2279;
    wire [63:0] _2276;
    wire [63:0] _2277;
    wire [62:0] _2278;
    wire [63:0] _2280;
    wire _2281;
    wire _2282;
    wire _2270;
    wire [63:0] _2267;
    wire [63:0] _2268;
    wire [62:0] _2269;
    wire [63:0] _2271;
    wire _2272;
    wire _2273;
    wire _2261;
    wire [63:0] _2258;
    wire [63:0] _2259;
    wire [62:0] _2260;
    wire [63:0] _2262;
    wire _2263;
    wire _2264;
    wire _2252;
    wire [63:0] _2249;
    wire [63:0] _2250;
    wire [62:0] _2251;
    wire [63:0] _2253;
    wire _2254;
    wire _2255;
    wire _2243;
    wire [63:0] _2240;
    wire [63:0] _2241;
    wire [62:0] _2242;
    wire [63:0] _2244;
    wire _2245;
    wire _2246;
    wire _2234;
    wire [63:0] _2231;
    wire [63:0] _2232;
    wire [62:0] _2233;
    wire [63:0] _2235;
    wire _2236;
    wire _2237;
    wire _2225;
    wire [63:0] _2222;
    wire [63:0] _2223;
    wire [62:0] _2224;
    wire [63:0] _2226;
    wire _2227;
    wire _2228;
    wire _2216;
    wire [63:0] _2213;
    wire [63:0] _2214;
    wire [62:0] _2215;
    wire [63:0] _2217;
    wire _2218;
    wire _2219;
    wire _2207;
    wire [63:0] _2204;
    wire [63:0] _2205;
    wire [62:0] _2206;
    wire [63:0] _2208;
    wire _2209;
    wire _2210;
    wire _2198;
    wire [63:0] _2195;
    wire [63:0] _2196;
    wire [62:0] _2197;
    wire [63:0] _2199;
    wire _2200;
    wire _2201;
    wire _2189;
    wire [63:0] _2186;
    wire [63:0] _2187;
    wire [62:0] _2188;
    wire [63:0] _2190;
    wire _2191;
    wire _2192;
    wire _2180;
    wire [63:0] _2177;
    wire [63:0] _2178;
    wire [62:0] _2179;
    wire [63:0] _2181;
    wire _2182;
    wire _2183;
    wire _2171;
    wire [63:0] _2168;
    wire [63:0] _2169;
    wire [62:0] _2170;
    wire [63:0] _2172;
    wire _2173;
    wire _2174;
    wire _2162;
    wire [63:0] _2159;
    wire [63:0] _2160;
    wire [62:0] _2161;
    wire [63:0] _2163;
    wire _2164;
    wire _2165;
    wire _2153;
    wire [63:0] _2150;
    wire [63:0] _2151;
    wire [62:0] _2152;
    wire [63:0] _2154;
    wire _2155;
    wire _2156;
    wire _2144;
    wire [63:0] _2141;
    wire [63:0] _2142;
    wire [62:0] _2143;
    wire [63:0] _2145;
    wire _2146;
    wire _2147;
    wire _2135;
    wire [63:0] _2132;
    wire [63:0] _2133;
    wire [62:0] _2134;
    wire [63:0] _2136;
    wire _2137;
    wire _2138;
    wire _2126;
    wire [63:0] _2123;
    wire [63:0] _2124;
    wire [62:0] _2125;
    wire [63:0] _2127;
    wire _2128;
    wire _2129;
    wire _2117;
    wire [63:0] _2114;
    wire [63:0] _2115;
    wire [62:0] _2116;
    wire [63:0] _2118;
    wire _2119;
    wire _2120;
    wire _2108;
    wire [63:0] _2105;
    wire [63:0] _2106;
    wire [62:0] _2107;
    wire [63:0] _2109;
    wire _2110;
    wire _2111;
    wire _2099;
    wire [63:0] _2096;
    wire [63:0] _2097;
    wire [62:0] _2098;
    wire [63:0] _2100;
    wire _2101;
    wire _2102;
    wire _2090;
    wire [63:0] _2087;
    wire [63:0] _2088;
    wire [62:0] _2089;
    wire [63:0] _2091;
    wire _2092;
    wire _2093;
    wire _2081;
    wire [63:0] _2078;
    wire [63:0] _2079;
    wire [62:0] _2080;
    wire [63:0] _2082;
    wire _2083;
    wire _2084;
    wire _2072;
    wire [63:0] _2069;
    wire [63:0] _2070;
    wire [62:0] _2071;
    wire [63:0] _2073;
    wire _2074;
    wire _2075;
    wire _2063;
    wire [63:0] _2060;
    wire [63:0] _2061;
    wire [62:0] _2062;
    wire [63:0] _2064;
    wire _2065;
    wire _2066;
    wire _2054;
    wire [63:0] _2051;
    wire [63:0] _2052;
    wire [62:0] _2053;
    wire [63:0] _2055;
    wire _2056;
    wire _2057;
    wire _2045;
    wire [63:0] _2042;
    wire [63:0] _2043;
    wire [62:0] _2044;
    wire [63:0] _2046;
    wire _2047;
    wire _2048;
    wire _2036;
    wire [63:0] _2033;
    wire [63:0] _2034;
    wire [62:0] _2035;
    wire [63:0] _2037;
    wire _2038;
    wire _2039;
    wire _2027;
    wire [63:0] _2024;
    wire [63:0] _2025;
    wire [62:0] _2026;
    wire [63:0] _2028;
    wire _2029;
    wire _2030;
    wire _2018;
    wire [63:0] _2015;
    wire [63:0] _2016;
    wire [62:0] _2017;
    wire [63:0] _2019;
    wire _2020;
    wire _2021;
    wire _2009;
    wire [63:0] _2006;
    wire [63:0] _2007;
    wire [62:0] _2008;
    wire [63:0] _2010;
    wire _2011;
    wire _2012;
    wire _2000;
    wire [63:0] _1997;
    wire [63:0] _1998;
    wire [62:0] _1999;
    wire [63:0] _2001;
    wire _2002;
    wire _2003;
    wire _1991;
    wire [63:0] _1988;
    wire [63:0] _1989;
    wire [62:0] _1990;
    wire [63:0] _1992;
    wire _1993;
    wire _1994;
    wire _1982;
    wire [63:0] _1979;
    wire [63:0] _1980;
    wire [62:0] _1981;
    wire [63:0] _1983;
    wire _1984;
    wire _1985;
    wire _1973;
    wire [63:0] _1970;
    wire [63:0] _1971;
    wire [62:0] _1972;
    wire [63:0] _1974;
    wire _1975;
    wire _1976;
    wire _1964;
    wire [63:0] _1961;
    wire [63:0] _1962;
    wire [62:0] _1963;
    wire [63:0] _1965;
    wire _1966;
    wire _1967;
    wire _1955;
    wire [63:0] _1952;
    wire [63:0] _1953;
    wire [62:0] _1954;
    wire [63:0] _1956;
    wire _1957;
    wire _1958;
    wire _1946;
    wire [63:0] _1943;
    wire [63:0] _1944;
    wire [62:0] _1945;
    wire [63:0] _1947;
    wire _1948;
    wire _1949;
    wire _1937;
    wire [63:0] _1934;
    wire [63:0] _1935;
    wire [62:0] _1936;
    wire [63:0] _1938;
    wire _1939;
    wire _1940;
    wire _1928;
    wire [63:0] _1925;
    wire [63:0] _1926;
    wire [62:0] _1927;
    wire [63:0] _1929;
    wire _1930;
    wire _1931;
    wire _1919;
    wire [63:0] _1916;
    wire [63:0] _1917;
    wire [62:0] _1918;
    wire [63:0] _1920;
    wire _1921;
    wire _1922;
    wire _1910;
    wire [63:0] _1907;
    wire [63:0] _1908;
    wire [62:0] _1909;
    wire [63:0] _1911;
    wire _1912;
    wire _1913;
    wire _1901;
    wire [63:0] _1898;
    wire [63:0] _1899;
    wire [62:0] _1900;
    wire [63:0] _1902;
    wire _1903;
    wire _1904;
    wire _1892;
    wire [63:0] _1889;
    wire [63:0] _1890;
    wire [62:0] _1891;
    wire [63:0] _1893;
    wire _1894;
    wire _1895;
    wire _1883;
    wire [63:0] _1880;
    wire [63:0] _1881;
    wire [62:0] _1882;
    wire [63:0] _1884;
    wire _1885;
    wire _1886;
    wire _1874;
    wire [63:0] _1871;
    wire [63:0] _1872;
    wire [62:0] _1873;
    wire [63:0] _1875;
    wire _1876;
    wire _1877;
    wire _1865;
    wire [63:0] _1862;
    wire [63:0] _1863;
    wire [62:0] _1864;
    wire [63:0] _1866;
    wire _1867;
    wire _1868;
    wire _1856;
    wire [63:0] _1853;
    wire [63:0] _1854;
    wire [62:0] _1855;
    wire [63:0] _1857;
    wire _1858;
    wire _1859;
    wire _1847;
    wire [63:0] _1844;
    wire [63:0] _1845;
    wire [62:0] _1846;
    wire [63:0] _1848;
    wire _1849;
    wire _1850;
    wire _1838;
    wire [63:0] _1835;
    wire [63:0] _1836;
    wire [62:0] _1837;
    wire [63:0] _1839;
    wire _1840;
    wire _1841;
    wire _1829;
    wire [63:0] _1826;
    wire [63:0] _1827;
    wire [62:0] _1828;
    wire [63:0] _1830;
    wire _1831;
    wire _1832;
    wire _1820;
    wire [63:0] _1817;
    wire [63:0] _1818;
    wire [62:0] _1819;
    wire [63:0] _1821;
    wire _1822;
    wire _1823;
    wire _1811;
    wire [63:0] _1808;
    wire [63:0] _1809;
    wire [62:0] _1810;
    wire [63:0] _1812;
    wire _1813;
    wire _1814;
    wire _1802;
    wire [63:0] _1799;
    wire [63:0] _1800;
    wire [62:0] _1801;
    wire [63:0] _1803;
    wire _1804;
    wire _1805;
    wire _1793;
    wire [63:0] _1790;
    wire [63:0] _1791;
    wire [62:0] _1792;
    wire [63:0] _1794;
    wire _1795;
    wire _1796;
    wire _1784;
    wire [63:0] _1781;
    wire [63:0] _1782;
    wire [62:0] _1783;
    wire [63:0] _1785;
    wire _1786;
    wire _1787;
    wire _1775;
    wire [63:0] _1772;
    wire [63:0] _1773;
    wire [62:0] _1774;
    wire [63:0] _1776;
    wire _1777;
    wire _1778;
    wire [63:0] _1767;
    wire [63:0] _1763;
    wire [63:0] _1764;
    wire _1765;
    wire [63:0] _1766;
    wire _1768;
    wire _1769;
    wire [63:0] _1770;
    wire [62:0] _1771;
    wire [63:0] _1779;
    wire [62:0] _1780;
    wire [63:0] _1788;
    wire [62:0] _1789;
    wire [63:0] _1797;
    wire [62:0] _1798;
    wire [63:0] _1806;
    wire [62:0] _1807;
    wire [63:0] _1815;
    wire [62:0] _1816;
    wire [63:0] _1824;
    wire [62:0] _1825;
    wire [63:0] _1833;
    wire [62:0] _1834;
    wire [63:0] _1842;
    wire [62:0] _1843;
    wire [63:0] _1851;
    wire [62:0] _1852;
    wire [63:0] _1860;
    wire [62:0] _1861;
    wire [63:0] _1869;
    wire [62:0] _1870;
    wire [63:0] _1878;
    wire [62:0] _1879;
    wire [63:0] _1887;
    wire [62:0] _1888;
    wire [63:0] _1896;
    wire [62:0] _1897;
    wire [63:0] _1905;
    wire [62:0] _1906;
    wire [63:0] _1914;
    wire [62:0] _1915;
    wire [63:0] _1923;
    wire [62:0] _1924;
    wire [63:0] _1932;
    wire [62:0] _1933;
    wire [63:0] _1941;
    wire [62:0] _1942;
    wire [63:0] _1950;
    wire [62:0] _1951;
    wire [63:0] _1959;
    wire [62:0] _1960;
    wire [63:0] _1968;
    wire [62:0] _1969;
    wire [63:0] _1977;
    wire [62:0] _1978;
    wire [63:0] _1986;
    wire [62:0] _1987;
    wire [63:0] _1995;
    wire [62:0] _1996;
    wire [63:0] _2004;
    wire [62:0] _2005;
    wire [63:0] _2013;
    wire [62:0] _2014;
    wire [63:0] _2022;
    wire [62:0] _2023;
    wire [63:0] _2031;
    wire [62:0] _2032;
    wire [63:0] _2040;
    wire [62:0] _2041;
    wire [63:0] _2049;
    wire [62:0] _2050;
    wire [63:0] _2058;
    wire [62:0] _2059;
    wire [63:0] _2067;
    wire [62:0] _2068;
    wire [63:0] _2076;
    wire [62:0] _2077;
    wire [63:0] _2085;
    wire [62:0] _2086;
    wire [63:0] _2094;
    wire [62:0] _2095;
    wire [63:0] _2103;
    wire [62:0] _2104;
    wire [63:0] _2112;
    wire [62:0] _2113;
    wire [63:0] _2121;
    wire [62:0] _2122;
    wire [63:0] _2130;
    wire [62:0] _2131;
    wire [63:0] _2139;
    wire [62:0] _2140;
    wire [63:0] _2148;
    wire [62:0] _2149;
    wire [63:0] _2157;
    wire [62:0] _2158;
    wire [63:0] _2166;
    wire [62:0] _2167;
    wire [63:0] _2175;
    wire [62:0] _2176;
    wire [63:0] _2184;
    wire [62:0] _2185;
    wire [63:0] _2193;
    wire [62:0] _2194;
    wire [63:0] _2202;
    wire [62:0] _2203;
    wire [63:0] _2211;
    wire [62:0] _2212;
    wire [63:0] _2220;
    wire [62:0] _2221;
    wire [63:0] _2229;
    wire [62:0] _2230;
    wire [63:0] _2238;
    wire [62:0] _2239;
    wire [63:0] _2247;
    wire [62:0] _2248;
    wire [63:0] _2256;
    wire [62:0] _2257;
    wire [63:0] _2265;
    wire [62:0] _2266;
    wire [63:0] _2274;
    wire [62:0] _2275;
    wire [63:0] _2283;
    wire [62:0] _2284;
    wire [63:0] _2292;
    wire [62:0] _2293;
    wire [63:0] _2301;
    wire [62:0] _2302;
    wire [63:0] _2310;
    wire [62:0] _2311;
    wire [63:0] _2319;
    wire [62:0] _2320;
    wire [63:0] _2328;
    wire [62:0] _2329;
    wire [63:0] _2337;
    wire [127:0] _2338;
    wire [63:0] _2339;
    wire [63:0] _1760;
    wire _2340;
    wire [63:0] _2341;
    wire [63:0] _1757;
    wire _1758;
    wire [63:0] _1759;
    wire _2342;
    wire _2343;
    wire [63:0] _3506;
    wire _1748;
    wire [63:0] _1745;
    wire [63:0] _1746;
    wire [62:0] _1747;
    wire [63:0] _1749;
    wire _1750;
    wire _1751;
    wire _1739;
    wire [63:0] _1736;
    wire [63:0] _1737;
    wire [62:0] _1738;
    wire [63:0] _1740;
    wire _1741;
    wire _1742;
    wire _1730;
    wire [63:0] _1727;
    wire [63:0] _1728;
    wire [62:0] _1729;
    wire [63:0] _1731;
    wire _1732;
    wire _1733;
    wire _1721;
    wire [63:0] _1718;
    wire [63:0] _1719;
    wire [62:0] _1720;
    wire [63:0] _1722;
    wire _1723;
    wire _1724;
    wire _1712;
    wire [63:0] _1709;
    wire [63:0] _1710;
    wire [62:0] _1711;
    wire [63:0] _1713;
    wire _1714;
    wire _1715;
    wire _1703;
    wire [63:0] _1700;
    wire [63:0] _1701;
    wire [62:0] _1702;
    wire [63:0] _1704;
    wire _1705;
    wire _1706;
    wire _1694;
    wire [63:0] _1691;
    wire [63:0] _1692;
    wire [62:0] _1693;
    wire [63:0] _1695;
    wire _1696;
    wire _1697;
    wire _1685;
    wire [63:0] _1682;
    wire [63:0] _1683;
    wire [62:0] _1684;
    wire [63:0] _1686;
    wire _1687;
    wire _1688;
    wire _1676;
    wire [63:0] _1673;
    wire [63:0] _1674;
    wire [62:0] _1675;
    wire [63:0] _1677;
    wire _1678;
    wire _1679;
    wire _1667;
    wire [63:0] _1664;
    wire [63:0] _1665;
    wire [62:0] _1666;
    wire [63:0] _1668;
    wire _1669;
    wire _1670;
    wire _1658;
    wire [63:0] _1655;
    wire [63:0] _1656;
    wire [62:0] _1657;
    wire [63:0] _1659;
    wire _1660;
    wire _1661;
    wire _1649;
    wire [63:0] _1646;
    wire [63:0] _1647;
    wire [62:0] _1648;
    wire [63:0] _1650;
    wire _1651;
    wire _1652;
    wire _1640;
    wire [63:0] _1637;
    wire [63:0] _1638;
    wire [62:0] _1639;
    wire [63:0] _1641;
    wire _1642;
    wire _1643;
    wire _1631;
    wire [63:0] _1628;
    wire [63:0] _1629;
    wire [62:0] _1630;
    wire [63:0] _1632;
    wire _1633;
    wire _1634;
    wire _1622;
    wire [63:0] _1619;
    wire [63:0] _1620;
    wire [62:0] _1621;
    wire [63:0] _1623;
    wire _1624;
    wire _1625;
    wire _1613;
    wire [63:0] _1610;
    wire [63:0] _1611;
    wire [62:0] _1612;
    wire [63:0] _1614;
    wire _1615;
    wire _1616;
    wire _1604;
    wire [63:0] _1601;
    wire [63:0] _1602;
    wire [62:0] _1603;
    wire [63:0] _1605;
    wire _1606;
    wire _1607;
    wire _1595;
    wire [63:0] _1592;
    wire [63:0] _1593;
    wire [62:0] _1594;
    wire [63:0] _1596;
    wire _1597;
    wire _1598;
    wire _1586;
    wire [63:0] _1583;
    wire [63:0] _1584;
    wire [62:0] _1585;
    wire [63:0] _1587;
    wire _1588;
    wire _1589;
    wire _1577;
    wire [63:0] _1574;
    wire [63:0] _1575;
    wire [62:0] _1576;
    wire [63:0] _1578;
    wire _1579;
    wire _1580;
    wire _1568;
    wire [63:0] _1565;
    wire [63:0] _1566;
    wire [62:0] _1567;
    wire [63:0] _1569;
    wire _1570;
    wire _1571;
    wire _1559;
    wire [63:0] _1556;
    wire [63:0] _1557;
    wire [62:0] _1558;
    wire [63:0] _1560;
    wire _1561;
    wire _1562;
    wire _1550;
    wire [63:0] _1547;
    wire [63:0] _1548;
    wire [62:0] _1549;
    wire [63:0] _1551;
    wire _1552;
    wire _1553;
    wire _1541;
    wire [63:0] _1538;
    wire [63:0] _1539;
    wire [62:0] _1540;
    wire [63:0] _1542;
    wire _1543;
    wire _1544;
    wire _1532;
    wire [63:0] _1529;
    wire [63:0] _1530;
    wire [62:0] _1531;
    wire [63:0] _1533;
    wire _1534;
    wire _1535;
    wire _1523;
    wire [63:0] _1520;
    wire [63:0] _1521;
    wire [62:0] _1522;
    wire [63:0] _1524;
    wire _1525;
    wire _1526;
    wire _1514;
    wire [63:0] _1511;
    wire [63:0] _1512;
    wire [62:0] _1513;
    wire [63:0] _1515;
    wire _1516;
    wire _1517;
    wire _1505;
    wire [63:0] _1502;
    wire [63:0] _1503;
    wire [62:0] _1504;
    wire [63:0] _1506;
    wire _1507;
    wire _1508;
    wire _1496;
    wire [63:0] _1493;
    wire [63:0] _1494;
    wire [62:0] _1495;
    wire [63:0] _1497;
    wire _1498;
    wire _1499;
    wire _1487;
    wire [63:0] _1484;
    wire [63:0] _1485;
    wire [62:0] _1486;
    wire [63:0] _1488;
    wire _1489;
    wire _1490;
    wire _1478;
    wire [63:0] _1475;
    wire [63:0] _1476;
    wire [62:0] _1477;
    wire [63:0] _1479;
    wire _1480;
    wire _1481;
    wire _1469;
    wire [63:0] _1466;
    wire [63:0] _1467;
    wire [62:0] _1468;
    wire [63:0] _1470;
    wire _1471;
    wire _1472;
    wire _1460;
    wire [63:0] _1457;
    wire [63:0] _1458;
    wire [62:0] _1459;
    wire [63:0] _1461;
    wire _1462;
    wire _1463;
    wire _1451;
    wire [63:0] _1448;
    wire [63:0] _1449;
    wire [62:0] _1450;
    wire [63:0] _1452;
    wire _1453;
    wire _1454;
    wire _1442;
    wire [63:0] _1439;
    wire [63:0] _1440;
    wire [62:0] _1441;
    wire [63:0] _1443;
    wire _1444;
    wire _1445;
    wire _1433;
    wire [63:0] _1430;
    wire [63:0] _1431;
    wire [62:0] _1432;
    wire [63:0] _1434;
    wire _1435;
    wire _1436;
    wire _1424;
    wire [63:0] _1421;
    wire [63:0] _1422;
    wire [62:0] _1423;
    wire [63:0] _1425;
    wire _1426;
    wire _1427;
    wire _1415;
    wire [63:0] _1412;
    wire [63:0] _1413;
    wire [62:0] _1414;
    wire [63:0] _1416;
    wire _1417;
    wire _1418;
    wire _1406;
    wire [63:0] _1403;
    wire [63:0] _1404;
    wire [62:0] _1405;
    wire [63:0] _1407;
    wire _1408;
    wire _1409;
    wire _1397;
    wire [63:0] _1394;
    wire [63:0] _1395;
    wire [62:0] _1396;
    wire [63:0] _1398;
    wire _1399;
    wire _1400;
    wire _1388;
    wire [63:0] _1385;
    wire [63:0] _1386;
    wire [62:0] _1387;
    wire [63:0] _1389;
    wire _1390;
    wire _1391;
    wire _1379;
    wire [63:0] _1376;
    wire [63:0] _1377;
    wire [62:0] _1378;
    wire [63:0] _1380;
    wire _1381;
    wire _1382;
    wire _1370;
    wire [63:0] _1367;
    wire [63:0] _1368;
    wire [62:0] _1369;
    wire [63:0] _1371;
    wire _1372;
    wire _1373;
    wire _1361;
    wire [63:0] _1358;
    wire [63:0] _1359;
    wire [62:0] _1360;
    wire [63:0] _1362;
    wire _1363;
    wire _1364;
    wire _1352;
    wire [63:0] _1349;
    wire [63:0] _1350;
    wire [62:0] _1351;
    wire [63:0] _1353;
    wire _1354;
    wire _1355;
    wire _1343;
    wire [63:0] _1340;
    wire [63:0] _1341;
    wire [62:0] _1342;
    wire [63:0] _1344;
    wire _1345;
    wire _1346;
    wire _1334;
    wire [63:0] _1331;
    wire [63:0] _1332;
    wire [62:0] _1333;
    wire [63:0] _1335;
    wire _1336;
    wire _1337;
    wire _1325;
    wire [63:0] _1322;
    wire [63:0] _1323;
    wire [62:0] _1324;
    wire [63:0] _1326;
    wire _1327;
    wire _1328;
    wire _1316;
    wire [63:0] _1313;
    wire [63:0] _1314;
    wire [62:0] _1315;
    wire [63:0] _1317;
    wire _1318;
    wire _1319;
    wire _1307;
    wire [63:0] _1304;
    wire [63:0] _1305;
    wire [62:0] _1306;
    wire [63:0] _1308;
    wire _1309;
    wire _1310;
    wire _1298;
    wire [63:0] _1295;
    wire [63:0] _1296;
    wire [62:0] _1297;
    wire [63:0] _1299;
    wire _1300;
    wire _1301;
    wire _1289;
    wire [63:0] _1286;
    wire [63:0] _1287;
    wire [62:0] _1288;
    wire [63:0] _1290;
    wire _1291;
    wire _1292;
    wire _1280;
    wire [63:0] _1277;
    wire [63:0] _1278;
    wire [62:0] _1279;
    wire [63:0] _1281;
    wire _1282;
    wire _1283;
    wire _1271;
    wire [63:0] _1268;
    wire [63:0] _1269;
    wire [62:0] _1270;
    wire [63:0] _1272;
    wire _1273;
    wire _1274;
    wire _1262;
    wire [63:0] _1259;
    wire [63:0] _1260;
    wire [62:0] _1261;
    wire [63:0] _1263;
    wire _1264;
    wire _1265;
    wire _1253;
    wire [63:0] _1250;
    wire [63:0] _1251;
    wire [62:0] _1252;
    wire [63:0] _1254;
    wire _1255;
    wire _1256;
    wire _1244;
    wire [63:0] _1241;
    wire [63:0] _1242;
    wire [62:0] _1243;
    wire [63:0] _1245;
    wire _1246;
    wire _1247;
    wire _1235;
    wire [63:0] _1232;
    wire [63:0] _1233;
    wire [62:0] _1234;
    wire [63:0] _1236;
    wire _1237;
    wire _1238;
    wire _1226;
    wire [63:0] _1223;
    wire [63:0] _1224;
    wire [62:0] _1225;
    wire [63:0] _1227;
    wire _1228;
    wire _1229;
    wire _1217;
    wire [63:0] _1214;
    wire [63:0] _1215;
    wire [62:0] _1216;
    wire [63:0] _1218;
    wire _1219;
    wire _1220;
    wire _1208;
    wire [63:0] _1205;
    wire [63:0] _1206;
    wire [62:0] _1207;
    wire [63:0] _1209;
    wire _1210;
    wire _1211;
    wire _1199;
    wire [63:0] _1196;
    wire [63:0] _1197;
    wire [62:0] _1198;
    wire [63:0] _1200;
    wire _1201;
    wire _1202;
    wire _1190;
    wire [63:0] _1187;
    wire [63:0] _1188;
    wire [62:0] _1189;
    wire [63:0] _1191;
    wire _1192;
    wire _1193;
    wire [63:0] _1177;
    wire [127:0] _1178;
    wire [63:0] _1179;
    wire _1180;
    wire [63:0] _1181;
    wire _1183;
    wire _1184;
    wire [63:0] _1185;
    wire [62:0] _1186;
    wire [63:0] _1194;
    wire [62:0] _1195;
    wire [63:0] _1203;
    wire [62:0] _1204;
    wire [63:0] _1212;
    wire [62:0] _1213;
    wire [63:0] _1221;
    wire [62:0] _1222;
    wire [63:0] _1230;
    wire [62:0] _1231;
    wire [63:0] _1239;
    wire [62:0] _1240;
    wire [63:0] _1248;
    wire [62:0] _1249;
    wire [63:0] _1257;
    wire [62:0] _1258;
    wire [63:0] _1266;
    wire [62:0] _1267;
    wire [63:0] _1275;
    wire [62:0] _1276;
    wire [63:0] _1284;
    wire [62:0] _1285;
    wire [63:0] _1293;
    wire [62:0] _1294;
    wire [63:0] _1302;
    wire [62:0] _1303;
    wire [63:0] _1311;
    wire [62:0] _1312;
    wire [63:0] _1320;
    wire [62:0] _1321;
    wire [63:0] _1329;
    wire [62:0] _1330;
    wire [63:0] _1338;
    wire [62:0] _1339;
    wire [63:0] _1347;
    wire [62:0] _1348;
    wire [63:0] _1356;
    wire [62:0] _1357;
    wire [63:0] _1365;
    wire [62:0] _1366;
    wire [63:0] _1374;
    wire [62:0] _1375;
    wire [63:0] _1383;
    wire [62:0] _1384;
    wire [63:0] _1392;
    wire [62:0] _1393;
    wire [63:0] _1401;
    wire [62:0] _1402;
    wire [63:0] _1410;
    wire [62:0] _1411;
    wire [63:0] _1419;
    wire [62:0] _1420;
    wire [63:0] _1428;
    wire [62:0] _1429;
    wire [63:0] _1437;
    wire [62:0] _1438;
    wire [63:0] _1446;
    wire [62:0] _1447;
    wire [63:0] _1455;
    wire [62:0] _1456;
    wire [63:0] _1464;
    wire [62:0] _1465;
    wire [63:0] _1473;
    wire [62:0] _1474;
    wire [63:0] _1482;
    wire [62:0] _1483;
    wire [63:0] _1491;
    wire [62:0] _1492;
    wire [63:0] _1500;
    wire [62:0] _1501;
    wire [63:0] _1509;
    wire [62:0] _1510;
    wire [63:0] _1518;
    wire [62:0] _1519;
    wire [63:0] _1527;
    wire [62:0] _1528;
    wire [63:0] _1536;
    wire [62:0] _1537;
    wire [63:0] _1545;
    wire [62:0] _1546;
    wire [63:0] _1554;
    wire [62:0] _1555;
    wire [63:0] _1563;
    wire [62:0] _1564;
    wire [63:0] _1572;
    wire [62:0] _1573;
    wire [63:0] _1581;
    wire [62:0] _1582;
    wire [63:0] _1590;
    wire [62:0] _1591;
    wire [63:0] _1599;
    wire [62:0] _1600;
    wire [63:0] _1608;
    wire [62:0] _1609;
    wire [63:0] _1617;
    wire [62:0] _1618;
    wire [63:0] _1626;
    wire [62:0] _1627;
    wire [63:0] _1635;
    wire [62:0] _1636;
    wire [63:0] _1644;
    wire [62:0] _1645;
    wire [63:0] _1653;
    wire [62:0] _1654;
    wire [63:0] _1662;
    wire [62:0] _1663;
    wire [63:0] _1671;
    wire [62:0] _1672;
    wire [63:0] _1680;
    wire [62:0] _1681;
    wire [63:0] _1689;
    wire [62:0] _1690;
    wire [63:0] _1698;
    wire [62:0] _1699;
    wire [63:0] _1707;
    wire [62:0] _1708;
    wire [63:0] _1716;
    wire [62:0] _1717;
    wire [63:0] _1725;
    wire [62:0] _1726;
    wire [63:0] _1734;
    wire [62:0] _1735;
    wire [63:0] _1743;
    wire [62:0] _1744;
    wire [63:0] _1752;
    wire [127:0] _1753;
    wire [63:0] _1754;
    wire _1165;
    wire [63:0] _1162;
    wire [63:0] _1163;
    wire [62:0] _1164;
    wire [63:0] _1166;
    wire _1167;
    wire _1168;
    wire _1156;
    wire [63:0] _1153;
    wire [63:0] _1154;
    wire [62:0] _1155;
    wire [63:0] _1157;
    wire _1158;
    wire _1159;
    wire _1147;
    wire [63:0] _1144;
    wire [63:0] _1145;
    wire [62:0] _1146;
    wire [63:0] _1148;
    wire _1149;
    wire _1150;
    wire _1138;
    wire [63:0] _1135;
    wire [63:0] _1136;
    wire [62:0] _1137;
    wire [63:0] _1139;
    wire _1140;
    wire _1141;
    wire _1129;
    wire [63:0] _1126;
    wire [63:0] _1127;
    wire [62:0] _1128;
    wire [63:0] _1130;
    wire _1131;
    wire _1132;
    wire _1120;
    wire [63:0] _1117;
    wire [63:0] _1118;
    wire [62:0] _1119;
    wire [63:0] _1121;
    wire _1122;
    wire _1123;
    wire _1111;
    wire [63:0] _1108;
    wire [63:0] _1109;
    wire [62:0] _1110;
    wire [63:0] _1112;
    wire _1113;
    wire _1114;
    wire _1102;
    wire [63:0] _1099;
    wire [63:0] _1100;
    wire [62:0] _1101;
    wire [63:0] _1103;
    wire _1104;
    wire _1105;
    wire _1093;
    wire [63:0] _1090;
    wire [63:0] _1091;
    wire [62:0] _1092;
    wire [63:0] _1094;
    wire _1095;
    wire _1096;
    wire _1084;
    wire [63:0] _1081;
    wire [63:0] _1082;
    wire [62:0] _1083;
    wire [63:0] _1085;
    wire _1086;
    wire _1087;
    wire _1075;
    wire [63:0] _1072;
    wire [63:0] _1073;
    wire [62:0] _1074;
    wire [63:0] _1076;
    wire _1077;
    wire _1078;
    wire _1066;
    wire [63:0] _1063;
    wire [63:0] _1064;
    wire [62:0] _1065;
    wire [63:0] _1067;
    wire _1068;
    wire _1069;
    wire _1057;
    wire [63:0] _1054;
    wire [63:0] _1055;
    wire [62:0] _1056;
    wire [63:0] _1058;
    wire _1059;
    wire _1060;
    wire _1048;
    wire [63:0] _1045;
    wire [63:0] _1046;
    wire [62:0] _1047;
    wire [63:0] _1049;
    wire _1050;
    wire _1051;
    wire _1039;
    wire [63:0] _1036;
    wire [63:0] _1037;
    wire [62:0] _1038;
    wire [63:0] _1040;
    wire _1041;
    wire _1042;
    wire _1030;
    wire [63:0] _1027;
    wire [63:0] _1028;
    wire [62:0] _1029;
    wire [63:0] _1031;
    wire _1032;
    wire _1033;
    wire _1021;
    wire [63:0] _1018;
    wire [63:0] _1019;
    wire [62:0] _1020;
    wire [63:0] _1022;
    wire _1023;
    wire _1024;
    wire _1012;
    wire [63:0] _1009;
    wire [63:0] _1010;
    wire [62:0] _1011;
    wire [63:0] _1013;
    wire _1014;
    wire _1015;
    wire _1003;
    wire [63:0] _1000;
    wire [63:0] _1001;
    wire [62:0] _1002;
    wire [63:0] _1004;
    wire _1005;
    wire _1006;
    wire _994;
    wire [63:0] _991;
    wire [63:0] _992;
    wire [62:0] _993;
    wire [63:0] _995;
    wire _996;
    wire _997;
    wire _985;
    wire [63:0] _982;
    wire [63:0] _983;
    wire [62:0] _984;
    wire [63:0] _986;
    wire _987;
    wire _988;
    wire _976;
    wire [63:0] _973;
    wire [63:0] _974;
    wire [62:0] _975;
    wire [63:0] _977;
    wire _978;
    wire _979;
    wire _967;
    wire [63:0] _964;
    wire [63:0] _965;
    wire [62:0] _966;
    wire [63:0] _968;
    wire _969;
    wire _970;
    wire _958;
    wire [63:0] _955;
    wire [63:0] _956;
    wire [62:0] _957;
    wire [63:0] _959;
    wire _960;
    wire _961;
    wire _949;
    wire [63:0] _946;
    wire [63:0] _947;
    wire [62:0] _948;
    wire [63:0] _950;
    wire _951;
    wire _952;
    wire _940;
    wire [63:0] _937;
    wire [63:0] _938;
    wire [62:0] _939;
    wire [63:0] _941;
    wire _942;
    wire _943;
    wire _931;
    wire [63:0] _928;
    wire [63:0] _929;
    wire [62:0] _930;
    wire [63:0] _932;
    wire _933;
    wire _934;
    wire _922;
    wire [63:0] _919;
    wire [63:0] _920;
    wire [62:0] _921;
    wire [63:0] _923;
    wire _924;
    wire _925;
    wire _913;
    wire [63:0] _910;
    wire [63:0] _911;
    wire [62:0] _912;
    wire [63:0] _914;
    wire _915;
    wire _916;
    wire _904;
    wire [63:0] _901;
    wire [63:0] _902;
    wire [62:0] _903;
    wire [63:0] _905;
    wire _906;
    wire _907;
    wire _895;
    wire [63:0] _892;
    wire [63:0] _893;
    wire [62:0] _894;
    wire [63:0] _896;
    wire _897;
    wire _898;
    wire _886;
    wire [63:0] _883;
    wire [63:0] _884;
    wire [62:0] _885;
    wire [63:0] _887;
    wire _888;
    wire _889;
    wire _877;
    wire [63:0] _874;
    wire [63:0] _875;
    wire [62:0] _876;
    wire [63:0] _878;
    wire _879;
    wire _880;
    wire _868;
    wire [63:0] _865;
    wire [63:0] _866;
    wire [62:0] _867;
    wire [63:0] _869;
    wire _870;
    wire _871;
    wire _859;
    wire [63:0] _856;
    wire [63:0] _857;
    wire [62:0] _858;
    wire [63:0] _860;
    wire _861;
    wire _862;
    wire _850;
    wire [63:0] _847;
    wire [63:0] _848;
    wire [62:0] _849;
    wire [63:0] _851;
    wire _852;
    wire _853;
    wire _841;
    wire [63:0] _838;
    wire [63:0] _839;
    wire [62:0] _840;
    wire [63:0] _842;
    wire _843;
    wire _844;
    wire _832;
    wire [63:0] _829;
    wire [63:0] _830;
    wire [62:0] _831;
    wire [63:0] _833;
    wire _834;
    wire _835;
    wire _823;
    wire [63:0] _820;
    wire [63:0] _821;
    wire [62:0] _822;
    wire [63:0] _824;
    wire _825;
    wire _826;
    wire _814;
    wire [63:0] _811;
    wire [63:0] _812;
    wire [62:0] _813;
    wire [63:0] _815;
    wire _816;
    wire _817;
    wire _805;
    wire [63:0] _802;
    wire [63:0] _803;
    wire [62:0] _804;
    wire [63:0] _806;
    wire _807;
    wire _808;
    wire _796;
    wire [63:0] _793;
    wire [63:0] _794;
    wire [62:0] _795;
    wire [63:0] _797;
    wire _798;
    wire _799;
    wire _787;
    wire [63:0] _784;
    wire [63:0] _785;
    wire [62:0] _786;
    wire [63:0] _788;
    wire _789;
    wire _790;
    wire _778;
    wire [63:0] _775;
    wire [63:0] _776;
    wire [62:0] _777;
    wire [63:0] _779;
    wire _780;
    wire _781;
    wire _769;
    wire [63:0] _766;
    wire [63:0] _767;
    wire [62:0] _768;
    wire [63:0] _770;
    wire _771;
    wire _772;
    wire _760;
    wire [63:0] _757;
    wire [63:0] _758;
    wire [62:0] _759;
    wire [63:0] _761;
    wire _762;
    wire _763;
    wire _751;
    wire [63:0] _748;
    wire [63:0] _749;
    wire [62:0] _750;
    wire [63:0] _752;
    wire _753;
    wire _754;
    wire _742;
    wire [63:0] _739;
    wire [63:0] _740;
    wire [62:0] _741;
    wire [63:0] _743;
    wire _744;
    wire _745;
    wire _733;
    wire [63:0] _730;
    wire [63:0] _731;
    wire [62:0] _732;
    wire [63:0] _734;
    wire _735;
    wire _736;
    wire _724;
    wire [63:0] _721;
    wire [63:0] _722;
    wire [62:0] _723;
    wire [63:0] _725;
    wire _726;
    wire _727;
    wire _715;
    wire [63:0] _712;
    wire [63:0] _713;
    wire [62:0] _714;
    wire [63:0] _716;
    wire _717;
    wire _718;
    wire _706;
    wire [63:0] _703;
    wire [63:0] _704;
    wire [62:0] _705;
    wire [63:0] _707;
    wire _708;
    wire _709;
    wire _697;
    wire [63:0] _694;
    wire [63:0] _695;
    wire [62:0] _696;
    wire [63:0] _698;
    wire _699;
    wire _700;
    wire _688;
    wire [63:0] _685;
    wire [63:0] _686;
    wire [62:0] _687;
    wire [63:0] _689;
    wire _690;
    wire _691;
    wire _679;
    wire [63:0] _676;
    wire [63:0] _677;
    wire [62:0] _678;
    wire [63:0] _680;
    wire _681;
    wire _682;
    wire _670;
    wire [63:0] _667;
    wire [63:0] _668;
    wire [62:0] _669;
    wire [63:0] _671;
    wire _672;
    wire _673;
    wire _661;
    wire [63:0] _658;
    wire [63:0] _659;
    wire [62:0] _660;
    wire [63:0] _662;
    wire _663;
    wire _664;
    wire _652;
    wire [63:0] _649;
    wire [63:0] _650;
    wire [62:0] _651;
    wire [63:0] _653;
    wire _654;
    wire _655;
    wire _643;
    wire [63:0] _640;
    wire [63:0] _641;
    wire [62:0] _642;
    wire [63:0] _644;
    wire _645;
    wire _646;
    wire _634;
    wire [63:0] _631;
    wire [63:0] _632;
    wire [62:0] _633;
    wire [63:0] _635;
    wire _636;
    wire _637;
    wire _625;
    wire [63:0] _622;
    wire [63:0] _623;
    wire [62:0] _624;
    wire [63:0] _626;
    wire _627;
    wire _628;
    wire _616;
    wire [63:0] _613;
    wire [63:0] _614;
    wire [62:0] _615;
    wire [63:0] _617;
    wire _618;
    wire _619;
    wire _607;
    wire [63:0] _604;
    wire [63:0] _605;
    wire [62:0] _606;
    wire [63:0] _608;
    wire _609;
    wire _610;
    wire [63:0] _597;
    wire _598;
    wire [63:0] _599;
    wire _600;
    wire _601;
    wire [63:0] _602;
    wire [62:0] _603;
    wire [63:0] _611;
    wire [62:0] _612;
    wire [63:0] _620;
    wire [62:0] _621;
    wire [63:0] _629;
    wire [62:0] _630;
    wire [63:0] _638;
    wire [62:0] _639;
    wire [63:0] _647;
    wire [62:0] _648;
    wire [63:0] _656;
    wire [62:0] _657;
    wire [63:0] _665;
    wire [62:0] _666;
    wire [63:0] _674;
    wire [62:0] _675;
    wire [63:0] _683;
    wire [62:0] _684;
    wire [63:0] _692;
    wire [62:0] _693;
    wire [63:0] _701;
    wire [62:0] _702;
    wire [63:0] _710;
    wire [62:0] _711;
    wire [63:0] _719;
    wire [62:0] _720;
    wire [63:0] _728;
    wire [62:0] _729;
    wire [63:0] _737;
    wire [62:0] _738;
    wire [63:0] _746;
    wire [62:0] _747;
    wire [63:0] _755;
    wire [62:0] _756;
    wire [63:0] _764;
    wire [62:0] _765;
    wire [63:0] _773;
    wire [62:0] _774;
    wire [63:0] _782;
    wire [62:0] _783;
    wire [63:0] _791;
    wire [62:0] _792;
    wire [63:0] _800;
    wire [62:0] _801;
    wire [63:0] _809;
    wire [62:0] _810;
    wire [63:0] _818;
    wire [62:0] _819;
    wire [63:0] _827;
    wire [62:0] _828;
    wire [63:0] _836;
    wire [62:0] _837;
    wire [63:0] _845;
    wire [62:0] _846;
    wire [63:0] _854;
    wire [62:0] _855;
    wire [63:0] _863;
    wire [62:0] _864;
    wire [63:0] _872;
    wire [62:0] _873;
    wire [63:0] _881;
    wire [62:0] _882;
    wire [63:0] _890;
    wire [62:0] _891;
    wire [63:0] _899;
    wire [62:0] _900;
    wire [63:0] _908;
    wire [62:0] _909;
    wire [63:0] _917;
    wire [62:0] _918;
    wire [63:0] _926;
    wire [62:0] _927;
    wire [63:0] _935;
    wire [62:0] _936;
    wire [63:0] _944;
    wire [62:0] _945;
    wire [63:0] _953;
    wire [62:0] _954;
    wire [63:0] _962;
    wire [62:0] _963;
    wire [63:0] _971;
    wire [62:0] _972;
    wire [63:0] _980;
    wire [62:0] _981;
    wire [63:0] _989;
    wire [62:0] _990;
    wire [63:0] _998;
    wire [62:0] _999;
    wire [63:0] _1007;
    wire [62:0] _1008;
    wire [63:0] _1016;
    wire [62:0] _1017;
    wire [63:0] _1025;
    wire [62:0] _1026;
    wire [63:0] _1034;
    wire [62:0] _1035;
    wire [63:0] _1043;
    wire [62:0] _1044;
    wire [63:0] _1052;
    wire [62:0] _1053;
    wire [63:0] _1061;
    wire [62:0] _1062;
    wire [63:0] _1070;
    wire [62:0] _1071;
    wire [63:0] _1079;
    wire [62:0] _1080;
    wire [63:0] _1088;
    wire [62:0] _1089;
    wire [63:0] _1097;
    wire [62:0] _1098;
    wire [63:0] _1106;
    wire [62:0] _1107;
    wire [63:0] _1115;
    wire [62:0] _1116;
    wire [63:0] _1124;
    wire [62:0] _1125;
    wire [63:0] _1133;
    wire [62:0] _1134;
    wire [63:0] _1142;
    wire [62:0] _1143;
    wire [63:0] _1151;
    wire [62:0] _1152;
    wire [63:0] _1160;
    wire [62:0] _1161;
    wire [63:0] _1169;
    wire [63:0] _1171;
    wire [127:0] _1172;
    wire [63:0] _1173;
    wire [63:0] _1755;
    wire _583;
    wire [63:0] _580;
    wire [63:0] _581;
    wire [62:0] _582;
    wire [63:0] _584;
    wire _585;
    wire _586;
    wire _574;
    wire [63:0] _571;
    wire [63:0] _572;
    wire [62:0] _573;
    wire [63:0] _575;
    wire _576;
    wire _577;
    wire _565;
    wire [63:0] _562;
    wire [63:0] _563;
    wire [62:0] _564;
    wire [63:0] _566;
    wire _567;
    wire _568;
    wire _556;
    wire [63:0] _553;
    wire [63:0] _554;
    wire [62:0] _555;
    wire [63:0] _557;
    wire _558;
    wire _559;
    wire _547;
    wire [63:0] _544;
    wire [63:0] _545;
    wire [62:0] _546;
    wire [63:0] _548;
    wire _549;
    wire _550;
    wire _538;
    wire [63:0] _535;
    wire [63:0] _536;
    wire [62:0] _537;
    wire [63:0] _539;
    wire _540;
    wire _541;
    wire _529;
    wire [63:0] _526;
    wire [63:0] _527;
    wire [62:0] _528;
    wire [63:0] _530;
    wire _531;
    wire _532;
    wire _520;
    wire [63:0] _517;
    wire [63:0] _518;
    wire [62:0] _519;
    wire [63:0] _521;
    wire _522;
    wire _523;
    wire _511;
    wire [63:0] _508;
    wire [63:0] _509;
    wire [62:0] _510;
    wire [63:0] _512;
    wire _513;
    wire _514;
    wire _502;
    wire [63:0] _499;
    wire [63:0] _500;
    wire [62:0] _501;
    wire [63:0] _503;
    wire _504;
    wire _505;
    wire _493;
    wire [63:0] _490;
    wire [63:0] _491;
    wire [62:0] _492;
    wire [63:0] _494;
    wire _495;
    wire _496;
    wire _484;
    wire [63:0] _481;
    wire [63:0] _482;
    wire [62:0] _483;
    wire [63:0] _485;
    wire _486;
    wire _487;
    wire _475;
    wire [63:0] _472;
    wire [63:0] _473;
    wire [62:0] _474;
    wire [63:0] _476;
    wire _477;
    wire _478;
    wire _466;
    wire [63:0] _463;
    wire [63:0] _464;
    wire [62:0] _465;
    wire [63:0] _467;
    wire _468;
    wire _469;
    wire _457;
    wire [63:0] _454;
    wire [63:0] _455;
    wire [62:0] _456;
    wire [63:0] _458;
    wire _459;
    wire _460;
    wire _448;
    wire [63:0] _445;
    wire [63:0] _446;
    wire [62:0] _447;
    wire [63:0] _449;
    wire _450;
    wire _451;
    wire _439;
    wire [63:0] _436;
    wire [63:0] _437;
    wire [62:0] _438;
    wire [63:0] _440;
    wire _441;
    wire _442;
    wire _430;
    wire [63:0] _427;
    wire [63:0] _428;
    wire [62:0] _429;
    wire [63:0] _431;
    wire _432;
    wire _433;
    wire _421;
    wire [63:0] _418;
    wire [63:0] _419;
    wire [62:0] _420;
    wire [63:0] _422;
    wire _423;
    wire _424;
    wire _412;
    wire [63:0] _409;
    wire [63:0] _410;
    wire [62:0] _411;
    wire [63:0] _413;
    wire _414;
    wire _415;
    wire _403;
    wire [63:0] _400;
    wire [63:0] _401;
    wire [62:0] _402;
    wire [63:0] _404;
    wire _405;
    wire _406;
    wire _394;
    wire [63:0] _391;
    wire [63:0] _392;
    wire [62:0] _393;
    wire [63:0] _395;
    wire _396;
    wire _397;
    wire _385;
    wire [63:0] _382;
    wire [63:0] _383;
    wire [62:0] _384;
    wire [63:0] _386;
    wire _387;
    wire _388;
    wire _376;
    wire [63:0] _373;
    wire [63:0] _374;
    wire [62:0] _375;
    wire [63:0] _377;
    wire _378;
    wire _379;
    wire _367;
    wire [63:0] _364;
    wire [63:0] _365;
    wire [62:0] _366;
    wire [63:0] _368;
    wire _369;
    wire _370;
    wire _358;
    wire [63:0] _355;
    wire [63:0] _356;
    wire [62:0] _357;
    wire [63:0] _359;
    wire _360;
    wire _361;
    wire _349;
    wire [63:0] _346;
    wire [63:0] _347;
    wire [62:0] _348;
    wire [63:0] _350;
    wire _351;
    wire _352;
    wire _340;
    wire [63:0] _337;
    wire [63:0] _338;
    wire [62:0] _339;
    wire [63:0] _341;
    wire _342;
    wire _343;
    wire _331;
    wire [63:0] _328;
    wire [63:0] _329;
    wire [62:0] _330;
    wire [63:0] _332;
    wire _333;
    wire _334;
    wire _322;
    wire [63:0] _319;
    wire [63:0] _320;
    wire [62:0] _321;
    wire [63:0] _323;
    wire _324;
    wire _325;
    wire _313;
    wire [63:0] _310;
    wire [63:0] _311;
    wire [62:0] _312;
    wire [63:0] _314;
    wire _315;
    wire _316;
    wire _304;
    wire [63:0] _301;
    wire [63:0] _302;
    wire [62:0] _303;
    wire [63:0] _305;
    wire _306;
    wire _307;
    wire _295;
    wire [63:0] _292;
    wire [63:0] _293;
    wire [62:0] _294;
    wire [63:0] _296;
    wire _297;
    wire _298;
    wire _286;
    wire [63:0] _283;
    wire [63:0] _284;
    wire [62:0] _285;
    wire [63:0] _287;
    wire _288;
    wire _289;
    wire _277;
    wire [63:0] _274;
    wire [63:0] _275;
    wire [62:0] _276;
    wire [63:0] _278;
    wire _279;
    wire _280;
    wire _268;
    wire [63:0] _265;
    wire [63:0] _266;
    wire [62:0] _267;
    wire [63:0] _269;
    wire _270;
    wire _271;
    wire _259;
    wire [63:0] _256;
    wire [63:0] _257;
    wire [62:0] _258;
    wire [63:0] _260;
    wire _261;
    wire _262;
    wire _250;
    wire [63:0] _247;
    wire [63:0] _248;
    wire [62:0] _249;
    wire [63:0] _251;
    wire _252;
    wire _253;
    wire _241;
    wire [63:0] _238;
    wire [63:0] _239;
    wire [62:0] _240;
    wire [63:0] _242;
    wire _243;
    wire _244;
    wire _232;
    wire [63:0] _229;
    wire [63:0] _230;
    wire [62:0] _231;
    wire [63:0] _233;
    wire _234;
    wire _235;
    wire _223;
    wire [63:0] _220;
    wire [63:0] _221;
    wire [62:0] _222;
    wire [63:0] _224;
    wire _225;
    wire _226;
    wire _214;
    wire [63:0] _211;
    wire [63:0] _212;
    wire [62:0] _213;
    wire [63:0] _215;
    wire _216;
    wire _217;
    wire _205;
    wire [63:0] _202;
    wire [63:0] _203;
    wire [62:0] _204;
    wire [63:0] _206;
    wire _207;
    wire _208;
    wire _196;
    wire [63:0] _193;
    wire [63:0] _194;
    wire [62:0] _195;
    wire [63:0] _197;
    wire _198;
    wire _199;
    wire _187;
    wire [63:0] _184;
    wire [63:0] _185;
    wire [62:0] _186;
    wire [63:0] _188;
    wire _189;
    wire _190;
    wire _178;
    wire [63:0] _175;
    wire [63:0] _176;
    wire [62:0] _177;
    wire [63:0] _179;
    wire _180;
    wire _181;
    wire _169;
    wire [63:0] _166;
    wire [63:0] _167;
    wire [62:0] _168;
    wire [63:0] _170;
    wire _171;
    wire _172;
    wire _160;
    wire [63:0] _157;
    wire [63:0] _158;
    wire [62:0] _159;
    wire [63:0] _161;
    wire _162;
    wire _163;
    wire _151;
    wire [63:0] _148;
    wire [63:0] _149;
    wire [62:0] _150;
    wire [63:0] _152;
    wire _153;
    wire _154;
    wire _142;
    wire [63:0] _139;
    wire [63:0] _140;
    wire [62:0] _141;
    wire [63:0] _143;
    wire _144;
    wire _145;
    wire _133;
    wire [63:0] _130;
    wire [63:0] _131;
    wire [62:0] _132;
    wire [63:0] _134;
    wire _135;
    wire _136;
    wire _124;
    wire [63:0] _121;
    wire [63:0] _122;
    wire [62:0] _123;
    wire [63:0] _125;
    wire _126;
    wire _127;
    wire _115;
    wire [63:0] _112;
    wire [63:0] _113;
    wire [62:0] _114;
    wire [63:0] _116;
    wire _117;
    wire _118;
    wire _106;
    wire [63:0] _103;
    wire [63:0] _104;
    wire [62:0] _105;
    wire [63:0] _107;
    wire _108;
    wire _109;
    wire _97;
    wire [63:0] _94;
    wire [63:0] _95;
    wire [62:0] _96;
    wire [63:0] _98;
    wire _99;
    wire _100;
    wire _88;
    wire [63:0] _85;
    wire [63:0] _86;
    wire [62:0] _87;
    wire [63:0] _89;
    wire _90;
    wire _91;
    wire _79;
    wire [63:0] _76;
    wire [63:0] _77;
    wire [62:0] _78;
    wire [63:0] _80;
    wire _81;
    wire _82;
    wire _70;
    wire [63:0] _67;
    wire [63:0] _68;
    wire [62:0] _69;
    wire [63:0] _71;
    wire _72;
    wire _73;
    wire _61;
    wire [63:0] _58;
    wire [63:0] _59;
    wire [62:0] _60;
    wire [63:0] _62;
    wire _63;
    wire _64;
    wire _52;
    wire [63:0] _49;
    wire [63:0] _50;
    wire [62:0] _51;
    wire [63:0] _53;
    wire _54;
    wire _55;
    wire _43;
    wire [63:0] _40;
    wire [63:0] _41;
    wire [62:0] _42;
    wire [63:0] _44;
    wire _45;
    wire _46;
    wire _34;
    wire [63:0] _31;
    wire [63:0] _32;
    wire [62:0] _33;
    wire [63:0] _35;
    wire _36;
    wire _37;
    wire _25;
    wire [63:0] _22;
    wire [63:0] _23;
    wire [62:0] _24;
    wire [63:0] _26;
    wire _27;
    wire _28;
    wire [63:0] _17;
    wire [63:0] _13;
    wire [63:0] _3;
    wire [63:0] _14;
    wire _15;
    wire [63:0] _16;
    wire _18;
    wire _19;
    wire [63:0] _20;
    wire [62:0] _21;
    wire [63:0] _29;
    wire [62:0] _30;
    wire [63:0] _38;
    wire [62:0] _39;
    wire [63:0] _47;
    wire [62:0] _48;
    wire [63:0] _56;
    wire [62:0] _57;
    wire [63:0] _65;
    wire [62:0] _66;
    wire [63:0] _74;
    wire [62:0] _75;
    wire [63:0] _83;
    wire [62:0] _84;
    wire [63:0] _92;
    wire [62:0] _93;
    wire [63:0] _101;
    wire [62:0] _102;
    wire [63:0] _110;
    wire [62:0] _111;
    wire [63:0] _119;
    wire [62:0] _120;
    wire [63:0] _128;
    wire [62:0] _129;
    wire [63:0] _137;
    wire [62:0] _138;
    wire [63:0] _146;
    wire [62:0] _147;
    wire [63:0] _155;
    wire [62:0] _156;
    wire [63:0] _164;
    wire [62:0] _165;
    wire [63:0] _173;
    wire [62:0] _174;
    wire [63:0] _182;
    wire [62:0] _183;
    wire [63:0] _191;
    wire [62:0] _192;
    wire [63:0] _200;
    wire [62:0] _201;
    wire [63:0] _209;
    wire [62:0] _210;
    wire [63:0] _218;
    wire [62:0] _219;
    wire [63:0] _227;
    wire [62:0] _228;
    wire [63:0] _236;
    wire [62:0] _237;
    wire [63:0] _245;
    wire [62:0] _246;
    wire [63:0] _254;
    wire [62:0] _255;
    wire [63:0] _263;
    wire [62:0] _264;
    wire [63:0] _272;
    wire [62:0] _273;
    wire [63:0] _281;
    wire [62:0] _282;
    wire [63:0] _290;
    wire [62:0] _291;
    wire [63:0] _299;
    wire [62:0] _300;
    wire [63:0] _308;
    wire [62:0] _309;
    wire [63:0] _317;
    wire [62:0] _318;
    wire [63:0] _326;
    wire [62:0] _327;
    wire [63:0] _335;
    wire [62:0] _336;
    wire [63:0] _344;
    wire [62:0] _345;
    wire [63:0] _353;
    wire [62:0] _354;
    wire [63:0] _362;
    wire [62:0] _363;
    wire [63:0] _371;
    wire [62:0] _372;
    wire [63:0] _380;
    wire [62:0] _381;
    wire [63:0] _389;
    wire [62:0] _390;
    wire [63:0] _398;
    wire [62:0] _399;
    wire [63:0] _407;
    wire [62:0] _408;
    wire [63:0] _416;
    wire [62:0] _417;
    wire [63:0] _425;
    wire [62:0] _426;
    wire [63:0] _434;
    wire [62:0] _435;
    wire [63:0] _443;
    wire [62:0] _444;
    wire [63:0] _452;
    wire [62:0] _453;
    wire [63:0] _461;
    wire [62:0] _462;
    wire [63:0] _470;
    wire [62:0] _471;
    wire [63:0] _479;
    wire [62:0] _480;
    wire [63:0] _488;
    wire [62:0] _489;
    wire [63:0] _497;
    wire [62:0] _498;
    wire [63:0] _506;
    wire [62:0] _507;
    wire [63:0] _515;
    wire [62:0] _516;
    wire [63:0] _524;
    wire [62:0] _525;
    wire [63:0] _533;
    wire [62:0] _534;
    wire [63:0] _542;
    wire [62:0] _543;
    wire [63:0] _551;
    wire [62:0] _552;
    wire [63:0] _560;
    wire [62:0] _561;
    wire [63:0] _569;
    wire [62:0] _570;
    wire [63:0] _578;
    wire [62:0] _579;
    wire [63:0] _587;
    wire [127:0] _588;
    wire [63:0] _589;
    wire _590;
    wire [63:0] _591;
    wire [63:0] _7;
    wire [63:0] _5;
    wire _8;
    wire [63:0] _9;
    wire _592;
    wire _593;
    wire [63:0] _1756;
    wire [63:0] _3507;
    wire [63:0] _5258;
    wire [63:0] _7009;
    wire [63:0] _8760;
    assign _22758 = _22189[0:0];
    assign _22755 = _22750 - _22192;
    assign _22756 = _22752 ? _22755 : _22750;
    assign _22757 = _22756[62:0];
    assign _22759 = { _22757,
                      _22758 };
    assign _22760 = _22759 < _22192;
    assign _22761 = ~ _22760;
    assign _22749 = _22189[1:1];
    assign _22746 = _22741 - _22192;
    assign _22747 = _22743 ? _22746 : _22741;
    assign _22748 = _22747[62:0];
    assign _22750 = { _22748,
                      _22749 };
    assign _22751 = _22750 < _22192;
    assign _22752 = ~ _22751;
    assign _22740 = _22189[2:2];
    assign _22737 = _22732 - _22192;
    assign _22738 = _22734 ? _22737 : _22732;
    assign _22739 = _22738[62:0];
    assign _22741 = { _22739,
                      _22740 };
    assign _22742 = _22741 < _22192;
    assign _22743 = ~ _22742;
    assign _22731 = _22189[3:3];
    assign _22728 = _22723 - _22192;
    assign _22729 = _22725 ? _22728 : _22723;
    assign _22730 = _22729[62:0];
    assign _22732 = { _22730,
                      _22731 };
    assign _22733 = _22732 < _22192;
    assign _22734 = ~ _22733;
    assign _22722 = _22189[4:4];
    assign _22719 = _22714 - _22192;
    assign _22720 = _22716 ? _22719 : _22714;
    assign _22721 = _22720[62:0];
    assign _22723 = { _22721,
                      _22722 };
    assign _22724 = _22723 < _22192;
    assign _22725 = ~ _22724;
    assign _22713 = _22189[5:5];
    assign _22710 = _22705 - _22192;
    assign _22711 = _22707 ? _22710 : _22705;
    assign _22712 = _22711[62:0];
    assign _22714 = { _22712,
                      _22713 };
    assign _22715 = _22714 < _22192;
    assign _22716 = ~ _22715;
    assign _22704 = _22189[6:6];
    assign _22701 = _22696 - _22192;
    assign _22702 = _22698 ? _22701 : _22696;
    assign _22703 = _22702[62:0];
    assign _22705 = { _22703,
                      _22704 };
    assign _22706 = _22705 < _22192;
    assign _22707 = ~ _22706;
    assign _22695 = _22189[7:7];
    assign _22692 = _22687 - _22192;
    assign _22693 = _22689 ? _22692 : _22687;
    assign _22694 = _22693[62:0];
    assign _22696 = { _22694,
                      _22695 };
    assign _22697 = _22696 < _22192;
    assign _22698 = ~ _22697;
    assign _22686 = _22189[8:8];
    assign _22683 = _22678 - _22192;
    assign _22684 = _22680 ? _22683 : _22678;
    assign _22685 = _22684[62:0];
    assign _22687 = { _22685,
                      _22686 };
    assign _22688 = _22687 < _22192;
    assign _22689 = ~ _22688;
    assign _22677 = _22189[9:9];
    assign _22674 = _22669 - _22192;
    assign _22675 = _22671 ? _22674 : _22669;
    assign _22676 = _22675[62:0];
    assign _22678 = { _22676,
                      _22677 };
    assign _22679 = _22678 < _22192;
    assign _22680 = ~ _22679;
    assign _22668 = _22189[10:10];
    assign _22665 = _22660 - _22192;
    assign _22666 = _22662 ? _22665 : _22660;
    assign _22667 = _22666[62:0];
    assign _22669 = { _22667,
                      _22668 };
    assign _22670 = _22669 < _22192;
    assign _22671 = ~ _22670;
    assign _22659 = _22189[11:11];
    assign _22656 = _22651 - _22192;
    assign _22657 = _22653 ? _22656 : _22651;
    assign _22658 = _22657[62:0];
    assign _22660 = { _22658,
                      _22659 };
    assign _22661 = _22660 < _22192;
    assign _22662 = ~ _22661;
    assign _22650 = _22189[12:12];
    assign _22647 = _22642 - _22192;
    assign _22648 = _22644 ? _22647 : _22642;
    assign _22649 = _22648[62:0];
    assign _22651 = { _22649,
                      _22650 };
    assign _22652 = _22651 < _22192;
    assign _22653 = ~ _22652;
    assign _22641 = _22189[13:13];
    assign _22638 = _22633 - _22192;
    assign _22639 = _22635 ? _22638 : _22633;
    assign _22640 = _22639[62:0];
    assign _22642 = { _22640,
                      _22641 };
    assign _22643 = _22642 < _22192;
    assign _22644 = ~ _22643;
    assign _22632 = _22189[14:14];
    assign _22629 = _22624 - _22192;
    assign _22630 = _22626 ? _22629 : _22624;
    assign _22631 = _22630[62:0];
    assign _22633 = { _22631,
                      _22632 };
    assign _22634 = _22633 < _22192;
    assign _22635 = ~ _22634;
    assign _22623 = _22189[15:15];
    assign _22620 = _22615 - _22192;
    assign _22621 = _22617 ? _22620 : _22615;
    assign _22622 = _22621[62:0];
    assign _22624 = { _22622,
                      _22623 };
    assign _22625 = _22624 < _22192;
    assign _22626 = ~ _22625;
    assign _22614 = _22189[16:16];
    assign _22611 = _22606 - _22192;
    assign _22612 = _22608 ? _22611 : _22606;
    assign _22613 = _22612[62:0];
    assign _22615 = { _22613,
                      _22614 };
    assign _22616 = _22615 < _22192;
    assign _22617 = ~ _22616;
    assign _22605 = _22189[17:17];
    assign _22602 = _22597 - _22192;
    assign _22603 = _22599 ? _22602 : _22597;
    assign _22604 = _22603[62:0];
    assign _22606 = { _22604,
                      _22605 };
    assign _22607 = _22606 < _22192;
    assign _22608 = ~ _22607;
    assign _22596 = _22189[18:18];
    assign _22593 = _22588 - _22192;
    assign _22594 = _22590 ? _22593 : _22588;
    assign _22595 = _22594[62:0];
    assign _22597 = { _22595,
                      _22596 };
    assign _22598 = _22597 < _22192;
    assign _22599 = ~ _22598;
    assign _22587 = _22189[19:19];
    assign _22584 = _22579 - _22192;
    assign _22585 = _22581 ? _22584 : _22579;
    assign _22586 = _22585[62:0];
    assign _22588 = { _22586,
                      _22587 };
    assign _22589 = _22588 < _22192;
    assign _22590 = ~ _22589;
    assign _22578 = _22189[20:20];
    assign _22575 = _22570 - _22192;
    assign _22576 = _22572 ? _22575 : _22570;
    assign _22577 = _22576[62:0];
    assign _22579 = { _22577,
                      _22578 };
    assign _22580 = _22579 < _22192;
    assign _22581 = ~ _22580;
    assign _22569 = _22189[21:21];
    assign _22566 = _22561 - _22192;
    assign _22567 = _22563 ? _22566 : _22561;
    assign _22568 = _22567[62:0];
    assign _22570 = { _22568,
                      _22569 };
    assign _22571 = _22570 < _22192;
    assign _22572 = ~ _22571;
    assign _22560 = _22189[22:22];
    assign _22557 = _22552 - _22192;
    assign _22558 = _22554 ? _22557 : _22552;
    assign _22559 = _22558[62:0];
    assign _22561 = { _22559,
                      _22560 };
    assign _22562 = _22561 < _22192;
    assign _22563 = ~ _22562;
    assign _22551 = _22189[23:23];
    assign _22548 = _22543 - _22192;
    assign _22549 = _22545 ? _22548 : _22543;
    assign _22550 = _22549[62:0];
    assign _22552 = { _22550,
                      _22551 };
    assign _22553 = _22552 < _22192;
    assign _22554 = ~ _22553;
    assign _22542 = _22189[24:24];
    assign _22539 = _22534 - _22192;
    assign _22540 = _22536 ? _22539 : _22534;
    assign _22541 = _22540[62:0];
    assign _22543 = { _22541,
                      _22542 };
    assign _22544 = _22543 < _22192;
    assign _22545 = ~ _22544;
    assign _22533 = _22189[25:25];
    assign _22530 = _22525 - _22192;
    assign _22531 = _22527 ? _22530 : _22525;
    assign _22532 = _22531[62:0];
    assign _22534 = { _22532,
                      _22533 };
    assign _22535 = _22534 < _22192;
    assign _22536 = ~ _22535;
    assign _22524 = _22189[26:26];
    assign _22521 = _22516 - _22192;
    assign _22522 = _22518 ? _22521 : _22516;
    assign _22523 = _22522[62:0];
    assign _22525 = { _22523,
                      _22524 };
    assign _22526 = _22525 < _22192;
    assign _22527 = ~ _22526;
    assign _22515 = _22189[27:27];
    assign _22512 = _22507 - _22192;
    assign _22513 = _22509 ? _22512 : _22507;
    assign _22514 = _22513[62:0];
    assign _22516 = { _22514,
                      _22515 };
    assign _22517 = _22516 < _22192;
    assign _22518 = ~ _22517;
    assign _22506 = _22189[28:28];
    assign _22503 = _22498 - _22192;
    assign _22504 = _22500 ? _22503 : _22498;
    assign _22505 = _22504[62:0];
    assign _22507 = { _22505,
                      _22506 };
    assign _22508 = _22507 < _22192;
    assign _22509 = ~ _22508;
    assign _22497 = _22189[29:29];
    assign _22494 = _22489 - _22192;
    assign _22495 = _22491 ? _22494 : _22489;
    assign _22496 = _22495[62:0];
    assign _22498 = { _22496,
                      _22497 };
    assign _22499 = _22498 < _22192;
    assign _22500 = ~ _22499;
    assign _22488 = _22189[30:30];
    assign _22485 = _22480 - _22192;
    assign _22486 = _22482 ? _22485 : _22480;
    assign _22487 = _22486[62:0];
    assign _22489 = { _22487,
                      _22488 };
    assign _22490 = _22489 < _22192;
    assign _22491 = ~ _22490;
    assign _22479 = _22189[31:31];
    assign _22476 = _22471 - _22192;
    assign _22477 = _22473 ? _22476 : _22471;
    assign _22478 = _22477[62:0];
    assign _22480 = { _22478,
                      _22479 };
    assign _22481 = _22480 < _22192;
    assign _22482 = ~ _22481;
    assign _22470 = _22189[32:32];
    assign _22467 = _22462 - _22192;
    assign _22468 = _22464 ? _22467 : _22462;
    assign _22469 = _22468[62:0];
    assign _22471 = { _22469,
                      _22470 };
    assign _22472 = _22471 < _22192;
    assign _22473 = ~ _22472;
    assign _22461 = _22189[33:33];
    assign _22458 = _22453 - _22192;
    assign _22459 = _22455 ? _22458 : _22453;
    assign _22460 = _22459[62:0];
    assign _22462 = { _22460,
                      _22461 };
    assign _22463 = _22462 < _22192;
    assign _22464 = ~ _22463;
    assign _22452 = _22189[34:34];
    assign _22449 = _22444 - _22192;
    assign _22450 = _22446 ? _22449 : _22444;
    assign _22451 = _22450[62:0];
    assign _22453 = { _22451,
                      _22452 };
    assign _22454 = _22453 < _22192;
    assign _22455 = ~ _22454;
    assign _22443 = _22189[35:35];
    assign _22440 = _22435 - _22192;
    assign _22441 = _22437 ? _22440 : _22435;
    assign _22442 = _22441[62:0];
    assign _22444 = { _22442,
                      _22443 };
    assign _22445 = _22444 < _22192;
    assign _22446 = ~ _22445;
    assign _22434 = _22189[36:36];
    assign _22431 = _22426 - _22192;
    assign _22432 = _22428 ? _22431 : _22426;
    assign _22433 = _22432[62:0];
    assign _22435 = { _22433,
                      _22434 };
    assign _22436 = _22435 < _22192;
    assign _22437 = ~ _22436;
    assign _22425 = _22189[37:37];
    assign _22422 = _22417 - _22192;
    assign _22423 = _22419 ? _22422 : _22417;
    assign _22424 = _22423[62:0];
    assign _22426 = { _22424,
                      _22425 };
    assign _22427 = _22426 < _22192;
    assign _22428 = ~ _22427;
    assign _22416 = _22189[38:38];
    assign _22413 = _22408 - _22192;
    assign _22414 = _22410 ? _22413 : _22408;
    assign _22415 = _22414[62:0];
    assign _22417 = { _22415,
                      _22416 };
    assign _22418 = _22417 < _22192;
    assign _22419 = ~ _22418;
    assign _22407 = _22189[39:39];
    assign _22404 = _22399 - _22192;
    assign _22405 = _22401 ? _22404 : _22399;
    assign _22406 = _22405[62:0];
    assign _22408 = { _22406,
                      _22407 };
    assign _22409 = _22408 < _22192;
    assign _22410 = ~ _22409;
    assign _22398 = _22189[40:40];
    assign _22395 = _22390 - _22192;
    assign _22396 = _22392 ? _22395 : _22390;
    assign _22397 = _22396[62:0];
    assign _22399 = { _22397,
                      _22398 };
    assign _22400 = _22399 < _22192;
    assign _22401 = ~ _22400;
    assign _22389 = _22189[41:41];
    assign _22386 = _22381 - _22192;
    assign _22387 = _22383 ? _22386 : _22381;
    assign _22388 = _22387[62:0];
    assign _22390 = { _22388,
                      _22389 };
    assign _22391 = _22390 < _22192;
    assign _22392 = ~ _22391;
    assign _22380 = _22189[42:42];
    assign _22377 = _22372 - _22192;
    assign _22378 = _22374 ? _22377 : _22372;
    assign _22379 = _22378[62:0];
    assign _22381 = { _22379,
                      _22380 };
    assign _22382 = _22381 < _22192;
    assign _22383 = ~ _22382;
    assign _22371 = _22189[43:43];
    assign _22368 = _22363 - _22192;
    assign _22369 = _22365 ? _22368 : _22363;
    assign _22370 = _22369[62:0];
    assign _22372 = { _22370,
                      _22371 };
    assign _22373 = _22372 < _22192;
    assign _22374 = ~ _22373;
    assign _22362 = _22189[44:44];
    assign _22359 = _22354 - _22192;
    assign _22360 = _22356 ? _22359 : _22354;
    assign _22361 = _22360[62:0];
    assign _22363 = { _22361,
                      _22362 };
    assign _22364 = _22363 < _22192;
    assign _22365 = ~ _22364;
    assign _22353 = _22189[45:45];
    assign _22350 = _22345 - _22192;
    assign _22351 = _22347 ? _22350 : _22345;
    assign _22352 = _22351[62:0];
    assign _22354 = { _22352,
                      _22353 };
    assign _22355 = _22354 < _22192;
    assign _22356 = ~ _22355;
    assign _22344 = _22189[46:46];
    assign _22341 = _22336 - _22192;
    assign _22342 = _22338 ? _22341 : _22336;
    assign _22343 = _22342[62:0];
    assign _22345 = { _22343,
                      _22344 };
    assign _22346 = _22345 < _22192;
    assign _22347 = ~ _22346;
    assign _22335 = _22189[47:47];
    assign _22332 = _22327 - _22192;
    assign _22333 = _22329 ? _22332 : _22327;
    assign _22334 = _22333[62:0];
    assign _22336 = { _22334,
                      _22335 };
    assign _22337 = _22336 < _22192;
    assign _22338 = ~ _22337;
    assign _22326 = _22189[48:48];
    assign _22323 = _22318 - _22192;
    assign _22324 = _22320 ? _22323 : _22318;
    assign _22325 = _22324[62:0];
    assign _22327 = { _22325,
                      _22326 };
    assign _22328 = _22327 < _22192;
    assign _22329 = ~ _22328;
    assign _22317 = _22189[49:49];
    assign _22314 = _22309 - _22192;
    assign _22315 = _22311 ? _22314 : _22309;
    assign _22316 = _22315[62:0];
    assign _22318 = { _22316,
                      _22317 };
    assign _22319 = _22318 < _22192;
    assign _22320 = ~ _22319;
    assign _22308 = _22189[50:50];
    assign _22305 = _22300 - _22192;
    assign _22306 = _22302 ? _22305 : _22300;
    assign _22307 = _22306[62:0];
    assign _22309 = { _22307,
                      _22308 };
    assign _22310 = _22309 < _22192;
    assign _22311 = ~ _22310;
    assign _22299 = _22189[51:51];
    assign _22296 = _22291 - _22192;
    assign _22297 = _22293 ? _22296 : _22291;
    assign _22298 = _22297[62:0];
    assign _22300 = { _22298,
                      _22299 };
    assign _22301 = _22300 < _22192;
    assign _22302 = ~ _22301;
    assign _22290 = _22189[52:52];
    assign _22287 = _22282 - _22192;
    assign _22288 = _22284 ? _22287 : _22282;
    assign _22289 = _22288[62:0];
    assign _22291 = { _22289,
                      _22290 };
    assign _22292 = _22291 < _22192;
    assign _22293 = ~ _22292;
    assign _22281 = _22189[53:53];
    assign _22278 = _22273 - _22192;
    assign _22279 = _22275 ? _22278 : _22273;
    assign _22280 = _22279[62:0];
    assign _22282 = { _22280,
                      _22281 };
    assign _22283 = _22282 < _22192;
    assign _22284 = ~ _22283;
    assign _22272 = _22189[54:54];
    assign _22269 = _22264 - _22192;
    assign _22270 = _22266 ? _22269 : _22264;
    assign _22271 = _22270[62:0];
    assign _22273 = { _22271,
                      _22272 };
    assign _22274 = _22273 < _22192;
    assign _22275 = ~ _22274;
    assign _22263 = _22189[55:55];
    assign _22260 = _22255 - _22192;
    assign _22261 = _22257 ? _22260 : _22255;
    assign _22262 = _22261[62:0];
    assign _22264 = { _22262,
                      _22263 };
    assign _22265 = _22264 < _22192;
    assign _22266 = ~ _22265;
    assign _22254 = _22189[56:56];
    assign _22251 = _22246 - _22192;
    assign _22252 = _22248 ? _22251 : _22246;
    assign _22253 = _22252[62:0];
    assign _22255 = { _22253,
                      _22254 };
    assign _22256 = _22255 < _22192;
    assign _22257 = ~ _22256;
    assign _22245 = _22189[57:57];
    assign _22242 = _22237 - _22192;
    assign _22243 = _22239 ? _22242 : _22237;
    assign _22244 = _22243[62:0];
    assign _22246 = { _22244,
                      _22245 };
    assign _22247 = _22246 < _22192;
    assign _22248 = ~ _22247;
    assign _22236 = _22189[58:58];
    assign _22233 = _22228 - _22192;
    assign _22234 = _22230 ? _22233 : _22228;
    assign _22235 = _22234[62:0];
    assign _22237 = { _22235,
                      _22236 };
    assign _22238 = _22237 < _22192;
    assign _22239 = ~ _22238;
    assign _22227 = _22189[59:59];
    assign _22224 = _22219 - _22192;
    assign _22225 = _22221 ? _22224 : _22219;
    assign _22226 = _22225[62:0];
    assign _22228 = { _22226,
                      _22227 };
    assign _22229 = _22228 < _22192;
    assign _22230 = ~ _22229;
    assign _22218 = _22189[60:60];
    assign _22215 = _22210 - _22192;
    assign _22216 = _22212 ? _22215 : _22210;
    assign _22217 = _22216[62:0];
    assign _22219 = { _22217,
                      _22218 };
    assign _22220 = _22219 < _22192;
    assign _22221 = ~ _22220;
    assign _22209 = _22189[61:61];
    assign _22206 = _22201 - _22192;
    assign _22207 = _22203 ? _22206 : _22201;
    assign _22208 = _22207[62:0];
    assign _22210 = { _22208,
                      _22209 };
    assign _22211 = _22210 < _22192;
    assign _22212 = ~ _22211;
    assign _22200 = _22189[62:62];
    assign _22197 = _22191 - _22192;
    assign _22198 = _22194 ? _22197 : _22191;
    assign _22199 = _22198[62:0];
    assign _22201 = { _22199,
                      _22200 };
    assign _22202 = _22201 < _22192;
    assign _22203 = ~ _22202;
    assign _22192 = 64'b0000000000000000000000000000000000000000000000000000000000000010;
    assign _22186 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    assign _22187 = _22179 + _22186;
    assign _22188 = _22179 * _22187;
    assign _22189 = _22188[63:0];
    assign _22190 = _22189[63:63];
    assign _22185 = 63'b000000000000000000000000000000000000000000000000000000000000000;
    assign _22191 = { _22185,
                      _22190 };
    assign _22193 = _22191 < _22192;
    assign _22194 = ~ _22193;
    assign _22195 = { _22185,
                      _22194 };
    assign _22196 = _22195[62:0];
    assign _22204 = { _22196,
                      _22203 };
    assign _22205 = _22204[62:0];
    assign _22213 = { _22205,
                      _22212 };
    assign _22214 = _22213[62:0];
    assign _22222 = { _22214,
                      _22221 };
    assign _22223 = _22222[62:0];
    assign _22231 = { _22223,
                      _22230 };
    assign _22232 = _22231[62:0];
    assign _22240 = { _22232,
                      _22239 };
    assign _22241 = _22240[62:0];
    assign _22249 = { _22241,
                      _22248 };
    assign _22250 = _22249[62:0];
    assign _22258 = { _22250,
                      _22257 };
    assign _22259 = _22258[62:0];
    assign _22267 = { _22259,
                      _22266 };
    assign _22268 = _22267[62:0];
    assign _22276 = { _22268,
                      _22275 };
    assign _22277 = _22276[62:0];
    assign _22285 = { _22277,
                      _22284 };
    assign _22286 = _22285[62:0];
    assign _22294 = { _22286,
                      _22293 };
    assign _22295 = _22294[62:0];
    assign _22303 = { _22295,
                      _22302 };
    assign _22304 = _22303[62:0];
    assign _22312 = { _22304,
                      _22311 };
    assign _22313 = _22312[62:0];
    assign _22321 = { _22313,
                      _22320 };
    assign _22322 = _22321[62:0];
    assign _22330 = { _22322,
                      _22329 };
    assign _22331 = _22330[62:0];
    assign _22339 = { _22331,
                      _22338 };
    assign _22340 = _22339[62:0];
    assign _22348 = { _22340,
                      _22347 };
    assign _22349 = _22348[62:0];
    assign _22357 = { _22349,
                      _22356 };
    assign _22358 = _22357[62:0];
    assign _22366 = { _22358,
                      _22365 };
    assign _22367 = _22366[62:0];
    assign _22375 = { _22367,
                      _22374 };
    assign _22376 = _22375[62:0];
    assign _22384 = { _22376,
                      _22383 };
    assign _22385 = _22384[62:0];
    assign _22393 = { _22385,
                      _22392 };
    assign _22394 = _22393[62:0];
    assign _22402 = { _22394,
                      _22401 };
    assign _22403 = _22402[62:0];
    assign _22411 = { _22403,
                      _22410 };
    assign _22412 = _22411[62:0];
    assign _22420 = { _22412,
                      _22419 };
    assign _22421 = _22420[62:0];
    assign _22429 = { _22421,
                      _22428 };
    assign _22430 = _22429[62:0];
    assign _22438 = { _22430,
                      _22437 };
    assign _22439 = _22438[62:0];
    assign _22447 = { _22439,
                      _22446 };
    assign _22448 = _22447[62:0];
    assign _22456 = { _22448,
                      _22455 };
    assign _22457 = _22456[62:0];
    assign _22465 = { _22457,
                      _22464 };
    assign _22466 = _22465[62:0];
    assign _22474 = { _22466,
                      _22473 };
    assign _22475 = _22474[62:0];
    assign _22483 = { _22475,
                      _22482 };
    assign _22484 = _22483[62:0];
    assign _22492 = { _22484,
                      _22491 };
    assign _22493 = _22492[62:0];
    assign _22501 = { _22493,
                      _22500 };
    assign _22502 = _22501[62:0];
    assign _22510 = { _22502,
                      _22509 };
    assign _22511 = _22510[62:0];
    assign _22519 = { _22511,
                      _22518 };
    assign _22520 = _22519[62:0];
    assign _22528 = { _22520,
                      _22527 };
    assign _22529 = _22528[62:0];
    assign _22537 = { _22529,
                      _22536 };
    assign _22538 = _22537[62:0];
    assign _22546 = { _22538,
                      _22545 };
    assign _22547 = _22546[62:0];
    assign _22555 = { _22547,
                      _22554 };
    assign _22556 = _22555[62:0];
    assign _22564 = { _22556,
                      _22563 };
    assign _22565 = _22564[62:0];
    assign _22573 = { _22565,
                      _22572 };
    assign _22574 = _22573[62:0];
    assign _22582 = { _22574,
                      _22581 };
    assign _22583 = _22582[62:0];
    assign _22591 = { _22583,
                      _22590 };
    assign _22592 = _22591[62:0];
    assign _22600 = { _22592,
                      _22599 };
    assign _22601 = _22600[62:0];
    assign _22609 = { _22601,
                      _22608 };
    assign _22610 = _22609[62:0];
    assign _22618 = { _22610,
                      _22617 };
    assign _22619 = _22618[62:0];
    assign _22627 = { _22619,
                      _22626 };
    assign _22628 = _22627[62:0];
    assign _22636 = { _22628,
                      _22635 };
    assign _22637 = _22636[62:0];
    assign _22645 = { _22637,
                      _22644 };
    assign _22646 = _22645[62:0];
    assign _22654 = { _22646,
                      _22653 };
    assign _22655 = _22654[62:0];
    assign _22663 = { _22655,
                      _22662 };
    assign _22664 = _22663[62:0];
    assign _22672 = { _22664,
                      _22671 };
    assign _22673 = _22672[62:0];
    assign _22681 = { _22673,
                      _22680 };
    assign _22682 = _22681[62:0];
    assign _22690 = { _22682,
                      _22689 };
    assign _22691 = _22690[62:0];
    assign _22699 = { _22691,
                      _22698 };
    assign _22700 = _22699[62:0];
    assign _22708 = { _22700,
                      _22707 };
    assign _22709 = _22708[62:0];
    assign _22717 = { _22709,
                      _22716 };
    assign _22718 = _22717[62:0];
    assign _22726 = { _22718,
                      _22725 };
    assign _22727 = _22726[62:0];
    assign _22735 = { _22727,
                      _22734 };
    assign _22736 = _22735[62:0];
    assign _22744 = { _22736,
                      _22743 };
    assign _22745 = _22744[62:0];
    assign _22753 = { _22745,
                      _22752 };
    assign _22754 = _22753[62:0];
    assign _22762 = { _22754,
                      _22761 };
    assign _22763 = _21027 * _22762;
    assign _22764 = _22763[63:0];
    assign _22175 = _21607[0:0];
    assign _22172 = _22167 - _21027;
    assign _22173 = _22169 ? _22172 : _22167;
    assign _22174 = _22173[62:0];
    assign _22176 = { _22174,
                      _22175 };
    assign _22177 = _22176 < _21027;
    assign _22178 = ~ _22177;
    assign _22166 = _21607[1:1];
    assign _22163 = _22158 - _21027;
    assign _22164 = _22160 ? _22163 : _22158;
    assign _22165 = _22164[62:0];
    assign _22167 = { _22165,
                      _22166 };
    assign _22168 = _22167 < _21027;
    assign _22169 = ~ _22168;
    assign _22157 = _21607[2:2];
    assign _22154 = _22149 - _21027;
    assign _22155 = _22151 ? _22154 : _22149;
    assign _22156 = _22155[62:0];
    assign _22158 = { _22156,
                      _22157 };
    assign _22159 = _22158 < _21027;
    assign _22160 = ~ _22159;
    assign _22148 = _21607[3:3];
    assign _22145 = _22140 - _21027;
    assign _22146 = _22142 ? _22145 : _22140;
    assign _22147 = _22146[62:0];
    assign _22149 = { _22147,
                      _22148 };
    assign _22150 = _22149 < _21027;
    assign _22151 = ~ _22150;
    assign _22139 = _21607[4:4];
    assign _22136 = _22131 - _21027;
    assign _22137 = _22133 ? _22136 : _22131;
    assign _22138 = _22137[62:0];
    assign _22140 = { _22138,
                      _22139 };
    assign _22141 = _22140 < _21027;
    assign _22142 = ~ _22141;
    assign _22130 = _21607[5:5];
    assign _22127 = _22122 - _21027;
    assign _22128 = _22124 ? _22127 : _22122;
    assign _22129 = _22128[62:0];
    assign _22131 = { _22129,
                      _22130 };
    assign _22132 = _22131 < _21027;
    assign _22133 = ~ _22132;
    assign _22121 = _21607[6:6];
    assign _22118 = _22113 - _21027;
    assign _22119 = _22115 ? _22118 : _22113;
    assign _22120 = _22119[62:0];
    assign _22122 = { _22120,
                      _22121 };
    assign _22123 = _22122 < _21027;
    assign _22124 = ~ _22123;
    assign _22112 = _21607[7:7];
    assign _22109 = _22104 - _21027;
    assign _22110 = _22106 ? _22109 : _22104;
    assign _22111 = _22110[62:0];
    assign _22113 = { _22111,
                      _22112 };
    assign _22114 = _22113 < _21027;
    assign _22115 = ~ _22114;
    assign _22103 = _21607[8:8];
    assign _22100 = _22095 - _21027;
    assign _22101 = _22097 ? _22100 : _22095;
    assign _22102 = _22101[62:0];
    assign _22104 = { _22102,
                      _22103 };
    assign _22105 = _22104 < _21027;
    assign _22106 = ~ _22105;
    assign _22094 = _21607[9:9];
    assign _22091 = _22086 - _21027;
    assign _22092 = _22088 ? _22091 : _22086;
    assign _22093 = _22092[62:0];
    assign _22095 = { _22093,
                      _22094 };
    assign _22096 = _22095 < _21027;
    assign _22097 = ~ _22096;
    assign _22085 = _21607[10:10];
    assign _22082 = _22077 - _21027;
    assign _22083 = _22079 ? _22082 : _22077;
    assign _22084 = _22083[62:0];
    assign _22086 = { _22084,
                      _22085 };
    assign _22087 = _22086 < _21027;
    assign _22088 = ~ _22087;
    assign _22076 = _21607[11:11];
    assign _22073 = _22068 - _21027;
    assign _22074 = _22070 ? _22073 : _22068;
    assign _22075 = _22074[62:0];
    assign _22077 = { _22075,
                      _22076 };
    assign _22078 = _22077 < _21027;
    assign _22079 = ~ _22078;
    assign _22067 = _21607[12:12];
    assign _22064 = _22059 - _21027;
    assign _22065 = _22061 ? _22064 : _22059;
    assign _22066 = _22065[62:0];
    assign _22068 = { _22066,
                      _22067 };
    assign _22069 = _22068 < _21027;
    assign _22070 = ~ _22069;
    assign _22058 = _21607[13:13];
    assign _22055 = _22050 - _21027;
    assign _22056 = _22052 ? _22055 : _22050;
    assign _22057 = _22056[62:0];
    assign _22059 = { _22057,
                      _22058 };
    assign _22060 = _22059 < _21027;
    assign _22061 = ~ _22060;
    assign _22049 = _21607[14:14];
    assign _22046 = _22041 - _21027;
    assign _22047 = _22043 ? _22046 : _22041;
    assign _22048 = _22047[62:0];
    assign _22050 = { _22048,
                      _22049 };
    assign _22051 = _22050 < _21027;
    assign _22052 = ~ _22051;
    assign _22040 = _21607[15:15];
    assign _22037 = _22032 - _21027;
    assign _22038 = _22034 ? _22037 : _22032;
    assign _22039 = _22038[62:0];
    assign _22041 = { _22039,
                      _22040 };
    assign _22042 = _22041 < _21027;
    assign _22043 = ~ _22042;
    assign _22031 = _21607[16:16];
    assign _22028 = _22023 - _21027;
    assign _22029 = _22025 ? _22028 : _22023;
    assign _22030 = _22029[62:0];
    assign _22032 = { _22030,
                      _22031 };
    assign _22033 = _22032 < _21027;
    assign _22034 = ~ _22033;
    assign _22022 = _21607[17:17];
    assign _22019 = _22014 - _21027;
    assign _22020 = _22016 ? _22019 : _22014;
    assign _22021 = _22020[62:0];
    assign _22023 = { _22021,
                      _22022 };
    assign _22024 = _22023 < _21027;
    assign _22025 = ~ _22024;
    assign _22013 = _21607[18:18];
    assign _22010 = _22005 - _21027;
    assign _22011 = _22007 ? _22010 : _22005;
    assign _22012 = _22011[62:0];
    assign _22014 = { _22012,
                      _22013 };
    assign _22015 = _22014 < _21027;
    assign _22016 = ~ _22015;
    assign _22004 = _21607[19:19];
    assign _22001 = _21996 - _21027;
    assign _22002 = _21998 ? _22001 : _21996;
    assign _22003 = _22002[62:0];
    assign _22005 = { _22003,
                      _22004 };
    assign _22006 = _22005 < _21027;
    assign _22007 = ~ _22006;
    assign _21995 = _21607[20:20];
    assign _21992 = _21987 - _21027;
    assign _21993 = _21989 ? _21992 : _21987;
    assign _21994 = _21993[62:0];
    assign _21996 = { _21994,
                      _21995 };
    assign _21997 = _21996 < _21027;
    assign _21998 = ~ _21997;
    assign _21986 = _21607[21:21];
    assign _21983 = _21978 - _21027;
    assign _21984 = _21980 ? _21983 : _21978;
    assign _21985 = _21984[62:0];
    assign _21987 = { _21985,
                      _21986 };
    assign _21988 = _21987 < _21027;
    assign _21989 = ~ _21988;
    assign _21977 = _21607[22:22];
    assign _21974 = _21969 - _21027;
    assign _21975 = _21971 ? _21974 : _21969;
    assign _21976 = _21975[62:0];
    assign _21978 = { _21976,
                      _21977 };
    assign _21979 = _21978 < _21027;
    assign _21980 = ~ _21979;
    assign _21968 = _21607[23:23];
    assign _21965 = _21960 - _21027;
    assign _21966 = _21962 ? _21965 : _21960;
    assign _21967 = _21966[62:0];
    assign _21969 = { _21967,
                      _21968 };
    assign _21970 = _21969 < _21027;
    assign _21971 = ~ _21970;
    assign _21959 = _21607[24:24];
    assign _21956 = _21951 - _21027;
    assign _21957 = _21953 ? _21956 : _21951;
    assign _21958 = _21957[62:0];
    assign _21960 = { _21958,
                      _21959 };
    assign _21961 = _21960 < _21027;
    assign _21962 = ~ _21961;
    assign _21950 = _21607[25:25];
    assign _21947 = _21942 - _21027;
    assign _21948 = _21944 ? _21947 : _21942;
    assign _21949 = _21948[62:0];
    assign _21951 = { _21949,
                      _21950 };
    assign _21952 = _21951 < _21027;
    assign _21953 = ~ _21952;
    assign _21941 = _21607[26:26];
    assign _21938 = _21933 - _21027;
    assign _21939 = _21935 ? _21938 : _21933;
    assign _21940 = _21939[62:0];
    assign _21942 = { _21940,
                      _21941 };
    assign _21943 = _21942 < _21027;
    assign _21944 = ~ _21943;
    assign _21932 = _21607[27:27];
    assign _21929 = _21924 - _21027;
    assign _21930 = _21926 ? _21929 : _21924;
    assign _21931 = _21930[62:0];
    assign _21933 = { _21931,
                      _21932 };
    assign _21934 = _21933 < _21027;
    assign _21935 = ~ _21934;
    assign _21923 = _21607[28:28];
    assign _21920 = _21915 - _21027;
    assign _21921 = _21917 ? _21920 : _21915;
    assign _21922 = _21921[62:0];
    assign _21924 = { _21922,
                      _21923 };
    assign _21925 = _21924 < _21027;
    assign _21926 = ~ _21925;
    assign _21914 = _21607[29:29];
    assign _21911 = _21906 - _21027;
    assign _21912 = _21908 ? _21911 : _21906;
    assign _21913 = _21912[62:0];
    assign _21915 = { _21913,
                      _21914 };
    assign _21916 = _21915 < _21027;
    assign _21917 = ~ _21916;
    assign _21905 = _21607[30:30];
    assign _21902 = _21897 - _21027;
    assign _21903 = _21899 ? _21902 : _21897;
    assign _21904 = _21903[62:0];
    assign _21906 = { _21904,
                      _21905 };
    assign _21907 = _21906 < _21027;
    assign _21908 = ~ _21907;
    assign _21896 = _21607[31:31];
    assign _21893 = _21888 - _21027;
    assign _21894 = _21890 ? _21893 : _21888;
    assign _21895 = _21894[62:0];
    assign _21897 = { _21895,
                      _21896 };
    assign _21898 = _21897 < _21027;
    assign _21899 = ~ _21898;
    assign _21887 = _21607[32:32];
    assign _21884 = _21879 - _21027;
    assign _21885 = _21881 ? _21884 : _21879;
    assign _21886 = _21885[62:0];
    assign _21888 = { _21886,
                      _21887 };
    assign _21889 = _21888 < _21027;
    assign _21890 = ~ _21889;
    assign _21878 = _21607[33:33];
    assign _21875 = _21870 - _21027;
    assign _21876 = _21872 ? _21875 : _21870;
    assign _21877 = _21876[62:0];
    assign _21879 = { _21877,
                      _21878 };
    assign _21880 = _21879 < _21027;
    assign _21881 = ~ _21880;
    assign _21869 = _21607[34:34];
    assign _21866 = _21861 - _21027;
    assign _21867 = _21863 ? _21866 : _21861;
    assign _21868 = _21867[62:0];
    assign _21870 = { _21868,
                      _21869 };
    assign _21871 = _21870 < _21027;
    assign _21872 = ~ _21871;
    assign _21860 = _21607[35:35];
    assign _21857 = _21852 - _21027;
    assign _21858 = _21854 ? _21857 : _21852;
    assign _21859 = _21858[62:0];
    assign _21861 = { _21859,
                      _21860 };
    assign _21862 = _21861 < _21027;
    assign _21863 = ~ _21862;
    assign _21851 = _21607[36:36];
    assign _21848 = _21843 - _21027;
    assign _21849 = _21845 ? _21848 : _21843;
    assign _21850 = _21849[62:0];
    assign _21852 = { _21850,
                      _21851 };
    assign _21853 = _21852 < _21027;
    assign _21854 = ~ _21853;
    assign _21842 = _21607[37:37];
    assign _21839 = _21834 - _21027;
    assign _21840 = _21836 ? _21839 : _21834;
    assign _21841 = _21840[62:0];
    assign _21843 = { _21841,
                      _21842 };
    assign _21844 = _21843 < _21027;
    assign _21845 = ~ _21844;
    assign _21833 = _21607[38:38];
    assign _21830 = _21825 - _21027;
    assign _21831 = _21827 ? _21830 : _21825;
    assign _21832 = _21831[62:0];
    assign _21834 = { _21832,
                      _21833 };
    assign _21835 = _21834 < _21027;
    assign _21836 = ~ _21835;
    assign _21824 = _21607[39:39];
    assign _21821 = _21816 - _21027;
    assign _21822 = _21818 ? _21821 : _21816;
    assign _21823 = _21822[62:0];
    assign _21825 = { _21823,
                      _21824 };
    assign _21826 = _21825 < _21027;
    assign _21827 = ~ _21826;
    assign _21815 = _21607[40:40];
    assign _21812 = _21807 - _21027;
    assign _21813 = _21809 ? _21812 : _21807;
    assign _21814 = _21813[62:0];
    assign _21816 = { _21814,
                      _21815 };
    assign _21817 = _21816 < _21027;
    assign _21818 = ~ _21817;
    assign _21806 = _21607[41:41];
    assign _21803 = _21798 - _21027;
    assign _21804 = _21800 ? _21803 : _21798;
    assign _21805 = _21804[62:0];
    assign _21807 = { _21805,
                      _21806 };
    assign _21808 = _21807 < _21027;
    assign _21809 = ~ _21808;
    assign _21797 = _21607[42:42];
    assign _21794 = _21789 - _21027;
    assign _21795 = _21791 ? _21794 : _21789;
    assign _21796 = _21795[62:0];
    assign _21798 = { _21796,
                      _21797 };
    assign _21799 = _21798 < _21027;
    assign _21800 = ~ _21799;
    assign _21788 = _21607[43:43];
    assign _21785 = _21780 - _21027;
    assign _21786 = _21782 ? _21785 : _21780;
    assign _21787 = _21786[62:0];
    assign _21789 = { _21787,
                      _21788 };
    assign _21790 = _21789 < _21027;
    assign _21791 = ~ _21790;
    assign _21779 = _21607[44:44];
    assign _21776 = _21771 - _21027;
    assign _21777 = _21773 ? _21776 : _21771;
    assign _21778 = _21777[62:0];
    assign _21780 = { _21778,
                      _21779 };
    assign _21781 = _21780 < _21027;
    assign _21782 = ~ _21781;
    assign _21770 = _21607[45:45];
    assign _21767 = _21762 - _21027;
    assign _21768 = _21764 ? _21767 : _21762;
    assign _21769 = _21768[62:0];
    assign _21771 = { _21769,
                      _21770 };
    assign _21772 = _21771 < _21027;
    assign _21773 = ~ _21772;
    assign _21761 = _21607[46:46];
    assign _21758 = _21753 - _21027;
    assign _21759 = _21755 ? _21758 : _21753;
    assign _21760 = _21759[62:0];
    assign _21762 = { _21760,
                      _21761 };
    assign _21763 = _21762 < _21027;
    assign _21764 = ~ _21763;
    assign _21752 = _21607[47:47];
    assign _21749 = _21744 - _21027;
    assign _21750 = _21746 ? _21749 : _21744;
    assign _21751 = _21750[62:0];
    assign _21753 = { _21751,
                      _21752 };
    assign _21754 = _21753 < _21027;
    assign _21755 = ~ _21754;
    assign _21743 = _21607[48:48];
    assign _21740 = _21735 - _21027;
    assign _21741 = _21737 ? _21740 : _21735;
    assign _21742 = _21741[62:0];
    assign _21744 = { _21742,
                      _21743 };
    assign _21745 = _21744 < _21027;
    assign _21746 = ~ _21745;
    assign _21734 = _21607[49:49];
    assign _21731 = _21726 - _21027;
    assign _21732 = _21728 ? _21731 : _21726;
    assign _21733 = _21732[62:0];
    assign _21735 = { _21733,
                      _21734 };
    assign _21736 = _21735 < _21027;
    assign _21737 = ~ _21736;
    assign _21725 = _21607[50:50];
    assign _21722 = _21717 - _21027;
    assign _21723 = _21719 ? _21722 : _21717;
    assign _21724 = _21723[62:0];
    assign _21726 = { _21724,
                      _21725 };
    assign _21727 = _21726 < _21027;
    assign _21728 = ~ _21727;
    assign _21716 = _21607[51:51];
    assign _21713 = _21708 - _21027;
    assign _21714 = _21710 ? _21713 : _21708;
    assign _21715 = _21714[62:0];
    assign _21717 = { _21715,
                      _21716 };
    assign _21718 = _21717 < _21027;
    assign _21719 = ~ _21718;
    assign _21707 = _21607[52:52];
    assign _21704 = _21699 - _21027;
    assign _21705 = _21701 ? _21704 : _21699;
    assign _21706 = _21705[62:0];
    assign _21708 = { _21706,
                      _21707 };
    assign _21709 = _21708 < _21027;
    assign _21710 = ~ _21709;
    assign _21698 = _21607[53:53];
    assign _21695 = _21690 - _21027;
    assign _21696 = _21692 ? _21695 : _21690;
    assign _21697 = _21696[62:0];
    assign _21699 = { _21697,
                      _21698 };
    assign _21700 = _21699 < _21027;
    assign _21701 = ~ _21700;
    assign _21689 = _21607[54:54];
    assign _21686 = _21681 - _21027;
    assign _21687 = _21683 ? _21686 : _21681;
    assign _21688 = _21687[62:0];
    assign _21690 = { _21688,
                      _21689 };
    assign _21691 = _21690 < _21027;
    assign _21692 = ~ _21691;
    assign _21680 = _21607[55:55];
    assign _21677 = _21672 - _21027;
    assign _21678 = _21674 ? _21677 : _21672;
    assign _21679 = _21678[62:0];
    assign _21681 = { _21679,
                      _21680 };
    assign _21682 = _21681 < _21027;
    assign _21683 = ~ _21682;
    assign _21671 = _21607[56:56];
    assign _21668 = _21663 - _21027;
    assign _21669 = _21665 ? _21668 : _21663;
    assign _21670 = _21669[62:0];
    assign _21672 = { _21670,
                      _21671 };
    assign _21673 = _21672 < _21027;
    assign _21674 = ~ _21673;
    assign _21662 = _21607[57:57];
    assign _21659 = _21654 - _21027;
    assign _21660 = _21656 ? _21659 : _21654;
    assign _21661 = _21660[62:0];
    assign _21663 = { _21661,
                      _21662 };
    assign _21664 = _21663 < _21027;
    assign _21665 = ~ _21664;
    assign _21653 = _21607[58:58];
    assign _21650 = _21645 - _21027;
    assign _21651 = _21647 ? _21650 : _21645;
    assign _21652 = _21651[62:0];
    assign _21654 = { _21652,
                      _21653 };
    assign _21655 = _21654 < _21027;
    assign _21656 = ~ _21655;
    assign _21644 = _21607[59:59];
    assign _21641 = _21636 - _21027;
    assign _21642 = _21638 ? _21641 : _21636;
    assign _21643 = _21642[62:0];
    assign _21645 = { _21643,
                      _21644 };
    assign _21646 = _21645 < _21027;
    assign _21647 = ~ _21646;
    assign _21635 = _21607[60:60];
    assign _21632 = _21627 - _21027;
    assign _21633 = _21629 ? _21632 : _21627;
    assign _21634 = _21633[62:0];
    assign _21636 = { _21634,
                      _21635 };
    assign _21637 = _21636 < _21027;
    assign _21638 = ~ _21637;
    assign _21626 = _21607[61:61];
    assign _21623 = _21618 - _21027;
    assign _21624 = _21620 ? _21623 : _21618;
    assign _21625 = _21624[62:0];
    assign _21627 = { _21625,
                      _21626 };
    assign _21628 = _21627 < _21027;
    assign _21629 = ~ _21628;
    assign _21617 = _21607[62:62];
    assign _21614 = _21609 - _21027;
    assign _21615 = _21611 ? _21614 : _21609;
    assign _21616 = _21615[62:0];
    assign _21618 = { _21616,
                      _21617 };
    assign _21619 = _21618 < _21027;
    assign _21620 = ~ _21619;
    assign _21607 = _21019 - _21601;
    assign _21608 = _21607[63:63];
    assign _21609 = { _22185,
                      _21608 };
    assign _21610 = _21609 < _21027;
    assign _21611 = ~ _21610;
    assign _21612 = { _22185,
                      _21611 };
    assign _21613 = _21612[62:0];
    assign _21621 = { _21613,
                      _21620 };
    assign _21622 = _21621[62:0];
    assign _21630 = { _21622,
                      _21629 };
    assign _21631 = _21630[62:0];
    assign _21639 = { _21631,
                      _21638 };
    assign _21640 = _21639[62:0];
    assign _21648 = { _21640,
                      _21647 };
    assign _21649 = _21648[62:0];
    assign _21657 = { _21649,
                      _21656 };
    assign _21658 = _21657[62:0];
    assign _21666 = { _21658,
                      _21665 };
    assign _21667 = _21666[62:0];
    assign _21675 = { _21667,
                      _21674 };
    assign _21676 = _21675[62:0];
    assign _21684 = { _21676,
                      _21683 };
    assign _21685 = _21684[62:0];
    assign _21693 = { _21685,
                      _21692 };
    assign _21694 = _21693[62:0];
    assign _21702 = { _21694,
                      _21701 };
    assign _21703 = _21702[62:0];
    assign _21711 = { _21703,
                      _21710 };
    assign _21712 = _21711[62:0];
    assign _21720 = { _21712,
                      _21719 };
    assign _21721 = _21720[62:0];
    assign _21729 = { _21721,
                      _21728 };
    assign _21730 = _21729[62:0];
    assign _21738 = { _21730,
                      _21737 };
    assign _21739 = _21738[62:0];
    assign _21747 = { _21739,
                      _21746 };
    assign _21748 = _21747[62:0];
    assign _21756 = { _21748,
                      _21755 };
    assign _21757 = _21756[62:0];
    assign _21765 = { _21757,
                      _21764 };
    assign _21766 = _21765[62:0];
    assign _21774 = { _21766,
                      _21773 };
    assign _21775 = _21774[62:0];
    assign _21783 = { _21775,
                      _21782 };
    assign _21784 = _21783[62:0];
    assign _21792 = { _21784,
                      _21791 };
    assign _21793 = _21792[62:0];
    assign _21801 = { _21793,
                      _21800 };
    assign _21802 = _21801[62:0];
    assign _21810 = { _21802,
                      _21809 };
    assign _21811 = _21810[62:0];
    assign _21819 = { _21811,
                      _21818 };
    assign _21820 = _21819[62:0];
    assign _21828 = { _21820,
                      _21827 };
    assign _21829 = _21828[62:0];
    assign _21837 = { _21829,
                      _21836 };
    assign _21838 = _21837[62:0];
    assign _21846 = { _21838,
                      _21845 };
    assign _21847 = _21846[62:0];
    assign _21855 = { _21847,
                      _21854 };
    assign _21856 = _21855[62:0];
    assign _21864 = { _21856,
                      _21863 };
    assign _21865 = _21864[62:0];
    assign _21873 = { _21865,
                      _21872 };
    assign _21874 = _21873[62:0];
    assign _21882 = { _21874,
                      _21881 };
    assign _21883 = _21882[62:0];
    assign _21891 = { _21883,
                      _21890 };
    assign _21892 = _21891[62:0];
    assign _21900 = { _21892,
                      _21899 };
    assign _21901 = _21900[62:0];
    assign _21909 = { _21901,
                      _21908 };
    assign _21910 = _21909[62:0];
    assign _21918 = { _21910,
                      _21917 };
    assign _21919 = _21918[62:0];
    assign _21927 = { _21919,
                      _21926 };
    assign _21928 = _21927[62:0];
    assign _21936 = { _21928,
                      _21935 };
    assign _21937 = _21936[62:0];
    assign _21945 = { _21937,
                      _21944 };
    assign _21946 = _21945[62:0];
    assign _21954 = { _21946,
                      _21953 };
    assign _21955 = _21954[62:0];
    assign _21963 = { _21955,
                      _21962 };
    assign _21964 = _21963[62:0];
    assign _21972 = { _21964,
                      _21971 };
    assign _21973 = _21972[62:0];
    assign _21981 = { _21973,
                      _21980 };
    assign _21982 = _21981[62:0];
    assign _21990 = { _21982,
                      _21989 };
    assign _21991 = _21990[62:0];
    assign _21999 = { _21991,
                      _21998 };
    assign _22000 = _21999[62:0];
    assign _22008 = { _22000,
                      _22007 };
    assign _22009 = _22008[62:0];
    assign _22017 = { _22009,
                      _22016 };
    assign _22018 = _22017[62:0];
    assign _22026 = { _22018,
                      _22025 };
    assign _22027 = _22026[62:0];
    assign _22035 = { _22027,
                      _22034 };
    assign _22036 = _22035[62:0];
    assign _22044 = { _22036,
                      _22043 };
    assign _22045 = _22044[62:0];
    assign _22053 = { _22045,
                      _22052 };
    assign _22054 = _22053[62:0];
    assign _22062 = { _22054,
                      _22061 };
    assign _22063 = _22062[62:0];
    assign _22071 = { _22063,
                      _22070 };
    assign _22072 = _22071[62:0];
    assign _22080 = { _22072,
                      _22079 };
    assign _22081 = _22080[62:0];
    assign _22089 = { _22081,
                      _22088 };
    assign _22090 = _22089[62:0];
    assign _22098 = { _22090,
                      _22097 };
    assign _22099 = _22098[62:0];
    assign _22107 = { _22099,
                      _22106 };
    assign _22108 = _22107[62:0];
    assign _22116 = { _22108,
                      _22115 };
    assign _22117 = _22116[62:0];
    assign _22125 = { _22117,
                      _22124 };
    assign _22126 = _22125[62:0];
    assign _22134 = { _22126,
                      _22133 };
    assign _22135 = _22134[62:0];
    assign _22143 = { _22135,
                      _22142 };
    assign _22144 = _22143[62:0];
    assign _22152 = { _22144,
                      _22151 };
    assign _22153 = _22152[62:0];
    assign _22161 = { _22153,
                      _22160 };
    assign _22162 = _22161[62:0];
    assign _22170 = { _22162,
                      _22169 };
    assign _22171 = _22170[62:0];
    assign _22179 = { _22171,
                      _22178 };
    assign _22181 = _22179 + _22186;
    assign _22182 = _22181 * _21601;
    assign _22183 = _22182[63:0];
    assign _22765 = _22183 + _22764;
    assign _21604 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign _21593 = _21024[0:0];
    assign _21590 = _21585 - _21027;
    assign _21591 = _21587 ? _21590 : _21585;
    assign _21592 = _21591[62:0];
    assign _21594 = { _21592,
                      _21593 };
    assign _21595 = _21594 < _21027;
    assign _21596 = ~ _21595;
    assign _21584 = _21024[1:1];
    assign _21581 = _21576 - _21027;
    assign _21582 = _21578 ? _21581 : _21576;
    assign _21583 = _21582[62:0];
    assign _21585 = { _21583,
                      _21584 };
    assign _21586 = _21585 < _21027;
    assign _21587 = ~ _21586;
    assign _21575 = _21024[2:2];
    assign _21572 = _21567 - _21027;
    assign _21573 = _21569 ? _21572 : _21567;
    assign _21574 = _21573[62:0];
    assign _21576 = { _21574,
                      _21575 };
    assign _21577 = _21576 < _21027;
    assign _21578 = ~ _21577;
    assign _21566 = _21024[3:3];
    assign _21563 = _21558 - _21027;
    assign _21564 = _21560 ? _21563 : _21558;
    assign _21565 = _21564[62:0];
    assign _21567 = { _21565,
                      _21566 };
    assign _21568 = _21567 < _21027;
    assign _21569 = ~ _21568;
    assign _21557 = _21024[4:4];
    assign _21554 = _21549 - _21027;
    assign _21555 = _21551 ? _21554 : _21549;
    assign _21556 = _21555[62:0];
    assign _21558 = { _21556,
                      _21557 };
    assign _21559 = _21558 < _21027;
    assign _21560 = ~ _21559;
    assign _21548 = _21024[5:5];
    assign _21545 = _21540 - _21027;
    assign _21546 = _21542 ? _21545 : _21540;
    assign _21547 = _21546[62:0];
    assign _21549 = { _21547,
                      _21548 };
    assign _21550 = _21549 < _21027;
    assign _21551 = ~ _21550;
    assign _21539 = _21024[6:6];
    assign _21536 = _21531 - _21027;
    assign _21537 = _21533 ? _21536 : _21531;
    assign _21538 = _21537[62:0];
    assign _21540 = { _21538,
                      _21539 };
    assign _21541 = _21540 < _21027;
    assign _21542 = ~ _21541;
    assign _21530 = _21024[7:7];
    assign _21527 = _21522 - _21027;
    assign _21528 = _21524 ? _21527 : _21522;
    assign _21529 = _21528[62:0];
    assign _21531 = { _21529,
                      _21530 };
    assign _21532 = _21531 < _21027;
    assign _21533 = ~ _21532;
    assign _21521 = _21024[8:8];
    assign _21518 = _21513 - _21027;
    assign _21519 = _21515 ? _21518 : _21513;
    assign _21520 = _21519[62:0];
    assign _21522 = { _21520,
                      _21521 };
    assign _21523 = _21522 < _21027;
    assign _21524 = ~ _21523;
    assign _21512 = _21024[9:9];
    assign _21509 = _21504 - _21027;
    assign _21510 = _21506 ? _21509 : _21504;
    assign _21511 = _21510[62:0];
    assign _21513 = { _21511,
                      _21512 };
    assign _21514 = _21513 < _21027;
    assign _21515 = ~ _21514;
    assign _21503 = _21024[10:10];
    assign _21500 = _21495 - _21027;
    assign _21501 = _21497 ? _21500 : _21495;
    assign _21502 = _21501[62:0];
    assign _21504 = { _21502,
                      _21503 };
    assign _21505 = _21504 < _21027;
    assign _21506 = ~ _21505;
    assign _21494 = _21024[11:11];
    assign _21491 = _21486 - _21027;
    assign _21492 = _21488 ? _21491 : _21486;
    assign _21493 = _21492[62:0];
    assign _21495 = { _21493,
                      _21494 };
    assign _21496 = _21495 < _21027;
    assign _21497 = ~ _21496;
    assign _21485 = _21024[12:12];
    assign _21482 = _21477 - _21027;
    assign _21483 = _21479 ? _21482 : _21477;
    assign _21484 = _21483[62:0];
    assign _21486 = { _21484,
                      _21485 };
    assign _21487 = _21486 < _21027;
    assign _21488 = ~ _21487;
    assign _21476 = _21024[13:13];
    assign _21473 = _21468 - _21027;
    assign _21474 = _21470 ? _21473 : _21468;
    assign _21475 = _21474[62:0];
    assign _21477 = { _21475,
                      _21476 };
    assign _21478 = _21477 < _21027;
    assign _21479 = ~ _21478;
    assign _21467 = _21024[14:14];
    assign _21464 = _21459 - _21027;
    assign _21465 = _21461 ? _21464 : _21459;
    assign _21466 = _21465[62:0];
    assign _21468 = { _21466,
                      _21467 };
    assign _21469 = _21468 < _21027;
    assign _21470 = ~ _21469;
    assign _21458 = _21024[15:15];
    assign _21455 = _21450 - _21027;
    assign _21456 = _21452 ? _21455 : _21450;
    assign _21457 = _21456[62:0];
    assign _21459 = { _21457,
                      _21458 };
    assign _21460 = _21459 < _21027;
    assign _21461 = ~ _21460;
    assign _21449 = _21024[16:16];
    assign _21446 = _21441 - _21027;
    assign _21447 = _21443 ? _21446 : _21441;
    assign _21448 = _21447[62:0];
    assign _21450 = { _21448,
                      _21449 };
    assign _21451 = _21450 < _21027;
    assign _21452 = ~ _21451;
    assign _21440 = _21024[17:17];
    assign _21437 = _21432 - _21027;
    assign _21438 = _21434 ? _21437 : _21432;
    assign _21439 = _21438[62:0];
    assign _21441 = { _21439,
                      _21440 };
    assign _21442 = _21441 < _21027;
    assign _21443 = ~ _21442;
    assign _21431 = _21024[18:18];
    assign _21428 = _21423 - _21027;
    assign _21429 = _21425 ? _21428 : _21423;
    assign _21430 = _21429[62:0];
    assign _21432 = { _21430,
                      _21431 };
    assign _21433 = _21432 < _21027;
    assign _21434 = ~ _21433;
    assign _21422 = _21024[19:19];
    assign _21419 = _21414 - _21027;
    assign _21420 = _21416 ? _21419 : _21414;
    assign _21421 = _21420[62:0];
    assign _21423 = { _21421,
                      _21422 };
    assign _21424 = _21423 < _21027;
    assign _21425 = ~ _21424;
    assign _21413 = _21024[20:20];
    assign _21410 = _21405 - _21027;
    assign _21411 = _21407 ? _21410 : _21405;
    assign _21412 = _21411[62:0];
    assign _21414 = { _21412,
                      _21413 };
    assign _21415 = _21414 < _21027;
    assign _21416 = ~ _21415;
    assign _21404 = _21024[21:21];
    assign _21401 = _21396 - _21027;
    assign _21402 = _21398 ? _21401 : _21396;
    assign _21403 = _21402[62:0];
    assign _21405 = { _21403,
                      _21404 };
    assign _21406 = _21405 < _21027;
    assign _21407 = ~ _21406;
    assign _21395 = _21024[22:22];
    assign _21392 = _21387 - _21027;
    assign _21393 = _21389 ? _21392 : _21387;
    assign _21394 = _21393[62:0];
    assign _21396 = { _21394,
                      _21395 };
    assign _21397 = _21396 < _21027;
    assign _21398 = ~ _21397;
    assign _21386 = _21024[23:23];
    assign _21383 = _21378 - _21027;
    assign _21384 = _21380 ? _21383 : _21378;
    assign _21385 = _21384[62:0];
    assign _21387 = { _21385,
                      _21386 };
    assign _21388 = _21387 < _21027;
    assign _21389 = ~ _21388;
    assign _21377 = _21024[24:24];
    assign _21374 = _21369 - _21027;
    assign _21375 = _21371 ? _21374 : _21369;
    assign _21376 = _21375[62:0];
    assign _21378 = { _21376,
                      _21377 };
    assign _21379 = _21378 < _21027;
    assign _21380 = ~ _21379;
    assign _21368 = _21024[25:25];
    assign _21365 = _21360 - _21027;
    assign _21366 = _21362 ? _21365 : _21360;
    assign _21367 = _21366[62:0];
    assign _21369 = { _21367,
                      _21368 };
    assign _21370 = _21369 < _21027;
    assign _21371 = ~ _21370;
    assign _21359 = _21024[26:26];
    assign _21356 = _21351 - _21027;
    assign _21357 = _21353 ? _21356 : _21351;
    assign _21358 = _21357[62:0];
    assign _21360 = { _21358,
                      _21359 };
    assign _21361 = _21360 < _21027;
    assign _21362 = ~ _21361;
    assign _21350 = _21024[27:27];
    assign _21347 = _21342 - _21027;
    assign _21348 = _21344 ? _21347 : _21342;
    assign _21349 = _21348[62:0];
    assign _21351 = { _21349,
                      _21350 };
    assign _21352 = _21351 < _21027;
    assign _21353 = ~ _21352;
    assign _21341 = _21024[28:28];
    assign _21338 = _21333 - _21027;
    assign _21339 = _21335 ? _21338 : _21333;
    assign _21340 = _21339[62:0];
    assign _21342 = { _21340,
                      _21341 };
    assign _21343 = _21342 < _21027;
    assign _21344 = ~ _21343;
    assign _21332 = _21024[29:29];
    assign _21329 = _21324 - _21027;
    assign _21330 = _21326 ? _21329 : _21324;
    assign _21331 = _21330[62:0];
    assign _21333 = { _21331,
                      _21332 };
    assign _21334 = _21333 < _21027;
    assign _21335 = ~ _21334;
    assign _21323 = _21024[30:30];
    assign _21320 = _21315 - _21027;
    assign _21321 = _21317 ? _21320 : _21315;
    assign _21322 = _21321[62:0];
    assign _21324 = { _21322,
                      _21323 };
    assign _21325 = _21324 < _21027;
    assign _21326 = ~ _21325;
    assign _21314 = _21024[31:31];
    assign _21311 = _21306 - _21027;
    assign _21312 = _21308 ? _21311 : _21306;
    assign _21313 = _21312[62:0];
    assign _21315 = { _21313,
                      _21314 };
    assign _21316 = _21315 < _21027;
    assign _21317 = ~ _21316;
    assign _21305 = _21024[32:32];
    assign _21302 = _21297 - _21027;
    assign _21303 = _21299 ? _21302 : _21297;
    assign _21304 = _21303[62:0];
    assign _21306 = { _21304,
                      _21305 };
    assign _21307 = _21306 < _21027;
    assign _21308 = ~ _21307;
    assign _21296 = _21024[33:33];
    assign _21293 = _21288 - _21027;
    assign _21294 = _21290 ? _21293 : _21288;
    assign _21295 = _21294[62:0];
    assign _21297 = { _21295,
                      _21296 };
    assign _21298 = _21297 < _21027;
    assign _21299 = ~ _21298;
    assign _21287 = _21024[34:34];
    assign _21284 = _21279 - _21027;
    assign _21285 = _21281 ? _21284 : _21279;
    assign _21286 = _21285[62:0];
    assign _21288 = { _21286,
                      _21287 };
    assign _21289 = _21288 < _21027;
    assign _21290 = ~ _21289;
    assign _21278 = _21024[35:35];
    assign _21275 = _21270 - _21027;
    assign _21276 = _21272 ? _21275 : _21270;
    assign _21277 = _21276[62:0];
    assign _21279 = { _21277,
                      _21278 };
    assign _21280 = _21279 < _21027;
    assign _21281 = ~ _21280;
    assign _21269 = _21024[36:36];
    assign _21266 = _21261 - _21027;
    assign _21267 = _21263 ? _21266 : _21261;
    assign _21268 = _21267[62:0];
    assign _21270 = { _21268,
                      _21269 };
    assign _21271 = _21270 < _21027;
    assign _21272 = ~ _21271;
    assign _21260 = _21024[37:37];
    assign _21257 = _21252 - _21027;
    assign _21258 = _21254 ? _21257 : _21252;
    assign _21259 = _21258[62:0];
    assign _21261 = { _21259,
                      _21260 };
    assign _21262 = _21261 < _21027;
    assign _21263 = ~ _21262;
    assign _21251 = _21024[38:38];
    assign _21248 = _21243 - _21027;
    assign _21249 = _21245 ? _21248 : _21243;
    assign _21250 = _21249[62:0];
    assign _21252 = { _21250,
                      _21251 };
    assign _21253 = _21252 < _21027;
    assign _21254 = ~ _21253;
    assign _21242 = _21024[39:39];
    assign _21239 = _21234 - _21027;
    assign _21240 = _21236 ? _21239 : _21234;
    assign _21241 = _21240[62:0];
    assign _21243 = { _21241,
                      _21242 };
    assign _21244 = _21243 < _21027;
    assign _21245 = ~ _21244;
    assign _21233 = _21024[40:40];
    assign _21230 = _21225 - _21027;
    assign _21231 = _21227 ? _21230 : _21225;
    assign _21232 = _21231[62:0];
    assign _21234 = { _21232,
                      _21233 };
    assign _21235 = _21234 < _21027;
    assign _21236 = ~ _21235;
    assign _21224 = _21024[41:41];
    assign _21221 = _21216 - _21027;
    assign _21222 = _21218 ? _21221 : _21216;
    assign _21223 = _21222[62:0];
    assign _21225 = { _21223,
                      _21224 };
    assign _21226 = _21225 < _21027;
    assign _21227 = ~ _21226;
    assign _21215 = _21024[42:42];
    assign _21212 = _21207 - _21027;
    assign _21213 = _21209 ? _21212 : _21207;
    assign _21214 = _21213[62:0];
    assign _21216 = { _21214,
                      _21215 };
    assign _21217 = _21216 < _21027;
    assign _21218 = ~ _21217;
    assign _21206 = _21024[43:43];
    assign _21203 = _21198 - _21027;
    assign _21204 = _21200 ? _21203 : _21198;
    assign _21205 = _21204[62:0];
    assign _21207 = { _21205,
                      _21206 };
    assign _21208 = _21207 < _21027;
    assign _21209 = ~ _21208;
    assign _21197 = _21024[44:44];
    assign _21194 = _21189 - _21027;
    assign _21195 = _21191 ? _21194 : _21189;
    assign _21196 = _21195[62:0];
    assign _21198 = { _21196,
                      _21197 };
    assign _21199 = _21198 < _21027;
    assign _21200 = ~ _21199;
    assign _21188 = _21024[45:45];
    assign _21185 = _21180 - _21027;
    assign _21186 = _21182 ? _21185 : _21180;
    assign _21187 = _21186[62:0];
    assign _21189 = { _21187,
                      _21188 };
    assign _21190 = _21189 < _21027;
    assign _21191 = ~ _21190;
    assign _21179 = _21024[46:46];
    assign _21176 = _21171 - _21027;
    assign _21177 = _21173 ? _21176 : _21171;
    assign _21178 = _21177[62:0];
    assign _21180 = { _21178,
                      _21179 };
    assign _21181 = _21180 < _21027;
    assign _21182 = ~ _21181;
    assign _21170 = _21024[47:47];
    assign _21167 = _21162 - _21027;
    assign _21168 = _21164 ? _21167 : _21162;
    assign _21169 = _21168[62:0];
    assign _21171 = { _21169,
                      _21170 };
    assign _21172 = _21171 < _21027;
    assign _21173 = ~ _21172;
    assign _21161 = _21024[48:48];
    assign _21158 = _21153 - _21027;
    assign _21159 = _21155 ? _21158 : _21153;
    assign _21160 = _21159[62:0];
    assign _21162 = { _21160,
                      _21161 };
    assign _21163 = _21162 < _21027;
    assign _21164 = ~ _21163;
    assign _21152 = _21024[49:49];
    assign _21149 = _21144 - _21027;
    assign _21150 = _21146 ? _21149 : _21144;
    assign _21151 = _21150[62:0];
    assign _21153 = { _21151,
                      _21152 };
    assign _21154 = _21153 < _21027;
    assign _21155 = ~ _21154;
    assign _21143 = _21024[50:50];
    assign _21140 = _21135 - _21027;
    assign _21141 = _21137 ? _21140 : _21135;
    assign _21142 = _21141[62:0];
    assign _21144 = { _21142,
                      _21143 };
    assign _21145 = _21144 < _21027;
    assign _21146 = ~ _21145;
    assign _21134 = _21024[51:51];
    assign _21131 = _21126 - _21027;
    assign _21132 = _21128 ? _21131 : _21126;
    assign _21133 = _21132[62:0];
    assign _21135 = { _21133,
                      _21134 };
    assign _21136 = _21135 < _21027;
    assign _21137 = ~ _21136;
    assign _21125 = _21024[52:52];
    assign _21122 = _21117 - _21027;
    assign _21123 = _21119 ? _21122 : _21117;
    assign _21124 = _21123[62:0];
    assign _21126 = { _21124,
                      _21125 };
    assign _21127 = _21126 < _21027;
    assign _21128 = ~ _21127;
    assign _21116 = _21024[53:53];
    assign _21113 = _21108 - _21027;
    assign _21114 = _21110 ? _21113 : _21108;
    assign _21115 = _21114[62:0];
    assign _21117 = { _21115,
                      _21116 };
    assign _21118 = _21117 < _21027;
    assign _21119 = ~ _21118;
    assign _21107 = _21024[54:54];
    assign _21104 = _21099 - _21027;
    assign _21105 = _21101 ? _21104 : _21099;
    assign _21106 = _21105[62:0];
    assign _21108 = { _21106,
                      _21107 };
    assign _21109 = _21108 < _21027;
    assign _21110 = ~ _21109;
    assign _21098 = _21024[55:55];
    assign _21095 = _21090 - _21027;
    assign _21096 = _21092 ? _21095 : _21090;
    assign _21097 = _21096[62:0];
    assign _21099 = { _21097,
                      _21098 };
    assign _21100 = _21099 < _21027;
    assign _21101 = ~ _21100;
    assign _21089 = _21024[56:56];
    assign _21086 = _21081 - _21027;
    assign _21087 = _21083 ? _21086 : _21081;
    assign _21088 = _21087[62:0];
    assign _21090 = { _21088,
                      _21089 };
    assign _21091 = _21090 < _21027;
    assign _21092 = ~ _21091;
    assign _21080 = _21024[57:57];
    assign _21077 = _21072 - _21027;
    assign _21078 = _21074 ? _21077 : _21072;
    assign _21079 = _21078[62:0];
    assign _21081 = { _21079,
                      _21080 };
    assign _21082 = _21081 < _21027;
    assign _21083 = ~ _21082;
    assign _21071 = _21024[58:58];
    assign _21068 = _21063 - _21027;
    assign _21069 = _21065 ? _21068 : _21063;
    assign _21070 = _21069[62:0];
    assign _21072 = { _21070,
                      _21071 };
    assign _21073 = _21072 < _21027;
    assign _21074 = ~ _21073;
    assign _21062 = _21024[59:59];
    assign _21059 = _21054 - _21027;
    assign _21060 = _21056 ? _21059 : _21054;
    assign _21061 = _21060[62:0];
    assign _21063 = { _21061,
                      _21062 };
    assign _21064 = _21063 < _21027;
    assign _21065 = ~ _21064;
    assign _21053 = _21024[60:60];
    assign _21050 = _21045 - _21027;
    assign _21051 = _21047 ? _21050 : _21045;
    assign _21052 = _21051[62:0];
    assign _21054 = { _21052,
                      _21053 };
    assign _21055 = _21054 < _21027;
    assign _21056 = ~ _21055;
    assign _21044 = _21024[61:61];
    assign _21041 = _21036 - _21027;
    assign _21042 = _21038 ? _21041 : _21036;
    assign _21043 = _21042[62:0];
    assign _21045 = { _21043,
                      _21044 };
    assign _21046 = _21045 < _21027;
    assign _21047 = ~ _21046;
    assign _21035 = _21024[62:62];
    assign _21032 = _21026 - _21027;
    assign _21033 = _21029 ? _21032 : _21026;
    assign _21034 = _21033[62:0];
    assign _21036 = { _21034,
                      _21035 };
    assign _21037 = _21036 < _21027;
    assign _21038 = ~ _21037;
    assign _21027 = 64'b0000000000000000000000000000000001000010001110100011010111000111;
    assign _21023 = 64'b0000000000000000000000000000000001000010001110100011010111000110;
    assign _21024 = _3 + _21023;
    assign _21025 = _21024[63:63];
    assign _21026 = { _22185,
                      _21025 };
    assign _21028 = _21026 < _21027;
    assign _21029 = ~ _21028;
    assign _21030 = { _22185,
                      _21029 };
    assign _21031 = _21030[62:0];
    assign _21039 = { _21031,
                      _21038 };
    assign _21040 = _21039[62:0];
    assign _21048 = { _21040,
                      _21047 };
    assign _21049 = _21048[62:0];
    assign _21057 = { _21049,
                      _21056 };
    assign _21058 = _21057[62:0];
    assign _21066 = { _21058,
                      _21065 };
    assign _21067 = _21066[62:0];
    assign _21075 = { _21067,
                      _21074 };
    assign _21076 = _21075[62:0];
    assign _21084 = { _21076,
                      _21083 };
    assign _21085 = _21084[62:0];
    assign _21093 = { _21085,
                      _21092 };
    assign _21094 = _21093[62:0];
    assign _21102 = { _21094,
                      _21101 };
    assign _21103 = _21102[62:0];
    assign _21111 = { _21103,
                      _21110 };
    assign _21112 = _21111[62:0];
    assign _21120 = { _21112,
                      _21119 };
    assign _21121 = _21120[62:0];
    assign _21129 = { _21121,
                      _21128 };
    assign _21130 = _21129[62:0];
    assign _21138 = { _21130,
                      _21137 };
    assign _21139 = _21138[62:0];
    assign _21147 = { _21139,
                      _21146 };
    assign _21148 = _21147[62:0];
    assign _21156 = { _21148,
                      _21155 };
    assign _21157 = _21156[62:0];
    assign _21165 = { _21157,
                      _21164 };
    assign _21166 = _21165[62:0];
    assign _21174 = { _21166,
                      _21173 };
    assign _21175 = _21174[62:0];
    assign _21183 = { _21175,
                      _21182 };
    assign _21184 = _21183[62:0];
    assign _21192 = { _21184,
                      _21191 };
    assign _21193 = _21192[62:0];
    assign _21201 = { _21193,
                      _21200 };
    assign _21202 = _21201[62:0];
    assign _21210 = { _21202,
                      _21209 };
    assign _21211 = _21210[62:0];
    assign _21219 = { _21211,
                      _21218 };
    assign _21220 = _21219[62:0];
    assign _21228 = { _21220,
                      _21227 };
    assign _21229 = _21228[62:0];
    assign _21237 = { _21229,
                      _21236 };
    assign _21238 = _21237[62:0];
    assign _21246 = { _21238,
                      _21245 };
    assign _21247 = _21246[62:0];
    assign _21255 = { _21247,
                      _21254 };
    assign _21256 = _21255[62:0];
    assign _21264 = { _21256,
                      _21263 };
    assign _21265 = _21264[62:0];
    assign _21273 = { _21265,
                      _21272 };
    assign _21274 = _21273[62:0];
    assign _21282 = { _21274,
                      _21281 };
    assign _21283 = _21282[62:0];
    assign _21291 = { _21283,
                      _21290 };
    assign _21292 = _21291[62:0];
    assign _21300 = { _21292,
                      _21299 };
    assign _21301 = _21300[62:0];
    assign _21309 = { _21301,
                      _21308 };
    assign _21310 = _21309[62:0];
    assign _21318 = { _21310,
                      _21317 };
    assign _21319 = _21318[62:0];
    assign _21327 = { _21319,
                      _21326 };
    assign _21328 = _21327[62:0];
    assign _21336 = { _21328,
                      _21335 };
    assign _21337 = _21336[62:0];
    assign _21345 = { _21337,
                      _21344 };
    assign _21346 = _21345[62:0];
    assign _21354 = { _21346,
                      _21353 };
    assign _21355 = _21354[62:0];
    assign _21363 = { _21355,
                      _21362 };
    assign _21364 = _21363[62:0];
    assign _21372 = { _21364,
                      _21371 };
    assign _21373 = _21372[62:0];
    assign _21381 = { _21373,
                      _21380 };
    assign _21382 = _21381[62:0];
    assign _21390 = { _21382,
                      _21389 };
    assign _21391 = _21390[62:0];
    assign _21399 = { _21391,
                      _21398 };
    assign _21400 = _21399[62:0];
    assign _21408 = { _21400,
                      _21407 };
    assign _21409 = _21408[62:0];
    assign _21417 = { _21409,
                      _21416 };
    assign _21418 = _21417[62:0];
    assign _21426 = { _21418,
                      _21425 };
    assign _21427 = _21426[62:0];
    assign _21435 = { _21427,
                      _21434 };
    assign _21436 = _21435[62:0];
    assign _21444 = { _21436,
                      _21443 };
    assign _21445 = _21444[62:0];
    assign _21453 = { _21445,
                      _21452 };
    assign _21454 = _21453[62:0];
    assign _21462 = { _21454,
                      _21461 };
    assign _21463 = _21462[62:0];
    assign _21471 = { _21463,
                      _21470 };
    assign _21472 = _21471[62:0];
    assign _21480 = { _21472,
                      _21479 };
    assign _21481 = _21480[62:0];
    assign _21489 = { _21481,
                      _21488 };
    assign _21490 = _21489[62:0];
    assign _21498 = { _21490,
                      _21497 };
    assign _21499 = _21498[62:0];
    assign _21507 = { _21499,
                      _21506 };
    assign _21508 = _21507[62:0];
    assign _21516 = { _21508,
                      _21515 };
    assign _21517 = _21516[62:0];
    assign _21525 = { _21517,
                      _21524 };
    assign _21526 = _21525[62:0];
    assign _21534 = { _21526,
                      _21533 };
    assign _21535 = _21534[62:0];
    assign _21543 = { _21535,
                      _21542 };
    assign _21544 = _21543[62:0];
    assign _21552 = { _21544,
                      _21551 };
    assign _21553 = _21552[62:0];
    assign _21561 = { _21553,
                      _21560 };
    assign _21562 = _21561[62:0];
    assign _21570 = { _21562,
                      _21569 };
    assign _21571 = _21570[62:0];
    assign _21579 = { _21571,
                      _21578 };
    assign _21580 = _21579[62:0];
    assign _21588 = { _21580,
                      _21587 };
    assign _21589 = _21588[62:0];
    assign _21597 = { _21589,
                      _21596 };
    assign _21598 = _21597 * _21027;
    assign _21599 = _21598[63:0];
    assign _21600 = _21027 < _21599;
    assign _21601 = _21600 ? _21599 : _21027;
    assign _21017 = 64'b0000000000000000000000000000001001010100000010111110001111111111;
    assign _21018 = _5 < _21017;
    assign _21019 = _21018 ? _5 : _21017;
    assign _21602 = _21019 < _21601;
    assign _21603 = ~ _21602;
    assign _22766 = _21603 ? _22765 : _21604;
    assign _21008 = _20439[0:0];
    assign _21005 = _21000 - _22192;
    assign _21006 = _21002 ? _21005 : _21000;
    assign _21007 = _21006[62:0];
    assign _21009 = { _21007,
                      _21008 };
    assign _21010 = _21009 < _22192;
    assign _21011 = ~ _21010;
    assign _20999 = _20439[1:1];
    assign _20996 = _20991 - _22192;
    assign _20997 = _20993 ? _20996 : _20991;
    assign _20998 = _20997[62:0];
    assign _21000 = { _20998,
                      _20999 };
    assign _21001 = _21000 < _22192;
    assign _21002 = ~ _21001;
    assign _20990 = _20439[2:2];
    assign _20987 = _20982 - _22192;
    assign _20988 = _20984 ? _20987 : _20982;
    assign _20989 = _20988[62:0];
    assign _20991 = { _20989,
                      _20990 };
    assign _20992 = _20991 < _22192;
    assign _20993 = ~ _20992;
    assign _20981 = _20439[3:3];
    assign _20978 = _20973 - _22192;
    assign _20979 = _20975 ? _20978 : _20973;
    assign _20980 = _20979[62:0];
    assign _20982 = { _20980,
                      _20981 };
    assign _20983 = _20982 < _22192;
    assign _20984 = ~ _20983;
    assign _20972 = _20439[4:4];
    assign _20969 = _20964 - _22192;
    assign _20970 = _20966 ? _20969 : _20964;
    assign _20971 = _20970[62:0];
    assign _20973 = { _20971,
                      _20972 };
    assign _20974 = _20973 < _22192;
    assign _20975 = ~ _20974;
    assign _20963 = _20439[5:5];
    assign _20960 = _20955 - _22192;
    assign _20961 = _20957 ? _20960 : _20955;
    assign _20962 = _20961[62:0];
    assign _20964 = { _20962,
                      _20963 };
    assign _20965 = _20964 < _22192;
    assign _20966 = ~ _20965;
    assign _20954 = _20439[6:6];
    assign _20951 = _20946 - _22192;
    assign _20952 = _20948 ? _20951 : _20946;
    assign _20953 = _20952[62:0];
    assign _20955 = { _20953,
                      _20954 };
    assign _20956 = _20955 < _22192;
    assign _20957 = ~ _20956;
    assign _20945 = _20439[7:7];
    assign _20942 = _20937 - _22192;
    assign _20943 = _20939 ? _20942 : _20937;
    assign _20944 = _20943[62:0];
    assign _20946 = { _20944,
                      _20945 };
    assign _20947 = _20946 < _22192;
    assign _20948 = ~ _20947;
    assign _20936 = _20439[8:8];
    assign _20933 = _20928 - _22192;
    assign _20934 = _20930 ? _20933 : _20928;
    assign _20935 = _20934[62:0];
    assign _20937 = { _20935,
                      _20936 };
    assign _20938 = _20937 < _22192;
    assign _20939 = ~ _20938;
    assign _20927 = _20439[9:9];
    assign _20924 = _20919 - _22192;
    assign _20925 = _20921 ? _20924 : _20919;
    assign _20926 = _20925[62:0];
    assign _20928 = { _20926,
                      _20927 };
    assign _20929 = _20928 < _22192;
    assign _20930 = ~ _20929;
    assign _20918 = _20439[10:10];
    assign _20915 = _20910 - _22192;
    assign _20916 = _20912 ? _20915 : _20910;
    assign _20917 = _20916[62:0];
    assign _20919 = { _20917,
                      _20918 };
    assign _20920 = _20919 < _22192;
    assign _20921 = ~ _20920;
    assign _20909 = _20439[11:11];
    assign _20906 = _20901 - _22192;
    assign _20907 = _20903 ? _20906 : _20901;
    assign _20908 = _20907[62:0];
    assign _20910 = { _20908,
                      _20909 };
    assign _20911 = _20910 < _22192;
    assign _20912 = ~ _20911;
    assign _20900 = _20439[12:12];
    assign _20897 = _20892 - _22192;
    assign _20898 = _20894 ? _20897 : _20892;
    assign _20899 = _20898[62:0];
    assign _20901 = { _20899,
                      _20900 };
    assign _20902 = _20901 < _22192;
    assign _20903 = ~ _20902;
    assign _20891 = _20439[13:13];
    assign _20888 = _20883 - _22192;
    assign _20889 = _20885 ? _20888 : _20883;
    assign _20890 = _20889[62:0];
    assign _20892 = { _20890,
                      _20891 };
    assign _20893 = _20892 < _22192;
    assign _20894 = ~ _20893;
    assign _20882 = _20439[14:14];
    assign _20879 = _20874 - _22192;
    assign _20880 = _20876 ? _20879 : _20874;
    assign _20881 = _20880[62:0];
    assign _20883 = { _20881,
                      _20882 };
    assign _20884 = _20883 < _22192;
    assign _20885 = ~ _20884;
    assign _20873 = _20439[15:15];
    assign _20870 = _20865 - _22192;
    assign _20871 = _20867 ? _20870 : _20865;
    assign _20872 = _20871[62:0];
    assign _20874 = { _20872,
                      _20873 };
    assign _20875 = _20874 < _22192;
    assign _20876 = ~ _20875;
    assign _20864 = _20439[16:16];
    assign _20861 = _20856 - _22192;
    assign _20862 = _20858 ? _20861 : _20856;
    assign _20863 = _20862[62:0];
    assign _20865 = { _20863,
                      _20864 };
    assign _20866 = _20865 < _22192;
    assign _20867 = ~ _20866;
    assign _20855 = _20439[17:17];
    assign _20852 = _20847 - _22192;
    assign _20853 = _20849 ? _20852 : _20847;
    assign _20854 = _20853[62:0];
    assign _20856 = { _20854,
                      _20855 };
    assign _20857 = _20856 < _22192;
    assign _20858 = ~ _20857;
    assign _20846 = _20439[18:18];
    assign _20843 = _20838 - _22192;
    assign _20844 = _20840 ? _20843 : _20838;
    assign _20845 = _20844[62:0];
    assign _20847 = { _20845,
                      _20846 };
    assign _20848 = _20847 < _22192;
    assign _20849 = ~ _20848;
    assign _20837 = _20439[19:19];
    assign _20834 = _20829 - _22192;
    assign _20835 = _20831 ? _20834 : _20829;
    assign _20836 = _20835[62:0];
    assign _20838 = { _20836,
                      _20837 };
    assign _20839 = _20838 < _22192;
    assign _20840 = ~ _20839;
    assign _20828 = _20439[20:20];
    assign _20825 = _20820 - _22192;
    assign _20826 = _20822 ? _20825 : _20820;
    assign _20827 = _20826[62:0];
    assign _20829 = { _20827,
                      _20828 };
    assign _20830 = _20829 < _22192;
    assign _20831 = ~ _20830;
    assign _20819 = _20439[21:21];
    assign _20816 = _20811 - _22192;
    assign _20817 = _20813 ? _20816 : _20811;
    assign _20818 = _20817[62:0];
    assign _20820 = { _20818,
                      _20819 };
    assign _20821 = _20820 < _22192;
    assign _20822 = ~ _20821;
    assign _20810 = _20439[22:22];
    assign _20807 = _20802 - _22192;
    assign _20808 = _20804 ? _20807 : _20802;
    assign _20809 = _20808[62:0];
    assign _20811 = { _20809,
                      _20810 };
    assign _20812 = _20811 < _22192;
    assign _20813 = ~ _20812;
    assign _20801 = _20439[23:23];
    assign _20798 = _20793 - _22192;
    assign _20799 = _20795 ? _20798 : _20793;
    assign _20800 = _20799[62:0];
    assign _20802 = { _20800,
                      _20801 };
    assign _20803 = _20802 < _22192;
    assign _20804 = ~ _20803;
    assign _20792 = _20439[24:24];
    assign _20789 = _20784 - _22192;
    assign _20790 = _20786 ? _20789 : _20784;
    assign _20791 = _20790[62:0];
    assign _20793 = { _20791,
                      _20792 };
    assign _20794 = _20793 < _22192;
    assign _20795 = ~ _20794;
    assign _20783 = _20439[25:25];
    assign _20780 = _20775 - _22192;
    assign _20781 = _20777 ? _20780 : _20775;
    assign _20782 = _20781[62:0];
    assign _20784 = { _20782,
                      _20783 };
    assign _20785 = _20784 < _22192;
    assign _20786 = ~ _20785;
    assign _20774 = _20439[26:26];
    assign _20771 = _20766 - _22192;
    assign _20772 = _20768 ? _20771 : _20766;
    assign _20773 = _20772[62:0];
    assign _20775 = { _20773,
                      _20774 };
    assign _20776 = _20775 < _22192;
    assign _20777 = ~ _20776;
    assign _20765 = _20439[27:27];
    assign _20762 = _20757 - _22192;
    assign _20763 = _20759 ? _20762 : _20757;
    assign _20764 = _20763[62:0];
    assign _20766 = { _20764,
                      _20765 };
    assign _20767 = _20766 < _22192;
    assign _20768 = ~ _20767;
    assign _20756 = _20439[28:28];
    assign _20753 = _20748 - _22192;
    assign _20754 = _20750 ? _20753 : _20748;
    assign _20755 = _20754[62:0];
    assign _20757 = { _20755,
                      _20756 };
    assign _20758 = _20757 < _22192;
    assign _20759 = ~ _20758;
    assign _20747 = _20439[29:29];
    assign _20744 = _20739 - _22192;
    assign _20745 = _20741 ? _20744 : _20739;
    assign _20746 = _20745[62:0];
    assign _20748 = { _20746,
                      _20747 };
    assign _20749 = _20748 < _22192;
    assign _20750 = ~ _20749;
    assign _20738 = _20439[30:30];
    assign _20735 = _20730 - _22192;
    assign _20736 = _20732 ? _20735 : _20730;
    assign _20737 = _20736[62:0];
    assign _20739 = { _20737,
                      _20738 };
    assign _20740 = _20739 < _22192;
    assign _20741 = ~ _20740;
    assign _20729 = _20439[31:31];
    assign _20726 = _20721 - _22192;
    assign _20727 = _20723 ? _20726 : _20721;
    assign _20728 = _20727[62:0];
    assign _20730 = { _20728,
                      _20729 };
    assign _20731 = _20730 < _22192;
    assign _20732 = ~ _20731;
    assign _20720 = _20439[32:32];
    assign _20717 = _20712 - _22192;
    assign _20718 = _20714 ? _20717 : _20712;
    assign _20719 = _20718[62:0];
    assign _20721 = { _20719,
                      _20720 };
    assign _20722 = _20721 < _22192;
    assign _20723 = ~ _20722;
    assign _20711 = _20439[33:33];
    assign _20708 = _20703 - _22192;
    assign _20709 = _20705 ? _20708 : _20703;
    assign _20710 = _20709[62:0];
    assign _20712 = { _20710,
                      _20711 };
    assign _20713 = _20712 < _22192;
    assign _20714 = ~ _20713;
    assign _20702 = _20439[34:34];
    assign _20699 = _20694 - _22192;
    assign _20700 = _20696 ? _20699 : _20694;
    assign _20701 = _20700[62:0];
    assign _20703 = { _20701,
                      _20702 };
    assign _20704 = _20703 < _22192;
    assign _20705 = ~ _20704;
    assign _20693 = _20439[35:35];
    assign _20690 = _20685 - _22192;
    assign _20691 = _20687 ? _20690 : _20685;
    assign _20692 = _20691[62:0];
    assign _20694 = { _20692,
                      _20693 };
    assign _20695 = _20694 < _22192;
    assign _20696 = ~ _20695;
    assign _20684 = _20439[36:36];
    assign _20681 = _20676 - _22192;
    assign _20682 = _20678 ? _20681 : _20676;
    assign _20683 = _20682[62:0];
    assign _20685 = { _20683,
                      _20684 };
    assign _20686 = _20685 < _22192;
    assign _20687 = ~ _20686;
    assign _20675 = _20439[37:37];
    assign _20672 = _20667 - _22192;
    assign _20673 = _20669 ? _20672 : _20667;
    assign _20674 = _20673[62:0];
    assign _20676 = { _20674,
                      _20675 };
    assign _20677 = _20676 < _22192;
    assign _20678 = ~ _20677;
    assign _20666 = _20439[38:38];
    assign _20663 = _20658 - _22192;
    assign _20664 = _20660 ? _20663 : _20658;
    assign _20665 = _20664[62:0];
    assign _20667 = { _20665,
                      _20666 };
    assign _20668 = _20667 < _22192;
    assign _20669 = ~ _20668;
    assign _20657 = _20439[39:39];
    assign _20654 = _20649 - _22192;
    assign _20655 = _20651 ? _20654 : _20649;
    assign _20656 = _20655[62:0];
    assign _20658 = { _20656,
                      _20657 };
    assign _20659 = _20658 < _22192;
    assign _20660 = ~ _20659;
    assign _20648 = _20439[40:40];
    assign _20645 = _20640 - _22192;
    assign _20646 = _20642 ? _20645 : _20640;
    assign _20647 = _20646[62:0];
    assign _20649 = { _20647,
                      _20648 };
    assign _20650 = _20649 < _22192;
    assign _20651 = ~ _20650;
    assign _20639 = _20439[41:41];
    assign _20636 = _20631 - _22192;
    assign _20637 = _20633 ? _20636 : _20631;
    assign _20638 = _20637[62:0];
    assign _20640 = { _20638,
                      _20639 };
    assign _20641 = _20640 < _22192;
    assign _20642 = ~ _20641;
    assign _20630 = _20439[42:42];
    assign _20627 = _20622 - _22192;
    assign _20628 = _20624 ? _20627 : _20622;
    assign _20629 = _20628[62:0];
    assign _20631 = { _20629,
                      _20630 };
    assign _20632 = _20631 < _22192;
    assign _20633 = ~ _20632;
    assign _20621 = _20439[43:43];
    assign _20618 = _20613 - _22192;
    assign _20619 = _20615 ? _20618 : _20613;
    assign _20620 = _20619[62:0];
    assign _20622 = { _20620,
                      _20621 };
    assign _20623 = _20622 < _22192;
    assign _20624 = ~ _20623;
    assign _20612 = _20439[44:44];
    assign _20609 = _20604 - _22192;
    assign _20610 = _20606 ? _20609 : _20604;
    assign _20611 = _20610[62:0];
    assign _20613 = { _20611,
                      _20612 };
    assign _20614 = _20613 < _22192;
    assign _20615 = ~ _20614;
    assign _20603 = _20439[45:45];
    assign _20600 = _20595 - _22192;
    assign _20601 = _20597 ? _20600 : _20595;
    assign _20602 = _20601[62:0];
    assign _20604 = { _20602,
                      _20603 };
    assign _20605 = _20604 < _22192;
    assign _20606 = ~ _20605;
    assign _20594 = _20439[46:46];
    assign _20591 = _20586 - _22192;
    assign _20592 = _20588 ? _20591 : _20586;
    assign _20593 = _20592[62:0];
    assign _20595 = { _20593,
                      _20594 };
    assign _20596 = _20595 < _22192;
    assign _20597 = ~ _20596;
    assign _20585 = _20439[47:47];
    assign _20582 = _20577 - _22192;
    assign _20583 = _20579 ? _20582 : _20577;
    assign _20584 = _20583[62:0];
    assign _20586 = { _20584,
                      _20585 };
    assign _20587 = _20586 < _22192;
    assign _20588 = ~ _20587;
    assign _20576 = _20439[48:48];
    assign _20573 = _20568 - _22192;
    assign _20574 = _20570 ? _20573 : _20568;
    assign _20575 = _20574[62:0];
    assign _20577 = { _20575,
                      _20576 };
    assign _20578 = _20577 < _22192;
    assign _20579 = ~ _20578;
    assign _20567 = _20439[49:49];
    assign _20564 = _20559 - _22192;
    assign _20565 = _20561 ? _20564 : _20559;
    assign _20566 = _20565[62:0];
    assign _20568 = { _20566,
                      _20567 };
    assign _20569 = _20568 < _22192;
    assign _20570 = ~ _20569;
    assign _20558 = _20439[50:50];
    assign _20555 = _20550 - _22192;
    assign _20556 = _20552 ? _20555 : _20550;
    assign _20557 = _20556[62:0];
    assign _20559 = { _20557,
                      _20558 };
    assign _20560 = _20559 < _22192;
    assign _20561 = ~ _20560;
    assign _20549 = _20439[51:51];
    assign _20546 = _20541 - _22192;
    assign _20547 = _20543 ? _20546 : _20541;
    assign _20548 = _20547[62:0];
    assign _20550 = { _20548,
                      _20549 };
    assign _20551 = _20550 < _22192;
    assign _20552 = ~ _20551;
    assign _20540 = _20439[52:52];
    assign _20537 = _20532 - _22192;
    assign _20538 = _20534 ? _20537 : _20532;
    assign _20539 = _20538[62:0];
    assign _20541 = { _20539,
                      _20540 };
    assign _20542 = _20541 < _22192;
    assign _20543 = ~ _20542;
    assign _20531 = _20439[53:53];
    assign _20528 = _20523 - _22192;
    assign _20529 = _20525 ? _20528 : _20523;
    assign _20530 = _20529[62:0];
    assign _20532 = { _20530,
                      _20531 };
    assign _20533 = _20532 < _22192;
    assign _20534 = ~ _20533;
    assign _20522 = _20439[54:54];
    assign _20519 = _20514 - _22192;
    assign _20520 = _20516 ? _20519 : _20514;
    assign _20521 = _20520[62:0];
    assign _20523 = { _20521,
                      _20522 };
    assign _20524 = _20523 < _22192;
    assign _20525 = ~ _20524;
    assign _20513 = _20439[55:55];
    assign _20510 = _20505 - _22192;
    assign _20511 = _20507 ? _20510 : _20505;
    assign _20512 = _20511[62:0];
    assign _20514 = { _20512,
                      _20513 };
    assign _20515 = _20514 < _22192;
    assign _20516 = ~ _20515;
    assign _20504 = _20439[56:56];
    assign _20501 = _20496 - _22192;
    assign _20502 = _20498 ? _20501 : _20496;
    assign _20503 = _20502[62:0];
    assign _20505 = { _20503,
                      _20504 };
    assign _20506 = _20505 < _22192;
    assign _20507 = ~ _20506;
    assign _20495 = _20439[57:57];
    assign _20492 = _20487 - _22192;
    assign _20493 = _20489 ? _20492 : _20487;
    assign _20494 = _20493[62:0];
    assign _20496 = { _20494,
                      _20495 };
    assign _20497 = _20496 < _22192;
    assign _20498 = ~ _20497;
    assign _20486 = _20439[58:58];
    assign _20483 = _20478 - _22192;
    assign _20484 = _20480 ? _20483 : _20478;
    assign _20485 = _20484[62:0];
    assign _20487 = { _20485,
                      _20486 };
    assign _20488 = _20487 < _22192;
    assign _20489 = ~ _20488;
    assign _20477 = _20439[59:59];
    assign _20474 = _20469 - _22192;
    assign _20475 = _20471 ? _20474 : _20469;
    assign _20476 = _20475[62:0];
    assign _20478 = { _20476,
                      _20477 };
    assign _20479 = _20478 < _22192;
    assign _20480 = ~ _20479;
    assign _20468 = _20439[60:60];
    assign _20465 = _20460 - _22192;
    assign _20466 = _20462 ? _20465 : _20460;
    assign _20467 = _20466[62:0];
    assign _20469 = { _20467,
                      _20468 };
    assign _20470 = _20469 < _22192;
    assign _20471 = ~ _20470;
    assign _20459 = _20439[61:61];
    assign _20456 = _20451 - _22192;
    assign _20457 = _20453 ? _20456 : _20451;
    assign _20458 = _20457[62:0];
    assign _20460 = { _20458,
                      _20459 };
    assign _20461 = _20460 < _22192;
    assign _20462 = ~ _20461;
    assign _20450 = _20439[62:62];
    assign _20447 = _20441 - _22192;
    assign _20448 = _20444 ? _20447 : _20441;
    assign _20449 = _20448[62:0];
    assign _20451 = { _20449,
                      _20450 };
    assign _20452 = _20451 < _22192;
    assign _20453 = ~ _20452;
    assign _20437 = _20429 + _22186;
    assign _20438 = _20429 * _20437;
    assign _20439 = _20438[63:0];
    assign _20440 = _20439[63:63];
    assign _20441 = { _22185,
                      _20440 };
    assign _20443 = _20441 < _22192;
    assign _20444 = ~ _20443;
    assign _20445 = { _22185,
                      _20444 };
    assign _20446 = _20445[62:0];
    assign _20454 = { _20446,
                      _20453 };
    assign _20455 = _20454[62:0];
    assign _20463 = { _20455,
                      _20462 };
    assign _20464 = _20463[62:0];
    assign _20472 = { _20464,
                      _20471 };
    assign _20473 = _20472[62:0];
    assign _20481 = { _20473,
                      _20480 };
    assign _20482 = _20481[62:0];
    assign _20490 = { _20482,
                      _20489 };
    assign _20491 = _20490[62:0];
    assign _20499 = { _20491,
                      _20498 };
    assign _20500 = _20499[62:0];
    assign _20508 = { _20500,
                      _20507 };
    assign _20509 = _20508[62:0];
    assign _20517 = { _20509,
                      _20516 };
    assign _20518 = _20517[62:0];
    assign _20526 = { _20518,
                      _20525 };
    assign _20527 = _20526[62:0];
    assign _20535 = { _20527,
                      _20534 };
    assign _20536 = _20535[62:0];
    assign _20544 = { _20536,
                      _20543 };
    assign _20545 = _20544[62:0];
    assign _20553 = { _20545,
                      _20552 };
    assign _20554 = _20553[62:0];
    assign _20562 = { _20554,
                      _20561 };
    assign _20563 = _20562[62:0];
    assign _20571 = { _20563,
                      _20570 };
    assign _20572 = _20571[62:0];
    assign _20580 = { _20572,
                      _20579 };
    assign _20581 = _20580[62:0];
    assign _20589 = { _20581,
                      _20588 };
    assign _20590 = _20589[62:0];
    assign _20598 = { _20590,
                      _20597 };
    assign _20599 = _20598[62:0];
    assign _20607 = { _20599,
                      _20606 };
    assign _20608 = _20607[62:0];
    assign _20616 = { _20608,
                      _20615 };
    assign _20617 = _20616[62:0];
    assign _20625 = { _20617,
                      _20624 };
    assign _20626 = _20625[62:0];
    assign _20634 = { _20626,
                      _20633 };
    assign _20635 = _20634[62:0];
    assign _20643 = { _20635,
                      _20642 };
    assign _20644 = _20643[62:0];
    assign _20652 = { _20644,
                      _20651 };
    assign _20653 = _20652[62:0];
    assign _20661 = { _20653,
                      _20660 };
    assign _20662 = _20661[62:0];
    assign _20670 = { _20662,
                      _20669 };
    assign _20671 = _20670[62:0];
    assign _20679 = { _20671,
                      _20678 };
    assign _20680 = _20679[62:0];
    assign _20688 = { _20680,
                      _20687 };
    assign _20689 = _20688[62:0];
    assign _20697 = { _20689,
                      _20696 };
    assign _20698 = _20697[62:0];
    assign _20706 = { _20698,
                      _20705 };
    assign _20707 = _20706[62:0];
    assign _20715 = { _20707,
                      _20714 };
    assign _20716 = _20715[62:0];
    assign _20724 = { _20716,
                      _20723 };
    assign _20725 = _20724[62:0];
    assign _20733 = { _20725,
                      _20732 };
    assign _20734 = _20733[62:0];
    assign _20742 = { _20734,
                      _20741 };
    assign _20743 = _20742[62:0];
    assign _20751 = { _20743,
                      _20750 };
    assign _20752 = _20751[62:0];
    assign _20760 = { _20752,
                      _20759 };
    assign _20761 = _20760[62:0];
    assign _20769 = { _20761,
                      _20768 };
    assign _20770 = _20769[62:0];
    assign _20778 = { _20770,
                      _20777 };
    assign _20779 = _20778[62:0];
    assign _20787 = { _20779,
                      _20786 };
    assign _20788 = _20787[62:0];
    assign _20796 = { _20788,
                      _20795 };
    assign _20797 = _20796[62:0];
    assign _20805 = { _20797,
                      _20804 };
    assign _20806 = _20805[62:0];
    assign _20814 = { _20806,
                      _20813 };
    assign _20815 = _20814[62:0];
    assign _20823 = { _20815,
                      _20822 };
    assign _20824 = _20823[62:0];
    assign _20832 = { _20824,
                      _20831 };
    assign _20833 = _20832[62:0];
    assign _20841 = { _20833,
                      _20840 };
    assign _20842 = _20841[62:0];
    assign _20850 = { _20842,
                      _20849 };
    assign _20851 = _20850[62:0];
    assign _20859 = { _20851,
                      _20858 };
    assign _20860 = _20859[62:0];
    assign _20868 = { _20860,
                      _20867 };
    assign _20869 = _20868[62:0];
    assign _20877 = { _20869,
                      _20876 };
    assign _20878 = _20877[62:0];
    assign _20886 = { _20878,
                      _20885 };
    assign _20887 = _20886[62:0];
    assign _20895 = { _20887,
                      _20894 };
    assign _20896 = _20895[62:0];
    assign _20904 = { _20896,
                      _20903 };
    assign _20905 = _20904[62:0];
    assign _20913 = { _20905,
                      _20912 };
    assign _20914 = _20913[62:0];
    assign _20922 = { _20914,
                      _20921 };
    assign _20923 = _20922[62:0];
    assign _20931 = { _20923,
                      _20930 };
    assign _20932 = _20931[62:0];
    assign _20940 = { _20932,
                      _20939 };
    assign _20941 = _20940[62:0];
    assign _20949 = { _20941,
                      _20948 };
    assign _20950 = _20949[62:0];
    assign _20958 = { _20950,
                      _20957 };
    assign _20959 = _20958[62:0];
    assign _20967 = { _20959,
                      _20966 };
    assign _20968 = _20967[62:0];
    assign _20976 = { _20968,
                      _20975 };
    assign _20977 = _20976[62:0];
    assign _20985 = { _20977,
                      _20984 };
    assign _20986 = _20985[62:0];
    assign _20994 = { _20986,
                      _20993 };
    assign _20995 = _20994[62:0];
    assign _21003 = { _20995,
                      _21002 };
    assign _21004 = _21003[62:0];
    assign _21012 = { _21004,
                      _21011 };
    assign _21013 = _19277 * _21012;
    assign _21014 = _21013[63:0];
    assign _20425 = _19857[0:0];
    assign _20422 = _20417 - _19277;
    assign _20423 = _20419 ? _20422 : _20417;
    assign _20424 = _20423[62:0];
    assign _20426 = { _20424,
                      _20425 };
    assign _20427 = _20426 < _19277;
    assign _20428 = ~ _20427;
    assign _20416 = _19857[1:1];
    assign _20413 = _20408 - _19277;
    assign _20414 = _20410 ? _20413 : _20408;
    assign _20415 = _20414[62:0];
    assign _20417 = { _20415,
                      _20416 };
    assign _20418 = _20417 < _19277;
    assign _20419 = ~ _20418;
    assign _20407 = _19857[2:2];
    assign _20404 = _20399 - _19277;
    assign _20405 = _20401 ? _20404 : _20399;
    assign _20406 = _20405[62:0];
    assign _20408 = { _20406,
                      _20407 };
    assign _20409 = _20408 < _19277;
    assign _20410 = ~ _20409;
    assign _20398 = _19857[3:3];
    assign _20395 = _20390 - _19277;
    assign _20396 = _20392 ? _20395 : _20390;
    assign _20397 = _20396[62:0];
    assign _20399 = { _20397,
                      _20398 };
    assign _20400 = _20399 < _19277;
    assign _20401 = ~ _20400;
    assign _20389 = _19857[4:4];
    assign _20386 = _20381 - _19277;
    assign _20387 = _20383 ? _20386 : _20381;
    assign _20388 = _20387[62:0];
    assign _20390 = { _20388,
                      _20389 };
    assign _20391 = _20390 < _19277;
    assign _20392 = ~ _20391;
    assign _20380 = _19857[5:5];
    assign _20377 = _20372 - _19277;
    assign _20378 = _20374 ? _20377 : _20372;
    assign _20379 = _20378[62:0];
    assign _20381 = { _20379,
                      _20380 };
    assign _20382 = _20381 < _19277;
    assign _20383 = ~ _20382;
    assign _20371 = _19857[6:6];
    assign _20368 = _20363 - _19277;
    assign _20369 = _20365 ? _20368 : _20363;
    assign _20370 = _20369[62:0];
    assign _20372 = { _20370,
                      _20371 };
    assign _20373 = _20372 < _19277;
    assign _20374 = ~ _20373;
    assign _20362 = _19857[7:7];
    assign _20359 = _20354 - _19277;
    assign _20360 = _20356 ? _20359 : _20354;
    assign _20361 = _20360[62:0];
    assign _20363 = { _20361,
                      _20362 };
    assign _20364 = _20363 < _19277;
    assign _20365 = ~ _20364;
    assign _20353 = _19857[8:8];
    assign _20350 = _20345 - _19277;
    assign _20351 = _20347 ? _20350 : _20345;
    assign _20352 = _20351[62:0];
    assign _20354 = { _20352,
                      _20353 };
    assign _20355 = _20354 < _19277;
    assign _20356 = ~ _20355;
    assign _20344 = _19857[9:9];
    assign _20341 = _20336 - _19277;
    assign _20342 = _20338 ? _20341 : _20336;
    assign _20343 = _20342[62:0];
    assign _20345 = { _20343,
                      _20344 };
    assign _20346 = _20345 < _19277;
    assign _20347 = ~ _20346;
    assign _20335 = _19857[10:10];
    assign _20332 = _20327 - _19277;
    assign _20333 = _20329 ? _20332 : _20327;
    assign _20334 = _20333[62:0];
    assign _20336 = { _20334,
                      _20335 };
    assign _20337 = _20336 < _19277;
    assign _20338 = ~ _20337;
    assign _20326 = _19857[11:11];
    assign _20323 = _20318 - _19277;
    assign _20324 = _20320 ? _20323 : _20318;
    assign _20325 = _20324[62:0];
    assign _20327 = { _20325,
                      _20326 };
    assign _20328 = _20327 < _19277;
    assign _20329 = ~ _20328;
    assign _20317 = _19857[12:12];
    assign _20314 = _20309 - _19277;
    assign _20315 = _20311 ? _20314 : _20309;
    assign _20316 = _20315[62:0];
    assign _20318 = { _20316,
                      _20317 };
    assign _20319 = _20318 < _19277;
    assign _20320 = ~ _20319;
    assign _20308 = _19857[13:13];
    assign _20305 = _20300 - _19277;
    assign _20306 = _20302 ? _20305 : _20300;
    assign _20307 = _20306[62:0];
    assign _20309 = { _20307,
                      _20308 };
    assign _20310 = _20309 < _19277;
    assign _20311 = ~ _20310;
    assign _20299 = _19857[14:14];
    assign _20296 = _20291 - _19277;
    assign _20297 = _20293 ? _20296 : _20291;
    assign _20298 = _20297[62:0];
    assign _20300 = { _20298,
                      _20299 };
    assign _20301 = _20300 < _19277;
    assign _20302 = ~ _20301;
    assign _20290 = _19857[15:15];
    assign _20287 = _20282 - _19277;
    assign _20288 = _20284 ? _20287 : _20282;
    assign _20289 = _20288[62:0];
    assign _20291 = { _20289,
                      _20290 };
    assign _20292 = _20291 < _19277;
    assign _20293 = ~ _20292;
    assign _20281 = _19857[16:16];
    assign _20278 = _20273 - _19277;
    assign _20279 = _20275 ? _20278 : _20273;
    assign _20280 = _20279[62:0];
    assign _20282 = { _20280,
                      _20281 };
    assign _20283 = _20282 < _19277;
    assign _20284 = ~ _20283;
    assign _20272 = _19857[17:17];
    assign _20269 = _20264 - _19277;
    assign _20270 = _20266 ? _20269 : _20264;
    assign _20271 = _20270[62:0];
    assign _20273 = { _20271,
                      _20272 };
    assign _20274 = _20273 < _19277;
    assign _20275 = ~ _20274;
    assign _20263 = _19857[18:18];
    assign _20260 = _20255 - _19277;
    assign _20261 = _20257 ? _20260 : _20255;
    assign _20262 = _20261[62:0];
    assign _20264 = { _20262,
                      _20263 };
    assign _20265 = _20264 < _19277;
    assign _20266 = ~ _20265;
    assign _20254 = _19857[19:19];
    assign _20251 = _20246 - _19277;
    assign _20252 = _20248 ? _20251 : _20246;
    assign _20253 = _20252[62:0];
    assign _20255 = { _20253,
                      _20254 };
    assign _20256 = _20255 < _19277;
    assign _20257 = ~ _20256;
    assign _20245 = _19857[20:20];
    assign _20242 = _20237 - _19277;
    assign _20243 = _20239 ? _20242 : _20237;
    assign _20244 = _20243[62:0];
    assign _20246 = { _20244,
                      _20245 };
    assign _20247 = _20246 < _19277;
    assign _20248 = ~ _20247;
    assign _20236 = _19857[21:21];
    assign _20233 = _20228 - _19277;
    assign _20234 = _20230 ? _20233 : _20228;
    assign _20235 = _20234[62:0];
    assign _20237 = { _20235,
                      _20236 };
    assign _20238 = _20237 < _19277;
    assign _20239 = ~ _20238;
    assign _20227 = _19857[22:22];
    assign _20224 = _20219 - _19277;
    assign _20225 = _20221 ? _20224 : _20219;
    assign _20226 = _20225[62:0];
    assign _20228 = { _20226,
                      _20227 };
    assign _20229 = _20228 < _19277;
    assign _20230 = ~ _20229;
    assign _20218 = _19857[23:23];
    assign _20215 = _20210 - _19277;
    assign _20216 = _20212 ? _20215 : _20210;
    assign _20217 = _20216[62:0];
    assign _20219 = { _20217,
                      _20218 };
    assign _20220 = _20219 < _19277;
    assign _20221 = ~ _20220;
    assign _20209 = _19857[24:24];
    assign _20206 = _20201 - _19277;
    assign _20207 = _20203 ? _20206 : _20201;
    assign _20208 = _20207[62:0];
    assign _20210 = { _20208,
                      _20209 };
    assign _20211 = _20210 < _19277;
    assign _20212 = ~ _20211;
    assign _20200 = _19857[25:25];
    assign _20197 = _20192 - _19277;
    assign _20198 = _20194 ? _20197 : _20192;
    assign _20199 = _20198[62:0];
    assign _20201 = { _20199,
                      _20200 };
    assign _20202 = _20201 < _19277;
    assign _20203 = ~ _20202;
    assign _20191 = _19857[26:26];
    assign _20188 = _20183 - _19277;
    assign _20189 = _20185 ? _20188 : _20183;
    assign _20190 = _20189[62:0];
    assign _20192 = { _20190,
                      _20191 };
    assign _20193 = _20192 < _19277;
    assign _20194 = ~ _20193;
    assign _20182 = _19857[27:27];
    assign _20179 = _20174 - _19277;
    assign _20180 = _20176 ? _20179 : _20174;
    assign _20181 = _20180[62:0];
    assign _20183 = { _20181,
                      _20182 };
    assign _20184 = _20183 < _19277;
    assign _20185 = ~ _20184;
    assign _20173 = _19857[28:28];
    assign _20170 = _20165 - _19277;
    assign _20171 = _20167 ? _20170 : _20165;
    assign _20172 = _20171[62:0];
    assign _20174 = { _20172,
                      _20173 };
    assign _20175 = _20174 < _19277;
    assign _20176 = ~ _20175;
    assign _20164 = _19857[29:29];
    assign _20161 = _20156 - _19277;
    assign _20162 = _20158 ? _20161 : _20156;
    assign _20163 = _20162[62:0];
    assign _20165 = { _20163,
                      _20164 };
    assign _20166 = _20165 < _19277;
    assign _20167 = ~ _20166;
    assign _20155 = _19857[30:30];
    assign _20152 = _20147 - _19277;
    assign _20153 = _20149 ? _20152 : _20147;
    assign _20154 = _20153[62:0];
    assign _20156 = { _20154,
                      _20155 };
    assign _20157 = _20156 < _19277;
    assign _20158 = ~ _20157;
    assign _20146 = _19857[31:31];
    assign _20143 = _20138 - _19277;
    assign _20144 = _20140 ? _20143 : _20138;
    assign _20145 = _20144[62:0];
    assign _20147 = { _20145,
                      _20146 };
    assign _20148 = _20147 < _19277;
    assign _20149 = ~ _20148;
    assign _20137 = _19857[32:32];
    assign _20134 = _20129 - _19277;
    assign _20135 = _20131 ? _20134 : _20129;
    assign _20136 = _20135[62:0];
    assign _20138 = { _20136,
                      _20137 };
    assign _20139 = _20138 < _19277;
    assign _20140 = ~ _20139;
    assign _20128 = _19857[33:33];
    assign _20125 = _20120 - _19277;
    assign _20126 = _20122 ? _20125 : _20120;
    assign _20127 = _20126[62:0];
    assign _20129 = { _20127,
                      _20128 };
    assign _20130 = _20129 < _19277;
    assign _20131 = ~ _20130;
    assign _20119 = _19857[34:34];
    assign _20116 = _20111 - _19277;
    assign _20117 = _20113 ? _20116 : _20111;
    assign _20118 = _20117[62:0];
    assign _20120 = { _20118,
                      _20119 };
    assign _20121 = _20120 < _19277;
    assign _20122 = ~ _20121;
    assign _20110 = _19857[35:35];
    assign _20107 = _20102 - _19277;
    assign _20108 = _20104 ? _20107 : _20102;
    assign _20109 = _20108[62:0];
    assign _20111 = { _20109,
                      _20110 };
    assign _20112 = _20111 < _19277;
    assign _20113 = ~ _20112;
    assign _20101 = _19857[36:36];
    assign _20098 = _20093 - _19277;
    assign _20099 = _20095 ? _20098 : _20093;
    assign _20100 = _20099[62:0];
    assign _20102 = { _20100,
                      _20101 };
    assign _20103 = _20102 < _19277;
    assign _20104 = ~ _20103;
    assign _20092 = _19857[37:37];
    assign _20089 = _20084 - _19277;
    assign _20090 = _20086 ? _20089 : _20084;
    assign _20091 = _20090[62:0];
    assign _20093 = { _20091,
                      _20092 };
    assign _20094 = _20093 < _19277;
    assign _20095 = ~ _20094;
    assign _20083 = _19857[38:38];
    assign _20080 = _20075 - _19277;
    assign _20081 = _20077 ? _20080 : _20075;
    assign _20082 = _20081[62:0];
    assign _20084 = { _20082,
                      _20083 };
    assign _20085 = _20084 < _19277;
    assign _20086 = ~ _20085;
    assign _20074 = _19857[39:39];
    assign _20071 = _20066 - _19277;
    assign _20072 = _20068 ? _20071 : _20066;
    assign _20073 = _20072[62:0];
    assign _20075 = { _20073,
                      _20074 };
    assign _20076 = _20075 < _19277;
    assign _20077 = ~ _20076;
    assign _20065 = _19857[40:40];
    assign _20062 = _20057 - _19277;
    assign _20063 = _20059 ? _20062 : _20057;
    assign _20064 = _20063[62:0];
    assign _20066 = { _20064,
                      _20065 };
    assign _20067 = _20066 < _19277;
    assign _20068 = ~ _20067;
    assign _20056 = _19857[41:41];
    assign _20053 = _20048 - _19277;
    assign _20054 = _20050 ? _20053 : _20048;
    assign _20055 = _20054[62:0];
    assign _20057 = { _20055,
                      _20056 };
    assign _20058 = _20057 < _19277;
    assign _20059 = ~ _20058;
    assign _20047 = _19857[42:42];
    assign _20044 = _20039 - _19277;
    assign _20045 = _20041 ? _20044 : _20039;
    assign _20046 = _20045[62:0];
    assign _20048 = { _20046,
                      _20047 };
    assign _20049 = _20048 < _19277;
    assign _20050 = ~ _20049;
    assign _20038 = _19857[43:43];
    assign _20035 = _20030 - _19277;
    assign _20036 = _20032 ? _20035 : _20030;
    assign _20037 = _20036[62:0];
    assign _20039 = { _20037,
                      _20038 };
    assign _20040 = _20039 < _19277;
    assign _20041 = ~ _20040;
    assign _20029 = _19857[44:44];
    assign _20026 = _20021 - _19277;
    assign _20027 = _20023 ? _20026 : _20021;
    assign _20028 = _20027[62:0];
    assign _20030 = { _20028,
                      _20029 };
    assign _20031 = _20030 < _19277;
    assign _20032 = ~ _20031;
    assign _20020 = _19857[45:45];
    assign _20017 = _20012 - _19277;
    assign _20018 = _20014 ? _20017 : _20012;
    assign _20019 = _20018[62:0];
    assign _20021 = { _20019,
                      _20020 };
    assign _20022 = _20021 < _19277;
    assign _20023 = ~ _20022;
    assign _20011 = _19857[46:46];
    assign _20008 = _20003 - _19277;
    assign _20009 = _20005 ? _20008 : _20003;
    assign _20010 = _20009[62:0];
    assign _20012 = { _20010,
                      _20011 };
    assign _20013 = _20012 < _19277;
    assign _20014 = ~ _20013;
    assign _20002 = _19857[47:47];
    assign _19999 = _19994 - _19277;
    assign _20000 = _19996 ? _19999 : _19994;
    assign _20001 = _20000[62:0];
    assign _20003 = { _20001,
                      _20002 };
    assign _20004 = _20003 < _19277;
    assign _20005 = ~ _20004;
    assign _19993 = _19857[48:48];
    assign _19990 = _19985 - _19277;
    assign _19991 = _19987 ? _19990 : _19985;
    assign _19992 = _19991[62:0];
    assign _19994 = { _19992,
                      _19993 };
    assign _19995 = _19994 < _19277;
    assign _19996 = ~ _19995;
    assign _19984 = _19857[49:49];
    assign _19981 = _19976 - _19277;
    assign _19982 = _19978 ? _19981 : _19976;
    assign _19983 = _19982[62:0];
    assign _19985 = { _19983,
                      _19984 };
    assign _19986 = _19985 < _19277;
    assign _19987 = ~ _19986;
    assign _19975 = _19857[50:50];
    assign _19972 = _19967 - _19277;
    assign _19973 = _19969 ? _19972 : _19967;
    assign _19974 = _19973[62:0];
    assign _19976 = { _19974,
                      _19975 };
    assign _19977 = _19976 < _19277;
    assign _19978 = ~ _19977;
    assign _19966 = _19857[51:51];
    assign _19963 = _19958 - _19277;
    assign _19964 = _19960 ? _19963 : _19958;
    assign _19965 = _19964[62:0];
    assign _19967 = { _19965,
                      _19966 };
    assign _19968 = _19967 < _19277;
    assign _19969 = ~ _19968;
    assign _19957 = _19857[52:52];
    assign _19954 = _19949 - _19277;
    assign _19955 = _19951 ? _19954 : _19949;
    assign _19956 = _19955[62:0];
    assign _19958 = { _19956,
                      _19957 };
    assign _19959 = _19958 < _19277;
    assign _19960 = ~ _19959;
    assign _19948 = _19857[53:53];
    assign _19945 = _19940 - _19277;
    assign _19946 = _19942 ? _19945 : _19940;
    assign _19947 = _19946[62:0];
    assign _19949 = { _19947,
                      _19948 };
    assign _19950 = _19949 < _19277;
    assign _19951 = ~ _19950;
    assign _19939 = _19857[54:54];
    assign _19936 = _19931 - _19277;
    assign _19937 = _19933 ? _19936 : _19931;
    assign _19938 = _19937[62:0];
    assign _19940 = { _19938,
                      _19939 };
    assign _19941 = _19940 < _19277;
    assign _19942 = ~ _19941;
    assign _19930 = _19857[55:55];
    assign _19927 = _19922 - _19277;
    assign _19928 = _19924 ? _19927 : _19922;
    assign _19929 = _19928[62:0];
    assign _19931 = { _19929,
                      _19930 };
    assign _19932 = _19931 < _19277;
    assign _19933 = ~ _19932;
    assign _19921 = _19857[56:56];
    assign _19918 = _19913 - _19277;
    assign _19919 = _19915 ? _19918 : _19913;
    assign _19920 = _19919[62:0];
    assign _19922 = { _19920,
                      _19921 };
    assign _19923 = _19922 < _19277;
    assign _19924 = ~ _19923;
    assign _19912 = _19857[57:57];
    assign _19909 = _19904 - _19277;
    assign _19910 = _19906 ? _19909 : _19904;
    assign _19911 = _19910[62:0];
    assign _19913 = { _19911,
                      _19912 };
    assign _19914 = _19913 < _19277;
    assign _19915 = ~ _19914;
    assign _19903 = _19857[58:58];
    assign _19900 = _19895 - _19277;
    assign _19901 = _19897 ? _19900 : _19895;
    assign _19902 = _19901[62:0];
    assign _19904 = { _19902,
                      _19903 };
    assign _19905 = _19904 < _19277;
    assign _19906 = ~ _19905;
    assign _19894 = _19857[59:59];
    assign _19891 = _19886 - _19277;
    assign _19892 = _19888 ? _19891 : _19886;
    assign _19893 = _19892[62:0];
    assign _19895 = { _19893,
                      _19894 };
    assign _19896 = _19895 < _19277;
    assign _19897 = ~ _19896;
    assign _19885 = _19857[60:60];
    assign _19882 = _19877 - _19277;
    assign _19883 = _19879 ? _19882 : _19877;
    assign _19884 = _19883[62:0];
    assign _19886 = { _19884,
                      _19885 };
    assign _19887 = _19886 < _19277;
    assign _19888 = ~ _19887;
    assign _19876 = _19857[61:61];
    assign _19873 = _19868 - _19277;
    assign _19874 = _19870 ? _19873 : _19868;
    assign _19875 = _19874[62:0];
    assign _19877 = { _19875,
                      _19876 };
    assign _19878 = _19877 < _19277;
    assign _19879 = ~ _19878;
    assign _19867 = _19857[62:62];
    assign _19864 = _19859 - _19277;
    assign _19865 = _19861 ? _19864 : _19859;
    assign _19866 = _19865[62:0];
    assign _19868 = { _19866,
                      _19867 };
    assign _19869 = _19868 < _19277;
    assign _19870 = ~ _19869;
    assign _19857 = _19269 - _19851;
    assign _19858 = _19857[63:63];
    assign _19859 = { _22185,
                      _19858 };
    assign _19860 = _19859 < _19277;
    assign _19861 = ~ _19860;
    assign _19862 = { _22185,
                      _19861 };
    assign _19863 = _19862[62:0];
    assign _19871 = { _19863,
                      _19870 };
    assign _19872 = _19871[62:0];
    assign _19880 = { _19872,
                      _19879 };
    assign _19881 = _19880[62:0];
    assign _19889 = { _19881,
                      _19888 };
    assign _19890 = _19889[62:0];
    assign _19898 = { _19890,
                      _19897 };
    assign _19899 = _19898[62:0];
    assign _19907 = { _19899,
                      _19906 };
    assign _19908 = _19907[62:0];
    assign _19916 = { _19908,
                      _19915 };
    assign _19917 = _19916[62:0];
    assign _19925 = { _19917,
                      _19924 };
    assign _19926 = _19925[62:0];
    assign _19934 = { _19926,
                      _19933 };
    assign _19935 = _19934[62:0];
    assign _19943 = { _19935,
                      _19942 };
    assign _19944 = _19943[62:0];
    assign _19952 = { _19944,
                      _19951 };
    assign _19953 = _19952[62:0];
    assign _19961 = { _19953,
                      _19960 };
    assign _19962 = _19961[62:0];
    assign _19970 = { _19962,
                      _19969 };
    assign _19971 = _19970[62:0];
    assign _19979 = { _19971,
                      _19978 };
    assign _19980 = _19979[62:0];
    assign _19988 = { _19980,
                      _19987 };
    assign _19989 = _19988[62:0];
    assign _19997 = { _19989,
                      _19996 };
    assign _19998 = _19997[62:0];
    assign _20006 = { _19998,
                      _20005 };
    assign _20007 = _20006[62:0];
    assign _20015 = { _20007,
                      _20014 };
    assign _20016 = _20015[62:0];
    assign _20024 = { _20016,
                      _20023 };
    assign _20025 = _20024[62:0];
    assign _20033 = { _20025,
                      _20032 };
    assign _20034 = _20033[62:0];
    assign _20042 = { _20034,
                      _20041 };
    assign _20043 = _20042[62:0];
    assign _20051 = { _20043,
                      _20050 };
    assign _20052 = _20051[62:0];
    assign _20060 = { _20052,
                      _20059 };
    assign _20061 = _20060[62:0];
    assign _20069 = { _20061,
                      _20068 };
    assign _20070 = _20069[62:0];
    assign _20078 = { _20070,
                      _20077 };
    assign _20079 = _20078[62:0];
    assign _20087 = { _20079,
                      _20086 };
    assign _20088 = _20087[62:0];
    assign _20096 = { _20088,
                      _20095 };
    assign _20097 = _20096[62:0];
    assign _20105 = { _20097,
                      _20104 };
    assign _20106 = _20105[62:0];
    assign _20114 = { _20106,
                      _20113 };
    assign _20115 = _20114[62:0];
    assign _20123 = { _20115,
                      _20122 };
    assign _20124 = _20123[62:0];
    assign _20132 = { _20124,
                      _20131 };
    assign _20133 = _20132[62:0];
    assign _20141 = { _20133,
                      _20140 };
    assign _20142 = _20141[62:0];
    assign _20150 = { _20142,
                      _20149 };
    assign _20151 = _20150[62:0];
    assign _20159 = { _20151,
                      _20158 };
    assign _20160 = _20159[62:0];
    assign _20168 = { _20160,
                      _20167 };
    assign _20169 = _20168[62:0];
    assign _20177 = { _20169,
                      _20176 };
    assign _20178 = _20177[62:0];
    assign _20186 = { _20178,
                      _20185 };
    assign _20187 = _20186[62:0];
    assign _20195 = { _20187,
                      _20194 };
    assign _20196 = _20195[62:0];
    assign _20204 = { _20196,
                      _20203 };
    assign _20205 = _20204[62:0];
    assign _20213 = { _20205,
                      _20212 };
    assign _20214 = _20213[62:0];
    assign _20222 = { _20214,
                      _20221 };
    assign _20223 = _20222[62:0];
    assign _20231 = { _20223,
                      _20230 };
    assign _20232 = _20231[62:0];
    assign _20240 = { _20232,
                      _20239 };
    assign _20241 = _20240[62:0];
    assign _20249 = { _20241,
                      _20248 };
    assign _20250 = _20249[62:0];
    assign _20258 = { _20250,
                      _20257 };
    assign _20259 = _20258[62:0];
    assign _20267 = { _20259,
                      _20266 };
    assign _20268 = _20267[62:0];
    assign _20276 = { _20268,
                      _20275 };
    assign _20277 = _20276[62:0];
    assign _20285 = { _20277,
                      _20284 };
    assign _20286 = _20285[62:0];
    assign _20294 = { _20286,
                      _20293 };
    assign _20295 = _20294[62:0];
    assign _20303 = { _20295,
                      _20302 };
    assign _20304 = _20303[62:0];
    assign _20312 = { _20304,
                      _20311 };
    assign _20313 = _20312[62:0];
    assign _20321 = { _20313,
                      _20320 };
    assign _20322 = _20321[62:0];
    assign _20330 = { _20322,
                      _20329 };
    assign _20331 = _20330[62:0];
    assign _20339 = { _20331,
                      _20338 };
    assign _20340 = _20339[62:0];
    assign _20348 = { _20340,
                      _20347 };
    assign _20349 = _20348[62:0];
    assign _20357 = { _20349,
                      _20356 };
    assign _20358 = _20357[62:0];
    assign _20366 = { _20358,
                      _20365 };
    assign _20367 = _20366[62:0];
    assign _20375 = { _20367,
                      _20374 };
    assign _20376 = _20375[62:0];
    assign _20384 = { _20376,
                      _20383 };
    assign _20385 = _20384[62:0];
    assign _20393 = { _20385,
                      _20392 };
    assign _20394 = _20393[62:0];
    assign _20402 = { _20394,
                      _20401 };
    assign _20403 = _20402[62:0];
    assign _20411 = { _20403,
                      _20410 };
    assign _20412 = _20411[62:0];
    assign _20420 = { _20412,
                      _20419 };
    assign _20421 = _20420[62:0];
    assign _20429 = { _20421,
                      _20428 };
    assign _20431 = _20429 + _22186;
    assign _20432 = _20431 * _19851;
    assign _20433 = _20432[63:0];
    assign _21015 = _20433 + _21014;
    assign _19843 = _19274[0:0];
    assign _19840 = _19835 - _19277;
    assign _19841 = _19837 ? _19840 : _19835;
    assign _19842 = _19841[62:0];
    assign _19844 = { _19842,
                      _19843 };
    assign _19845 = _19844 < _19277;
    assign _19846 = ~ _19845;
    assign _19834 = _19274[1:1];
    assign _19831 = _19826 - _19277;
    assign _19832 = _19828 ? _19831 : _19826;
    assign _19833 = _19832[62:0];
    assign _19835 = { _19833,
                      _19834 };
    assign _19836 = _19835 < _19277;
    assign _19837 = ~ _19836;
    assign _19825 = _19274[2:2];
    assign _19822 = _19817 - _19277;
    assign _19823 = _19819 ? _19822 : _19817;
    assign _19824 = _19823[62:0];
    assign _19826 = { _19824,
                      _19825 };
    assign _19827 = _19826 < _19277;
    assign _19828 = ~ _19827;
    assign _19816 = _19274[3:3];
    assign _19813 = _19808 - _19277;
    assign _19814 = _19810 ? _19813 : _19808;
    assign _19815 = _19814[62:0];
    assign _19817 = { _19815,
                      _19816 };
    assign _19818 = _19817 < _19277;
    assign _19819 = ~ _19818;
    assign _19807 = _19274[4:4];
    assign _19804 = _19799 - _19277;
    assign _19805 = _19801 ? _19804 : _19799;
    assign _19806 = _19805[62:0];
    assign _19808 = { _19806,
                      _19807 };
    assign _19809 = _19808 < _19277;
    assign _19810 = ~ _19809;
    assign _19798 = _19274[5:5];
    assign _19795 = _19790 - _19277;
    assign _19796 = _19792 ? _19795 : _19790;
    assign _19797 = _19796[62:0];
    assign _19799 = { _19797,
                      _19798 };
    assign _19800 = _19799 < _19277;
    assign _19801 = ~ _19800;
    assign _19789 = _19274[6:6];
    assign _19786 = _19781 - _19277;
    assign _19787 = _19783 ? _19786 : _19781;
    assign _19788 = _19787[62:0];
    assign _19790 = { _19788,
                      _19789 };
    assign _19791 = _19790 < _19277;
    assign _19792 = ~ _19791;
    assign _19780 = _19274[7:7];
    assign _19777 = _19772 - _19277;
    assign _19778 = _19774 ? _19777 : _19772;
    assign _19779 = _19778[62:0];
    assign _19781 = { _19779,
                      _19780 };
    assign _19782 = _19781 < _19277;
    assign _19783 = ~ _19782;
    assign _19771 = _19274[8:8];
    assign _19768 = _19763 - _19277;
    assign _19769 = _19765 ? _19768 : _19763;
    assign _19770 = _19769[62:0];
    assign _19772 = { _19770,
                      _19771 };
    assign _19773 = _19772 < _19277;
    assign _19774 = ~ _19773;
    assign _19762 = _19274[9:9];
    assign _19759 = _19754 - _19277;
    assign _19760 = _19756 ? _19759 : _19754;
    assign _19761 = _19760[62:0];
    assign _19763 = { _19761,
                      _19762 };
    assign _19764 = _19763 < _19277;
    assign _19765 = ~ _19764;
    assign _19753 = _19274[10:10];
    assign _19750 = _19745 - _19277;
    assign _19751 = _19747 ? _19750 : _19745;
    assign _19752 = _19751[62:0];
    assign _19754 = { _19752,
                      _19753 };
    assign _19755 = _19754 < _19277;
    assign _19756 = ~ _19755;
    assign _19744 = _19274[11:11];
    assign _19741 = _19736 - _19277;
    assign _19742 = _19738 ? _19741 : _19736;
    assign _19743 = _19742[62:0];
    assign _19745 = { _19743,
                      _19744 };
    assign _19746 = _19745 < _19277;
    assign _19747 = ~ _19746;
    assign _19735 = _19274[12:12];
    assign _19732 = _19727 - _19277;
    assign _19733 = _19729 ? _19732 : _19727;
    assign _19734 = _19733[62:0];
    assign _19736 = { _19734,
                      _19735 };
    assign _19737 = _19736 < _19277;
    assign _19738 = ~ _19737;
    assign _19726 = _19274[13:13];
    assign _19723 = _19718 - _19277;
    assign _19724 = _19720 ? _19723 : _19718;
    assign _19725 = _19724[62:0];
    assign _19727 = { _19725,
                      _19726 };
    assign _19728 = _19727 < _19277;
    assign _19729 = ~ _19728;
    assign _19717 = _19274[14:14];
    assign _19714 = _19709 - _19277;
    assign _19715 = _19711 ? _19714 : _19709;
    assign _19716 = _19715[62:0];
    assign _19718 = { _19716,
                      _19717 };
    assign _19719 = _19718 < _19277;
    assign _19720 = ~ _19719;
    assign _19708 = _19274[15:15];
    assign _19705 = _19700 - _19277;
    assign _19706 = _19702 ? _19705 : _19700;
    assign _19707 = _19706[62:0];
    assign _19709 = { _19707,
                      _19708 };
    assign _19710 = _19709 < _19277;
    assign _19711 = ~ _19710;
    assign _19699 = _19274[16:16];
    assign _19696 = _19691 - _19277;
    assign _19697 = _19693 ? _19696 : _19691;
    assign _19698 = _19697[62:0];
    assign _19700 = { _19698,
                      _19699 };
    assign _19701 = _19700 < _19277;
    assign _19702 = ~ _19701;
    assign _19690 = _19274[17:17];
    assign _19687 = _19682 - _19277;
    assign _19688 = _19684 ? _19687 : _19682;
    assign _19689 = _19688[62:0];
    assign _19691 = { _19689,
                      _19690 };
    assign _19692 = _19691 < _19277;
    assign _19693 = ~ _19692;
    assign _19681 = _19274[18:18];
    assign _19678 = _19673 - _19277;
    assign _19679 = _19675 ? _19678 : _19673;
    assign _19680 = _19679[62:0];
    assign _19682 = { _19680,
                      _19681 };
    assign _19683 = _19682 < _19277;
    assign _19684 = ~ _19683;
    assign _19672 = _19274[19:19];
    assign _19669 = _19664 - _19277;
    assign _19670 = _19666 ? _19669 : _19664;
    assign _19671 = _19670[62:0];
    assign _19673 = { _19671,
                      _19672 };
    assign _19674 = _19673 < _19277;
    assign _19675 = ~ _19674;
    assign _19663 = _19274[20:20];
    assign _19660 = _19655 - _19277;
    assign _19661 = _19657 ? _19660 : _19655;
    assign _19662 = _19661[62:0];
    assign _19664 = { _19662,
                      _19663 };
    assign _19665 = _19664 < _19277;
    assign _19666 = ~ _19665;
    assign _19654 = _19274[21:21];
    assign _19651 = _19646 - _19277;
    assign _19652 = _19648 ? _19651 : _19646;
    assign _19653 = _19652[62:0];
    assign _19655 = { _19653,
                      _19654 };
    assign _19656 = _19655 < _19277;
    assign _19657 = ~ _19656;
    assign _19645 = _19274[22:22];
    assign _19642 = _19637 - _19277;
    assign _19643 = _19639 ? _19642 : _19637;
    assign _19644 = _19643[62:0];
    assign _19646 = { _19644,
                      _19645 };
    assign _19647 = _19646 < _19277;
    assign _19648 = ~ _19647;
    assign _19636 = _19274[23:23];
    assign _19633 = _19628 - _19277;
    assign _19634 = _19630 ? _19633 : _19628;
    assign _19635 = _19634[62:0];
    assign _19637 = { _19635,
                      _19636 };
    assign _19638 = _19637 < _19277;
    assign _19639 = ~ _19638;
    assign _19627 = _19274[24:24];
    assign _19624 = _19619 - _19277;
    assign _19625 = _19621 ? _19624 : _19619;
    assign _19626 = _19625[62:0];
    assign _19628 = { _19626,
                      _19627 };
    assign _19629 = _19628 < _19277;
    assign _19630 = ~ _19629;
    assign _19618 = _19274[25:25];
    assign _19615 = _19610 - _19277;
    assign _19616 = _19612 ? _19615 : _19610;
    assign _19617 = _19616[62:0];
    assign _19619 = { _19617,
                      _19618 };
    assign _19620 = _19619 < _19277;
    assign _19621 = ~ _19620;
    assign _19609 = _19274[26:26];
    assign _19606 = _19601 - _19277;
    assign _19607 = _19603 ? _19606 : _19601;
    assign _19608 = _19607[62:0];
    assign _19610 = { _19608,
                      _19609 };
    assign _19611 = _19610 < _19277;
    assign _19612 = ~ _19611;
    assign _19600 = _19274[27:27];
    assign _19597 = _19592 - _19277;
    assign _19598 = _19594 ? _19597 : _19592;
    assign _19599 = _19598[62:0];
    assign _19601 = { _19599,
                      _19600 };
    assign _19602 = _19601 < _19277;
    assign _19603 = ~ _19602;
    assign _19591 = _19274[28:28];
    assign _19588 = _19583 - _19277;
    assign _19589 = _19585 ? _19588 : _19583;
    assign _19590 = _19589[62:0];
    assign _19592 = { _19590,
                      _19591 };
    assign _19593 = _19592 < _19277;
    assign _19594 = ~ _19593;
    assign _19582 = _19274[29:29];
    assign _19579 = _19574 - _19277;
    assign _19580 = _19576 ? _19579 : _19574;
    assign _19581 = _19580[62:0];
    assign _19583 = { _19581,
                      _19582 };
    assign _19584 = _19583 < _19277;
    assign _19585 = ~ _19584;
    assign _19573 = _19274[30:30];
    assign _19570 = _19565 - _19277;
    assign _19571 = _19567 ? _19570 : _19565;
    assign _19572 = _19571[62:0];
    assign _19574 = { _19572,
                      _19573 };
    assign _19575 = _19574 < _19277;
    assign _19576 = ~ _19575;
    assign _19564 = _19274[31:31];
    assign _19561 = _19556 - _19277;
    assign _19562 = _19558 ? _19561 : _19556;
    assign _19563 = _19562[62:0];
    assign _19565 = { _19563,
                      _19564 };
    assign _19566 = _19565 < _19277;
    assign _19567 = ~ _19566;
    assign _19555 = _19274[32:32];
    assign _19552 = _19547 - _19277;
    assign _19553 = _19549 ? _19552 : _19547;
    assign _19554 = _19553[62:0];
    assign _19556 = { _19554,
                      _19555 };
    assign _19557 = _19556 < _19277;
    assign _19558 = ~ _19557;
    assign _19546 = _19274[33:33];
    assign _19543 = _19538 - _19277;
    assign _19544 = _19540 ? _19543 : _19538;
    assign _19545 = _19544[62:0];
    assign _19547 = { _19545,
                      _19546 };
    assign _19548 = _19547 < _19277;
    assign _19549 = ~ _19548;
    assign _19537 = _19274[34:34];
    assign _19534 = _19529 - _19277;
    assign _19535 = _19531 ? _19534 : _19529;
    assign _19536 = _19535[62:0];
    assign _19538 = { _19536,
                      _19537 };
    assign _19539 = _19538 < _19277;
    assign _19540 = ~ _19539;
    assign _19528 = _19274[35:35];
    assign _19525 = _19520 - _19277;
    assign _19526 = _19522 ? _19525 : _19520;
    assign _19527 = _19526[62:0];
    assign _19529 = { _19527,
                      _19528 };
    assign _19530 = _19529 < _19277;
    assign _19531 = ~ _19530;
    assign _19519 = _19274[36:36];
    assign _19516 = _19511 - _19277;
    assign _19517 = _19513 ? _19516 : _19511;
    assign _19518 = _19517[62:0];
    assign _19520 = { _19518,
                      _19519 };
    assign _19521 = _19520 < _19277;
    assign _19522 = ~ _19521;
    assign _19510 = _19274[37:37];
    assign _19507 = _19502 - _19277;
    assign _19508 = _19504 ? _19507 : _19502;
    assign _19509 = _19508[62:0];
    assign _19511 = { _19509,
                      _19510 };
    assign _19512 = _19511 < _19277;
    assign _19513 = ~ _19512;
    assign _19501 = _19274[38:38];
    assign _19498 = _19493 - _19277;
    assign _19499 = _19495 ? _19498 : _19493;
    assign _19500 = _19499[62:0];
    assign _19502 = { _19500,
                      _19501 };
    assign _19503 = _19502 < _19277;
    assign _19504 = ~ _19503;
    assign _19492 = _19274[39:39];
    assign _19489 = _19484 - _19277;
    assign _19490 = _19486 ? _19489 : _19484;
    assign _19491 = _19490[62:0];
    assign _19493 = { _19491,
                      _19492 };
    assign _19494 = _19493 < _19277;
    assign _19495 = ~ _19494;
    assign _19483 = _19274[40:40];
    assign _19480 = _19475 - _19277;
    assign _19481 = _19477 ? _19480 : _19475;
    assign _19482 = _19481[62:0];
    assign _19484 = { _19482,
                      _19483 };
    assign _19485 = _19484 < _19277;
    assign _19486 = ~ _19485;
    assign _19474 = _19274[41:41];
    assign _19471 = _19466 - _19277;
    assign _19472 = _19468 ? _19471 : _19466;
    assign _19473 = _19472[62:0];
    assign _19475 = { _19473,
                      _19474 };
    assign _19476 = _19475 < _19277;
    assign _19477 = ~ _19476;
    assign _19465 = _19274[42:42];
    assign _19462 = _19457 - _19277;
    assign _19463 = _19459 ? _19462 : _19457;
    assign _19464 = _19463[62:0];
    assign _19466 = { _19464,
                      _19465 };
    assign _19467 = _19466 < _19277;
    assign _19468 = ~ _19467;
    assign _19456 = _19274[43:43];
    assign _19453 = _19448 - _19277;
    assign _19454 = _19450 ? _19453 : _19448;
    assign _19455 = _19454[62:0];
    assign _19457 = { _19455,
                      _19456 };
    assign _19458 = _19457 < _19277;
    assign _19459 = ~ _19458;
    assign _19447 = _19274[44:44];
    assign _19444 = _19439 - _19277;
    assign _19445 = _19441 ? _19444 : _19439;
    assign _19446 = _19445[62:0];
    assign _19448 = { _19446,
                      _19447 };
    assign _19449 = _19448 < _19277;
    assign _19450 = ~ _19449;
    assign _19438 = _19274[45:45];
    assign _19435 = _19430 - _19277;
    assign _19436 = _19432 ? _19435 : _19430;
    assign _19437 = _19436[62:0];
    assign _19439 = { _19437,
                      _19438 };
    assign _19440 = _19439 < _19277;
    assign _19441 = ~ _19440;
    assign _19429 = _19274[46:46];
    assign _19426 = _19421 - _19277;
    assign _19427 = _19423 ? _19426 : _19421;
    assign _19428 = _19427[62:0];
    assign _19430 = { _19428,
                      _19429 };
    assign _19431 = _19430 < _19277;
    assign _19432 = ~ _19431;
    assign _19420 = _19274[47:47];
    assign _19417 = _19412 - _19277;
    assign _19418 = _19414 ? _19417 : _19412;
    assign _19419 = _19418[62:0];
    assign _19421 = { _19419,
                      _19420 };
    assign _19422 = _19421 < _19277;
    assign _19423 = ~ _19422;
    assign _19411 = _19274[48:48];
    assign _19408 = _19403 - _19277;
    assign _19409 = _19405 ? _19408 : _19403;
    assign _19410 = _19409[62:0];
    assign _19412 = { _19410,
                      _19411 };
    assign _19413 = _19412 < _19277;
    assign _19414 = ~ _19413;
    assign _19402 = _19274[49:49];
    assign _19399 = _19394 - _19277;
    assign _19400 = _19396 ? _19399 : _19394;
    assign _19401 = _19400[62:0];
    assign _19403 = { _19401,
                      _19402 };
    assign _19404 = _19403 < _19277;
    assign _19405 = ~ _19404;
    assign _19393 = _19274[50:50];
    assign _19390 = _19385 - _19277;
    assign _19391 = _19387 ? _19390 : _19385;
    assign _19392 = _19391[62:0];
    assign _19394 = { _19392,
                      _19393 };
    assign _19395 = _19394 < _19277;
    assign _19396 = ~ _19395;
    assign _19384 = _19274[51:51];
    assign _19381 = _19376 - _19277;
    assign _19382 = _19378 ? _19381 : _19376;
    assign _19383 = _19382[62:0];
    assign _19385 = { _19383,
                      _19384 };
    assign _19386 = _19385 < _19277;
    assign _19387 = ~ _19386;
    assign _19375 = _19274[52:52];
    assign _19372 = _19367 - _19277;
    assign _19373 = _19369 ? _19372 : _19367;
    assign _19374 = _19373[62:0];
    assign _19376 = { _19374,
                      _19375 };
    assign _19377 = _19376 < _19277;
    assign _19378 = ~ _19377;
    assign _19366 = _19274[53:53];
    assign _19363 = _19358 - _19277;
    assign _19364 = _19360 ? _19363 : _19358;
    assign _19365 = _19364[62:0];
    assign _19367 = { _19365,
                      _19366 };
    assign _19368 = _19367 < _19277;
    assign _19369 = ~ _19368;
    assign _19357 = _19274[54:54];
    assign _19354 = _19349 - _19277;
    assign _19355 = _19351 ? _19354 : _19349;
    assign _19356 = _19355[62:0];
    assign _19358 = { _19356,
                      _19357 };
    assign _19359 = _19358 < _19277;
    assign _19360 = ~ _19359;
    assign _19348 = _19274[55:55];
    assign _19345 = _19340 - _19277;
    assign _19346 = _19342 ? _19345 : _19340;
    assign _19347 = _19346[62:0];
    assign _19349 = { _19347,
                      _19348 };
    assign _19350 = _19349 < _19277;
    assign _19351 = ~ _19350;
    assign _19339 = _19274[56:56];
    assign _19336 = _19331 - _19277;
    assign _19337 = _19333 ? _19336 : _19331;
    assign _19338 = _19337[62:0];
    assign _19340 = { _19338,
                      _19339 };
    assign _19341 = _19340 < _19277;
    assign _19342 = ~ _19341;
    assign _19330 = _19274[57:57];
    assign _19327 = _19322 - _19277;
    assign _19328 = _19324 ? _19327 : _19322;
    assign _19329 = _19328[62:0];
    assign _19331 = { _19329,
                      _19330 };
    assign _19332 = _19331 < _19277;
    assign _19333 = ~ _19332;
    assign _19321 = _19274[58:58];
    assign _19318 = _19313 - _19277;
    assign _19319 = _19315 ? _19318 : _19313;
    assign _19320 = _19319[62:0];
    assign _19322 = { _19320,
                      _19321 };
    assign _19323 = _19322 < _19277;
    assign _19324 = ~ _19323;
    assign _19312 = _19274[59:59];
    assign _19309 = _19304 - _19277;
    assign _19310 = _19306 ? _19309 : _19304;
    assign _19311 = _19310[62:0];
    assign _19313 = { _19311,
                      _19312 };
    assign _19314 = _19313 < _19277;
    assign _19315 = ~ _19314;
    assign _19303 = _19274[60:60];
    assign _19300 = _19295 - _19277;
    assign _19301 = _19297 ? _19300 : _19295;
    assign _19302 = _19301[62:0];
    assign _19304 = { _19302,
                      _19303 };
    assign _19305 = _19304 < _19277;
    assign _19306 = ~ _19305;
    assign _19294 = _19274[61:61];
    assign _19291 = _19286 - _19277;
    assign _19292 = _19288 ? _19291 : _19286;
    assign _19293 = _19292[62:0];
    assign _19295 = { _19293,
                      _19294 };
    assign _19296 = _19295 < _19277;
    assign _19297 = ~ _19296;
    assign _19285 = _19274[62:62];
    assign _19282 = _19276 - _19277;
    assign _19283 = _19279 ? _19282 : _19276;
    assign _19284 = _19283[62:0];
    assign _19286 = { _19284,
                      _19285 };
    assign _19287 = _19286 < _19277;
    assign _19288 = ~ _19287;
    assign _19277 = 64'b0000000000000000000000000000000000000000000000011011001000000111;
    assign _19273 = 64'b0000000000000000000000000000000000000000000000011011001000000110;
    assign _19274 = _3 + _19273;
    assign _19275 = _19274[63:63];
    assign _19276 = { _22185,
                      _19275 };
    assign _19278 = _19276 < _19277;
    assign _19279 = ~ _19278;
    assign _19280 = { _22185,
                      _19279 };
    assign _19281 = _19280[62:0];
    assign _19289 = { _19281,
                      _19288 };
    assign _19290 = _19289[62:0];
    assign _19298 = { _19290,
                      _19297 };
    assign _19299 = _19298[62:0];
    assign _19307 = { _19299,
                      _19306 };
    assign _19308 = _19307[62:0];
    assign _19316 = { _19308,
                      _19315 };
    assign _19317 = _19316[62:0];
    assign _19325 = { _19317,
                      _19324 };
    assign _19326 = _19325[62:0];
    assign _19334 = { _19326,
                      _19333 };
    assign _19335 = _19334[62:0];
    assign _19343 = { _19335,
                      _19342 };
    assign _19344 = _19343[62:0];
    assign _19352 = { _19344,
                      _19351 };
    assign _19353 = _19352[62:0];
    assign _19361 = { _19353,
                      _19360 };
    assign _19362 = _19361[62:0];
    assign _19370 = { _19362,
                      _19369 };
    assign _19371 = _19370[62:0];
    assign _19379 = { _19371,
                      _19378 };
    assign _19380 = _19379[62:0];
    assign _19388 = { _19380,
                      _19387 };
    assign _19389 = _19388[62:0];
    assign _19397 = { _19389,
                      _19396 };
    assign _19398 = _19397[62:0];
    assign _19406 = { _19398,
                      _19405 };
    assign _19407 = _19406[62:0];
    assign _19415 = { _19407,
                      _19414 };
    assign _19416 = _19415[62:0];
    assign _19424 = { _19416,
                      _19423 };
    assign _19425 = _19424[62:0];
    assign _19433 = { _19425,
                      _19432 };
    assign _19434 = _19433[62:0];
    assign _19442 = { _19434,
                      _19441 };
    assign _19443 = _19442[62:0];
    assign _19451 = { _19443,
                      _19450 };
    assign _19452 = _19451[62:0];
    assign _19460 = { _19452,
                      _19459 };
    assign _19461 = _19460[62:0];
    assign _19469 = { _19461,
                      _19468 };
    assign _19470 = _19469[62:0];
    assign _19478 = { _19470,
                      _19477 };
    assign _19479 = _19478[62:0];
    assign _19487 = { _19479,
                      _19486 };
    assign _19488 = _19487[62:0];
    assign _19496 = { _19488,
                      _19495 };
    assign _19497 = _19496[62:0];
    assign _19505 = { _19497,
                      _19504 };
    assign _19506 = _19505[62:0];
    assign _19514 = { _19506,
                      _19513 };
    assign _19515 = _19514[62:0];
    assign _19523 = { _19515,
                      _19522 };
    assign _19524 = _19523[62:0];
    assign _19532 = { _19524,
                      _19531 };
    assign _19533 = _19532[62:0];
    assign _19541 = { _19533,
                      _19540 };
    assign _19542 = _19541[62:0];
    assign _19550 = { _19542,
                      _19549 };
    assign _19551 = _19550[62:0];
    assign _19559 = { _19551,
                      _19558 };
    assign _19560 = _19559[62:0];
    assign _19568 = { _19560,
                      _19567 };
    assign _19569 = _19568[62:0];
    assign _19577 = { _19569,
                      _19576 };
    assign _19578 = _19577[62:0];
    assign _19586 = { _19578,
                      _19585 };
    assign _19587 = _19586[62:0];
    assign _19595 = { _19587,
                      _19594 };
    assign _19596 = _19595[62:0];
    assign _19604 = { _19596,
                      _19603 };
    assign _19605 = _19604[62:0];
    assign _19613 = { _19605,
                      _19612 };
    assign _19614 = _19613[62:0];
    assign _19622 = { _19614,
                      _19621 };
    assign _19623 = _19622[62:0];
    assign _19631 = { _19623,
                      _19630 };
    assign _19632 = _19631[62:0];
    assign _19640 = { _19632,
                      _19639 };
    assign _19641 = _19640[62:0];
    assign _19649 = { _19641,
                      _19648 };
    assign _19650 = _19649[62:0];
    assign _19658 = { _19650,
                      _19657 };
    assign _19659 = _19658[62:0];
    assign _19667 = { _19659,
                      _19666 };
    assign _19668 = _19667[62:0];
    assign _19676 = { _19668,
                      _19675 };
    assign _19677 = _19676[62:0];
    assign _19685 = { _19677,
                      _19684 };
    assign _19686 = _19685[62:0];
    assign _19694 = { _19686,
                      _19693 };
    assign _19695 = _19694[62:0];
    assign _19703 = { _19695,
                      _19702 };
    assign _19704 = _19703[62:0];
    assign _19712 = { _19704,
                      _19711 };
    assign _19713 = _19712[62:0];
    assign _19721 = { _19713,
                      _19720 };
    assign _19722 = _19721[62:0];
    assign _19730 = { _19722,
                      _19729 };
    assign _19731 = _19730[62:0];
    assign _19739 = { _19731,
                      _19738 };
    assign _19740 = _19739[62:0];
    assign _19748 = { _19740,
                      _19747 };
    assign _19749 = _19748[62:0];
    assign _19757 = { _19749,
                      _19756 };
    assign _19758 = _19757[62:0];
    assign _19766 = { _19758,
                      _19765 };
    assign _19767 = _19766[62:0];
    assign _19775 = { _19767,
                      _19774 };
    assign _19776 = _19775[62:0];
    assign _19784 = { _19776,
                      _19783 };
    assign _19785 = _19784[62:0];
    assign _19793 = { _19785,
                      _19792 };
    assign _19794 = _19793[62:0];
    assign _19802 = { _19794,
                      _19801 };
    assign _19803 = _19802[62:0];
    assign _19811 = { _19803,
                      _19810 };
    assign _19812 = _19811[62:0];
    assign _19820 = { _19812,
                      _19819 };
    assign _19821 = _19820[62:0];
    assign _19829 = { _19821,
                      _19828 };
    assign _19830 = _19829[62:0];
    assign _19838 = { _19830,
                      _19837 };
    assign _19839 = _19838[62:0];
    assign _19847 = { _19839,
                      _19846 };
    assign _19848 = _19847 * _19277;
    assign _19849 = _19848[63:0];
    assign _19850 = _19277 < _19849;
    assign _19851 = _19850 ? _19849 : _19277;
    assign _19267 = 64'b0000000000000000000000000000000000000000000011110100001000111111;
    assign _19268 = _5 < _19267;
    assign _19269 = _19268 ? _5 : _19267;
    assign _19852 = _19269 < _19851;
    assign _19853 = ~ _19852;
    assign _21016 = _19853 ? _21015 : _21604;
    assign _22767 = _21016 + _22766;
    assign _19256 = _18687[0:0];
    assign _19253 = _19248 - _22192;
    assign _19254 = _19250 ? _19253 : _19248;
    assign _19255 = _19254[62:0];
    assign _19257 = { _19255,
                      _19256 };
    assign _19258 = _19257 < _22192;
    assign _19259 = ~ _19258;
    assign _19247 = _18687[1:1];
    assign _19244 = _19239 - _22192;
    assign _19245 = _19241 ? _19244 : _19239;
    assign _19246 = _19245[62:0];
    assign _19248 = { _19246,
                      _19247 };
    assign _19249 = _19248 < _22192;
    assign _19250 = ~ _19249;
    assign _19238 = _18687[2:2];
    assign _19235 = _19230 - _22192;
    assign _19236 = _19232 ? _19235 : _19230;
    assign _19237 = _19236[62:0];
    assign _19239 = { _19237,
                      _19238 };
    assign _19240 = _19239 < _22192;
    assign _19241 = ~ _19240;
    assign _19229 = _18687[3:3];
    assign _19226 = _19221 - _22192;
    assign _19227 = _19223 ? _19226 : _19221;
    assign _19228 = _19227[62:0];
    assign _19230 = { _19228,
                      _19229 };
    assign _19231 = _19230 < _22192;
    assign _19232 = ~ _19231;
    assign _19220 = _18687[4:4];
    assign _19217 = _19212 - _22192;
    assign _19218 = _19214 ? _19217 : _19212;
    assign _19219 = _19218[62:0];
    assign _19221 = { _19219,
                      _19220 };
    assign _19222 = _19221 < _22192;
    assign _19223 = ~ _19222;
    assign _19211 = _18687[5:5];
    assign _19208 = _19203 - _22192;
    assign _19209 = _19205 ? _19208 : _19203;
    assign _19210 = _19209[62:0];
    assign _19212 = { _19210,
                      _19211 };
    assign _19213 = _19212 < _22192;
    assign _19214 = ~ _19213;
    assign _19202 = _18687[6:6];
    assign _19199 = _19194 - _22192;
    assign _19200 = _19196 ? _19199 : _19194;
    assign _19201 = _19200[62:0];
    assign _19203 = { _19201,
                      _19202 };
    assign _19204 = _19203 < _22192;
    assign _19205 = ~ _19204;
    assign _19193 = _18687[7:7];
    assign _19190 = _19185 - _22192;
    assign _19191 = _19187 ? _19190 : _19185;
    assign _19192 = _19191[62:0];
    assign _19194 = { _19192,
                      _19193 };
    assign _19195 = _19194 < _22192;
    assign _19196 = ~ _19195;
    assign _19184 = _18687[8:8];
    assign _19181 = _19176 - _22192;
    assign _19182 = _19178 ? _19181 : _19176;
    assign _19183 = _19182[62:0];
    assign _19185 = { _19183,
                      _19184 };
    assign _19186 = _19185 < _22192;
    assign _19187 = ~ _19186;
    assign _19175 = _18687[9:9];
    assign _19172 = _19167 - _22192;
    assign _19173 = _19169 ? _19172 : _19167;
    assign _19174 = _19173[62:0];
    assign _19176 = { _19174,
                      _19175 };
    assign _19177 = _19176 < _22192;
    assign _19178 = ~ _19177;
    assign _19166 = _18687[10:10];
    assign _19163 = _19158 - _22192;
    assign _19164 = _19160 ? _19163 : _19158;
    assign _19165 = _19164[62:0];
    assign _19167 = { _19165,
                      _19166 };
    assign _19168 = _19167 < _22192;
    assign _19169 = ~ _19168;
    assign _19157 = _18687[11:11];
    assign _19154 = _19149 - _22192;
    assign _19155 = _19151 ? _19154 : _19149;
    assign _19156 = _19155[62:0];
    assign _19158 = { _19156,
                      _19157 };
    assign _19159 = _19158 < _22192;
    assign _19160 = ~ _19159;
    assign _19148 = _18687[12:12];
    assign _19145 = _19140 - _22192;
    assign _19146 = _19142 ? _19145 : _19140;
    assign _19147 = _19146[62:0];
    assign _19149 = { _19147,
                      _19148 };
    assign _19150 = _19149 < _22192;
    assign _19151 = ~ _19150;
    assign _19139 = _18687[13:13];
    assign _19136 = _19131 - _22192;
    assign _19137 = _19133 ? _19136 : _19131;
    assign _19138 = _19137[62:0];
    assign _19140 = { _19138,
                      _19139 };
    assign _19141 = _19140 < _22192;
    assign _19142 = ~ _19141;
    assign _19130 = _18687[14:14];
    assign _19127 = _19122 - _22192;
    assign _19128 = _19124 ? _19127 : _19122;
    assign _19129 = _19128[62:0];
    assign _19131 = { _19129,
                      _19130 };
    assign _19132 = _19131 < _22192;
    assign _19133 = ~ _19132;
    assign _19121 = _18687[15:15];
    assign _19118 = _19113 - _22192;
    assign _19119 = _19115 ? _19118 : _19113;
    assign _19120 = _19119[62:0];
    assign _19122 = { _19120,
                      _19121 };
    assign _19123 = _19122 < _22192;
    assign _19124 = ~ _19123;
    assign _19112 = _18687[16:16];
    assign _19109 = _19104 - _22192;
    assign _19110 = _19106 ? _19109 : _19104;
    assign _19111 = _19110[62:0];
    assign _19113 = { _19111,
                      _19112 };
    assign _19114 = _19113 < _22192;
    assign _19115 = ~ _19114;
    assign _19103 = _18687[17:17];
    assign _19100 = _19095 - _22192;
    assign _19101 = _19097 ? _19100 : _19095;
    assign _19102 = _19101[62:0];
    assign _19104 = { _19102,
                      _19103 };
    assign _19105 = _19104 < _22192;
    assign _19106 = ~ _19105;
    assign _19094 = _18687[18:18];
    assign _19091 = _19086 - _22192;
    assign _19092 = _19088 ? _19091 : _19086;
    assign _19093 = _19092[62:0];
    assign _19095 = { _19093,
                      _19094 };
    assign _19096 = _19095 < _22192;
    assign _19097 = ~ _19096;
    assign _19085 = _18687[19:19];
    assign _19082 = _19077 - _22192;
    assign _19083 = _19079 ? _19082 : _19077;
    assign _19084 = _19083[62:0];
    assign _19086 = { _19084,
                      _19085 };
    assign _19087 = _19086 < _22192;
    assign _19088 = ~ _19087;
    assign _19076 = _18687[20:20];
    assign _19073 = _19068 - _22192;
    assign _19074 = _19070 ? _19073 : _19068;
    assign _19075 = _19074[62:0];
    assign _19077 = { _19075,
                      _19076 };
    assign _19078 = _19077 < _22192;
    assign _19079 = ~ _19078;
    assign _19067 = _18687[21:21];
    assign _19064 = _19059 - _22192;
    assign _19065 = _19061 ? _19064 : _19059;
    assign _19066 = _19065[62:0];
    assign _19068 = { _19066,
                      _19067 };
    assign _19069 = _19068 < _22192;
    assign _19070 = ~ _19069;
    assign _19058 = _18687[22:22];
    assign _19055 = _19050 - _22192;
    assign _19056 = _19052 ? _19055 : _19050;
    assign _19057 = _19056[62:0];
    assign _19059 = { _19057,
                      _19058 };
    assign _19060 = _19059 < _22192;
    assign _19061 = ~ _19060;
    assign _19049 = _18687[23:23];
    assign _19046 = _19041 - _22192;
    assign _19047 = _19043 ? _19046 : _19041;
    assign _19048 = _19047[62:0];
    assign _19050 = { _19048,
                      _19049 };
    assign _19051 = _19050 < _22192;
    assign _19052 = ~ _19051;
    assign _19040 = _18687[24:24];
    assign _19037 = _19032 - _22192;
    assign _19038 = _19034 ? _19037 : _19032;
    assign _19039 = _19038[62:0];
    assign _19041 = { _19039,
                      _19040 };
    assign _19042 = _19041 < _22192;
    assign _19043 = ~ _19042;
    assign _19031 = _18687[25:25];
    assign _19028 = _19023 - _22192;
    assign _19029 = _19025 ? _19028 : _19023;
    assign _19030 = _19029[62:0];
    assign _19032 = { _19030,
                      _19031 };
    assign _19033 = _19032 < _22192;
    assign _19034 = ~ _19033;
    assign _19022 = _18687[26:26];
    assign _19019 = _19014 - _22192;
    assign _19020 = _19016 ? _19019 : _19014;
    assign _19021 = _19020[62:0];
    assign _19023 = { _19021,
                      _19022 };
    assign _19024 = _19023 < _22192;
    assign _19025 = ~ _19024;
    assign _19013 = _18687[27:27];
    assign _19010 = _19005 - _22192;
    assign _19011 = _19007 ? _19010 : _19005;
    assign _19012 = _19011[62:0];
    assign _19014 = { _19012,
                      _19013 };
    assign _19015 = _19014 < _22192;
    assign _19016 = ~ _19015;
    assign _19004 = _18687[28:28];
    assign _19001 = _18996 - _22192;
    assign _19002 = _18998 ? _19001 : _18996;
    assign _19003 = _19002[62:0];
    assign _19005 = { _19003,
                      _19004 };
    assign _19006 = _19005 < _22192;
    assign _19007 = ~ _19006;
    assign _18995 = _18687[29:29];
    assign _18992 = _18987 - _22192;
    assign _18993 = _18989 ? _18992 : _18987;
    assign _18994 = _18993[62:0];
    assign _18996 = { _18994,
                      _18995 };
    assign _18997 = _18996 < _22192;
    assign _18998 = ~ _18997;
    assign _18986 = _18687[30:30];
    assign _18983 = _18978 - _22192;
    assign _18984 = _18980 ? _18983 : _18978;
    assign _18985 = _18984[62:0];
    assign _18987 = { _18985,
                      _18986 };
    assign _18988 = _18987 < _22192;
    assign _18989 = ~ _18988;
    assign _18977 = _18687[31:31];
    assign _18974 = _18969 - _22192;
    assign _18975 = _18971 ? _18974 : _18969;
    assign _18976 = _18975[62:0];
    assign _18978 = { _18976,
                      _18977 };
    assign _18979 = _18978 < _22192;
    assign _18980 = ~ _18979;
    assign _18968 = _18687[32:32];
    assign _18965 = _18960 - _22192;
    assign _18966 = _18962 ? _18965 : _18960;
    assign _18967 = _18966[62:0];
    assign _18969 = { _18967,
                      _18968 };
    assign _18970 = _18969 < _22192;
    assign _18971 = ~ _18970;
    assign _18959 = _18687[33:33];
    assign _18956 = _18951 - _22192;
    assign _18957 = _18953 ? _18956 : _18951;
    assign _18958 = _18957[62:0];
    assign _18960 = { _18958,
                      _18959 };
    assign _18961 = _18960 < _22192;
    assign _18962 = ~ _18961;
    assign _18950 = _18687[34:34];
    assign _18947 = _18942 - _22192;
    assign _18948 = _18944 ? _18947 : _18942;
    assign _18949 = _18948[62:0];
    assign _18951 = { _18949,
                      _18950 };
    assign _18952 = _18951 < _22192;
    assign _18953 = ~ _18952;
    assign _18941 = _18687[35:35];
    assign _18938 = _18933 - _22192;
    assign _18939 = _18935 ? _18938 : _18933;
    assign _18940 = _18939[62:0];
    assign _18942 = { _18940,
                      _18941 };
    assign _18943 = _18942 < _22192;
    assign _18944 = ~ _18943;
    assign _18932 = _18687[36:36];
    assign _18929 = _18924 - _22192;
    assign _18930 = _18926 ? _18929 : _18924;
    assign _18931 = _18930[62:0];
    assign _18933 = { _18931,
                      _18932 };
    assign _18934 = _18933 < _22192;
    assign _18935 = ~ _18934;
    assign _18923 = _18687[37:37];
    assign _18920 = _18915 - _22192;
    assign _18921 = _18917 ? _18920 : _18915;
    assign _18922 = _18921[62:0];
    assign _18924 = { _18922,
                      _18923 };
    assign _18925 = _18924 < _22192;
    assign _18926 = ~ _18925;
    assign _18914 = _18687[38:38];
    assign _18911 = _18906 - _22192;
    assign _18912 = _18908 ? _18911 : _18906;
    assign _18913 = _18912[62:0];
    assign _18915 = { _18913,
                      _18914 };
    assign _18916 = _18915 < _22192;
    assign _18917 = ~ _18916;
    assign _18905 = _18687[39:39];
    assign _18902 = _18897 - _22192;
    assign _18903 = _18899 ? _18902 : _18897;
    assign _18904 = _18903[62:0];
    assign _18906 = { _18904,
                      _18905 };
    assign _18907 = _18906 < _22192;
    assign _18908 = ~ _18907;
    assign _18896 = _18687[40:40];
    assign _18893 = _18888 - _22192;
    assign _18894 = _18890 ? _18893 : _18888;
    assign _18895 = _18894[62:0];
    assign _18897 = { _18895,
                      _18896 };
    assign _18898 = _18897 < _22192;
    assign _18899 = ~ _18898;
    assign _18887 = _18687[41:41];
    assign _18884 = _18879 - _22192;
    assign _18885 = _18881 ? _18884 : _18879;
    assign _18886 = _18885[62:0];
    assign _18888 = { _18886,
                      _18887 };
    assign _18889 = _18888 < _22192;
    assign _18890 = ~ _18889;
    assign _18878 = _18687[42:42];
    assign _18875 = _18870 - _22192;
    assign _18876 = _18872 ? _18875 : _18870;
    assign _18877 = _18876[62:0];
    assign _18879 = { _18877,
                      _18878 };
    assign _18880 = _18879 < _22192;
    assign _18881 = ~ _18880;
    assign _18869 = _18687[43:43];
    assign _18866 = _18861 - _22192;
    assign _18867 = _18863 ? _18866 : _18861;
    assign _18868 = _18867[62:0];
    assign _18870 = { _18868,
                      _18869 };
    assign _18871 = _18870 < _22192;
    assign _18872 = ~ _18871;
    assign _18860 = _18687[44:44];
    assign _18857 = _18852 - _22192;
    assign _18858 = _18854 ? _18857 : _18852;
    assign _18859 = _18858[62:0];
    assign _18861 = { _18859,
                      _18860 };
    assign _18862 = _18861 < _22192;
    assign _18863 = ~ _18862;
    assign _18851 = _18687[45:45];
    assign _18848 = _18843 - _22192;
    assign _18849 = _18845 ? _18848 : _18843;
    assign _18850 = _18849[62:0];
    assign _18852 = { _18850,
                      _18851 };
    assign _18853 = _18852 < _22192;
    assign _18854 = ~ _18853;
    assign _18842 = _18687[46:46];
    assign _18839 = _18834 - _22192;
    assign _18840 = _18836 ? _18839 : _18834;
    assign _18841 = _18840[62:0];
    assign _18843 = { _18841,
                      _18842 };
    assign _18844 = _18843 < _22192;
    assign _18845 = ~ _18844;
    assign _18833 = _18687[47:47];
    assign _18830 = _18825 - _22192;
    assign _18831 = _18827 ? _18830 : _18825;
    assign _18832 = _18831[62:0];
    assign _18834 = { _18832,
                      _18833 };
    assign _18835 = _18834 < _22192;
    assign _18836 = ~ _18835;
    assign _18824 = _18687[48:48];
    assign _18821 = _18816 - _22192;
    assign _18822 = _18818 ? _18821 : _18816;
    assign _18823 = _18822[62:0];
    assign _18825 = { _18823,
                      _18824 };
    assign _18826 = _18825 < _22192;
    assign _18827 = ~ _18826;
    assign _18815 = _18687[49:49];
    assign _18812 = _18807 - _22192;
    assign _18813 = _18809 ? _18812 : _18807;
    assign _18814 = _18813[62:0];
    assign _18816 = { _18814,
                      _18815 };
    assign _18817 = _18816 < _22192;
    assign _18818 = ~ _18817;
    assign _18806 = _18687[50:50];
    assign _18803 = _18798 - _22192;
    assign _18804 = _18800 ? _18803 : _18798;
    assign _18805 = _18804[62:0];
    assign _18807 = { _18805,
                      _18806 };
    assign _18808 = _18807 < _22192;
    assign _18809 = ~ _18808;
    assign _18797 = _18687[51:51];
    assign _18794 = _18789 - _22192;
    assign _18795 = _18791 ? _18794 : _18789;
    assign _18796 = _18795[62:0];
    assign _18798 = { _18796,
                      _18797 };
    assign _18799 = _18798 < _22192;
    assign _18800 = ~ _18799;
    assign _18788 = _18687[52:52];
    assign _18785 = _18780 - _22192;
    assign _18786 = _18782 ? _18785 : _18780;
    assign _18787 = _18786[62:0];
    assign _18789 = { _18787,
                      _18788 };
    assign _18790 = _18789 < _22192;
    assign _18791 = ~ _18790;
    assign _18779 = _18687[53:53];
    assign _18776 = _18771 - _22192;
    assign _18777 = _18773 ? _18776 : _18771;
    assign _18778 = _18777[62:0];
    assign _18780 = { _18778,
                      _18779 };
    assign _18781 = _18780 < _22192;
    assign _18782 = ~ _18781;
    assign _18770 = _18687[54:54];
    assign _18767 = _18762 - _22192;
    assign _18768 = _18764 ? _18767 : _18762;
    assign _18769 = _18768[62:0];
    assign _18771 = { _18769,
                      _18770 };
    assign _18772 = _18771 < _22192;
    assign _18773 = ~ _18772;
    assign _18761 = _18687[55:55];
    assign _18758 = _18753 - _22192;
    assign _18759 = _18755 ? _18758 : _18753;
    assign _18760 = _18759[62:0];
    assign _18762 = { _18760,
                      _18761 };
    assign _18763 = _18762 < _22192;
    assign _18764 = ~ _18763;
    assign _18752 = _18687[56:56];
    assign _18749 = _18744 - _22192;
    assign _18750 = _18746 ? _18749 : _18744;
    assign _18751 = _18750[62:0];
    assign _18753 = { _18751,
                      _18752 };
    assign _18754 = _18753 < _22192;
    assign _18755 = ~ _18754;
    assign _18743 = _18687[57:57];
    assign _18740 = _18735 - _22192;
    assign _18741 = _18737 ? _18740 : _18735;
    assign _18742 = _18741[62:0];
    assign _18744 = { _18742,
                      _18743 };
    assign _18745 = _18744 < _22192;
    assign _18746 = ~ _18745;
    assign _18734 = _18687[58:58];
    assign _18731 = _18726 - _22192;
    assign _18732 = _18728 ? _18731 : _18726;
    assign _18733 = _18732[62:0];
    assign _18735 = { _18733,
                      _18734 };
    assign _18736 = _18735 < _22192;
    assign _18737 = ~ _18736;
    assign _18725 = _18687[59:59];
    assign _18722 = _18717 - _22192;
    assign _18723 = _18719 ? _18722 : _18717;
    assign _18724 = _18723[62:0];
    assign _18726 = { _18724,
                      _18725 };
    assign _18727 = _18726 < _22192;
    assign _18728 = ~ _18727;
    assign _18716 = _18687[60:60];
    assign _18713 = _18708 - _22192;
    assign _18714 = _18710 ? _18713 : _18708;
    assign _18715 = _18714[62:0];
    assign _18717 = { _18715,
                      _18716 };
    assign _18718 = _18717 < _22192;
    assign _18719 = ~ _18718;
    assign _18707 = _18687[61:61];
    assign _18704 = _18699 - _22192;
    assign _18705 = _18701 ? _18704 : _18699;
    assign _18706 = _18705[62:0];
    assign _18708 = { _18706,
                      _18707 };
    assign _18709 = _18708 < _22192;
    assign _18710 = ~ _18709;
    assign _18698 = _18687[62:62];
    assign _18695 = _18689 - _22192;
    assign _18696 = _18692 ? _18695 : _18689;
    assign _18697 = _18696[62:0];
    assign _18699 = { _18697,
                      _18698 };
    assign _18700 = _18699 < _22192;
    assign _18701 = ~ _18700;
    assign _18685 = _18677 + _22186;
    assign _18686 = _18677 * _18685;
    assign _18687 = _18686[63:0];
    assign _18688 = _18687[63:63];
    assign _18689 = { _22185,
                      _18688 };
    assign _18691 = _18689 < _22192;
    assign _18692 = ~ _18691;
    assign _18693 = { _22185,
                      _18692 };
    assign _18694 = _18693[62:0];
    assign _18702 = { _18694,
                      _18701 };
    assign _18703 = _18702[62:0];
    assign _18711 = { _18703,
                      _18710 };
    assign _18712 = _18711[62:0];
    assign _18720 = { _18712,
                      _18719 };
    assign _18721 = _18720[62:0];
    assign _18729 = { _18721,
                      _18728 };
    assign _18730 = _18729[62:0];
    assign _18738 = { _18730,
                      _18737 };
    assign _18739 = _18738[62:0];
    assign _18747 = { _18739,
                      _18746 };
    assign _18748 = _18747[62:0];
    assign _18756 = { _18748,
                      _18755 };
    assign _18757 = _18756[62:0];
    assign _18765 = { _18757,
                      _18764 };
    assign _18766 = _18765[62:0];
    assign _18774 = { _18766,
                      _18773 };
    assign _18775 = _18774[62:0];
    assign _18783 = { _18775,
                      _18782 };
    assign _18784 = _18783[62:0];
    assign _18792 = { _18784,
                      _18791 };
    assign _18793 = _18792[62:0];
    assign _18801 = { _18793,
                      _18800 };
    assign _18802 = _18801[62:0];
    assign _18810 = { _18802,
                      _18809 };
    assign _18811 = _18810[62:0];
    assign _18819 = { _18811,
                      _18818 };
    assign _18820 = _18819[62:0];
    assign _18828 = { _18820,
                      _18827 };
    assign _18829 = _18828[62:0];
    assign _18837 = { _18829,
                      _18836 };
    assign _18838 = _18837[62:0];
    assign _18846 = { _18838,
                      _18845 };
    assign _18847 = _18846[62:0];
    assign _18855 = { _18847,
                      _18854 };
    assign _18856 = _18855[62:0];
    assign _18864 = { _18856,
                      _18863 };
    assign _18865 = _18864[62:0];
    assign _18873 = { _18865,
                      _18872 };
    assign _18874 = _18873[62:0];
    assign _18882 = { _18874,
                      _18881 };
    assign _18883 = _18882[62:0];
    assign _18891 = { _18883,
                      _18890 };
    assign _18892 = _18891[62:0];
    assign _18900 = { _18892,
                      _18899 };
    assign _18901 = _18900[62:0];
    assign _18909 = { _18901,
                      _18908 };
    assign _18910 = _18909[62:0];
    assign _18918 = { _18910,
                      _18917 };
    assign _18919 = _18918[62:0];
    assign _18927 = { _18919,
                      _18926 };
    assign _18928 = _18927[62:0];
    assign _18936 = { _18928,
                      _18935 };
    assign _18937 = _18936[62:0];
    assign _18945 = { _18937,
                      _18944 };
    assign _18946 = _18945[62:0];
    assign _18954 = { _18946,
                      _18953 };
    assign _18955 = _18954[62:0];
    assign _18963 = { _18955,
                      _18962 };
    assign _18964 = _18963[62:0];
    assign _18972 = { _18964,
                      _18971 };
    assign _18973 = _18972[62:0];
    assign _18981 = { _18973,
                      _18980 };
    assign _18982 = _18981[62:0];
    assign _18990 = { _18982,
                      _18989 };
    assign _18991 = _18990[62:0];
    assign _18999 = { _18991,
                      _18998 };
    assign _19000 = _18999[62:0];
    assign _19008 = { _19000,
                      _19007 };
    assign _19009 = _19008[62:0];
    assign _19017 = { _19009,
                      _19016 };
    assign _19018 = _19017[62:0];
    assign _19026 = { _19018,
                      _19025 };
    assign _19027 = _19026[62:0];
    assign _19035 = { _19027,
                      _19034 };
    assign _19036 = _19035[62:0];
    assign _19044 = { _19036,
                      _19043 };
    assign _19045 = _19044[62:0];
    assign _19053 = { _19045,
                      _19052 };
    assign _19054 = _19053[62:0];
    assign _19062 = { _19054,
                      _19061 };
    assign _19063 = _19062[62:0];
    assign _19071 = { _19063,
                      _19070 };
    assign _19072 = _19071[62:0];
    assign _19080 = { _19072,
                      _19079 };
    assign _19081 = _19080[62:0];
    assign _19089 = { _19081,
                      _19088 };
    assign _19090 = _19089[62:0];
    assign _19098 = { _19090,
                      _19097 };
    assign _19099 = _19098[62:0];
    assign _19107 = { _19099,
                      _19106 };
    assign _19108 = _19107[62:0];
    assign _19116 = { _19108,
                      _19115 };
    assign _19117 = _19116[62:0];
    assign _19125 = { _19117,
                      _19124 };
    assign _19126 = _19125[62:0];
    assign _19134 = { _19126,
                      _19133 };
    assign _19135 = _19134[62:0];
    assign _19143 = { _19135,
                      _19142 };
    assign _19144 = _19143[62:0];
    assign _19152 = { _19144,
                      _19151 };
    assign _19153 = _19152[62:0];
    assign _19161 = { _19153,
                      _19160 };
    assign _19162 = _19161[62:0];
    assign _19170 = { _19162,
                      _19169 };
    assign _19171 = _19170[62:0];
    assign _19179 = { _19171,
                      _19178 };
    assign _19180 = _19179[62:0];
    assign _19188 = { _19180,
                      _19187 };
    assign _19189 = _19188[62:0];
    assign _19197 = { _19189,
                      _19196 };
    assign _19198 = _19197[62:0];
    assign _19206 = { _19198,
                      _19205 };
    assign _19207 = _19206[62:0];
    assign _19215 = { _19207,
                      _19214 };
    assign _19216 = _19215[62:0];
    assign _19224 = { _19216,
                      _19223 };
    assign _19225 = _19224[62:0];
    assign _19233 = { _19225,
                      _19232 };
    assign _19234 = _19233[62:0];
    assign _19242 = { _19234,
                      _19241 };
    assign _19243 = _19242[62:0];
    assign _19251 = { _19243,
                      _19250 };
    assign _19252 = _19251[62:0];
    assign _19260 = { _19252,
                      _19259 };
    assign _19261 = _17525 * _19260;
    assign _19262 = _19261[63:0];
    assign _18673 = _18105[0:0];
    assign _18670 = _18665 - _17525;
    assign _18671 = _18667 ? _18670 : _18665;
    assign _18672 = _18671[62:0];
    assign _18674 = { _18672,
                      _18673 };
    assign _18675 = _18674 < _17525;
    assign _18676 = ~ _18675;
    assign _18664 = _18105[1:1];
    assign _18661 = _18656 - _17525;
    assign _18662 = _18658 ? _18661 : _18656;
    assign _18663 = _18662[62:0];
    assign _18665 = { _18663,
                      _18664 };
    assign _18666 = _18665 < _17525;
    assign _18667 = ~ _18666;
    assign _18655 = _18105[2:2];
    assign _18652 = _18647 - _17525;
    assign _18653 = _18649 ? _18652 : _18647;
    assign _18654 = _18653[62:0];
    assign _18656 = { _18654,
                      _18655 };
    assign _18657 = _18656 < _17525;
    assign _18658 = ~ _18657;
    assign _18646 = _18105[3:3];
    assign _18643 = _18638 - _17525;
    assign _18644 = _18640 ? _18643 : _18638;
    assign _18645 = _18644[62:0];
    assign _18647 = { _18645,
                      _18646 };
    assign _18648 = _18647 < _17525;
    assign _18649 = ~ _18648;
    assign _18637 = _18105[4:4];
    assign _18634 = _18629 - _17525;
    assign _18635 = _18631 ? _18634 : _18629;
    assign _18636 = _18635[62:0];
    assign _18638 = { _18636,
                      _18637 };
    assign _18639 = _18638 < _17525;
    assign _18640 = ~ _18639;
    assign _18628 = _18105[5:5];
    assign _18625 = _18620 - _17525;
    assign _18626 = _18622 ? _18625 : _18620;
    assign _18627 = _18626[62:0];
    assign _18629 = { _18627,
                      _18628 };
    assign _18630 = _18629 < _17525;
    assign _18631 = ~ _18630;
    assign _18619 = _18105[6:6];
    assign _18616 = _18611 - _17525;
    assign _18617 = _18613 ? _18616 : _18611;
    assign _18618 = _18617[62:0];
    assign _18620 = { _18618,
                      _18619 };
    assign _18621 = _18620 < _17525;
    assign _18622 = ~ _18621;
    assign _18610 = _18105[7:7];
    assign _18607 = _18602 - _17525;
    assign _18608 = _18604 ? _18607 : _18602;
    assign _18609 = _18608[62:0];
    assign _18611 = { _18609,
                      _18610 };
    assign _18612 = _18611 < _17525;
    assign _18613 = ~ _18612;
    assign _18601 = _18105[8:8];
    assign _18598 = _18593 - _17525;
    assign _18599 = _18595 ? _18598 : _18593;
    assign _18600 = _18599[62:0];
    assign _18602 = { _18600,
                      _18601 };
    assign _18603 = _18602 < _17525;
    assign _18604 = ~ _18603;
    assign _18592 = _18105[9:9];
    assign _18589 = _18584 - _17525;
    assign _18590 = _18586 ? _18589 : _18584;
    assign _18591 = _18590[62:0];
    assign _18593 = { _18591,
                      _18592 };
    assign _18594 = _18593 < _17525;
    assign _18595 = ~ _18594;
    assign _18583 = _18105[10:10];
    assign _18580 = _18575 - _17525;
    assign _18581 = _18577 ? _18580 : _18575;
    assign _18582 = _18581[62:0];
    assign _18584 = { _18582,
                      _18583 };
    assign _18585 = _18584 < _17525;
    assign _18586 = ~ _18585;
    assign _18574 = _18105[11:11];
    assign _18571 = _18566 - _17525;
    assign _18572 = _18568 ? _18571 : _18566;
    assign _18573 = _18572[62:0];
    assign _18575 = { _18573,
                      _18574 };
    assign _18576 = _18575 < _17525;
    assign _18577 = ~ _18576;
    assign _18565 = _18105[12:12];
    assign _18562 = _18557 - _17525;
    assign _18563 = _18559 ? _18562 : _18557;
    assign _18564 = _18563[62:0];
    assign _18566 = { _18564,
                      _18565 };
    assign _18567 = _18566 < _17525;
    assign _18568 = ~ _18567;
    assign _18556 = _18105[13:13];
    assign _18553 = _18548 - _17525;
    assign _18554 = _18550 ? _18553 : _18548;
    assign _18555 = _18554[62:0];
    assign _18557 = { _18555,
                      _18556 };
    assign _18558 = _18557 < _17525;
    assign _18559 = ~ _18558;
    assign _18547 = _18105[14:14];
    assign _18544 = _18539 - _17525;
    assign _18545 = _18541 ? _18544 : _18539;
    assign _18546 = _18545[62:0];
    assign _18548 = { _18546,
                      _18547 };
    assign _18549 = _18548 < _17525;
    assign _18550 = ~ _18549;
    assign _18538 = _18105[15:15];
    assign _18535 = _18530 - _17525;
    assign _18536 = _18532 ? _18535 : _18530;
    assign _18537 = _18536[62:0];
    assign _18539 = { _18537,
                      _18538 };
    assign _18540 = _18539 < _17525;
    assign _18541 = ~ _18540;
    assign _18529 = _18105[16:16];
    assign _18526 = _18521 - _17525;
    assign _18527 = _18523 ? _18526 : _18521;
    assign _18528 = _18527[62:0];
    assign _18530 = { _18528,
                      _18529 };
    assign _18531 = _18530 < _17525;
    assign _18532 = ~ _18531;
    assign _18520 = _18105[17:17];
    assign _18517 = _18512 - _17525;
    assign _18518 = _18514 ? _18517 : _18512;
    assign _18519 = _18518[62:0];
    assign _18521 = { _18519,
                      _18520 };
    assign _18522 = _18521 < _17525;
    assign _18523 = ~ _18522;
    assign _18511 = _18105[18:18];
    assign _18508 = _18503 - _17525;
    assign _18509 = _18505 ? _18508 : _18503;
    assign _18510 = _18509[62:0];
    assign _18512 = { _18510,
                      _18511 };
    assign _18513 = _18512 < _17525;
    assign _18514 = ~ _18513;
    assign _18502 = _18105[19:19];
    assign _18499 = _18494 - _17525;
    assign _18500 = _18496 ? _18499 : _18494;
    assign _18501 = _18500[62:0];
    assign _18503 = { _18501,
                      _18502 };
    assign _18504 = _18503 < _17525;
    assign _18505 = ~ _18504;
    assign _18493 = _18105[20:20];
    assign _18490 = _18485 - _17525;
    assign _18491 = _18487 ? _18490 : _18485;
    assign _18492 = _18491[62:0];
    assign _18494 = { _18492,
                      _18493 };
    assign _18495 = _18494 < _17525;
    assign _18496 = ~ _18495;
    assign _18484 = _18105[21:21];
    assign _18481 = _18476 - _17525;
    assign _18482 = _18478 ? _18481 : _18476;
    assign _18483 = _18482[62:0];
    assign _18485 = { _18483,
                      _18484 };
    assign _18486 = _18485 < _17525;
    assign _18487 = ~ _18486;
    assign _18475 = _18105[22:22];
    assign _18472 = _18467 - _17525;
    assign _18473 = _18469 ? _18472 : _18467;
    assign _18474 = _18473[62:0];
    assign _18476 = { _18474,
                      _18475 };
    assign _18477 = _18476 < _17525;
    assign _18478 = ~ _18477;
    assign _18466 = _18105[23:23];
    assign _18463 = _18458 - _17525;
    assign _18464 = _18460 ? _18463 : _18458;
    assign _18465 = _18464[62:0];
    assign _18467 = { _18465,
                      _18466 };
    assign _18468 = _18467 < _17525;
    assign _18469 = ~ _18468;
    assign _18457 = _18105[24:24];
    assign _18454 = _18449 - _17525;
    assign _18455 = _18451 ? _18454 : _18449;
    assign _18456 = _18455[62:0];
    assign _18458 = { _18456,
                      _18457 };
    assign _18459 = _18458 < _17525;
    assign _18460 = ~ _18459;
    assign _18448 = _18105[25:25];
    assign _18445 = _18440 - _17525;
    assign _18446 = _18442 ? _18445 : _18440;
    assign _18447 = _18446[62:0];
    assign _18449 = { _18447,
                      _18448 };
    assign _18450 = _18449 < _17525;
    assign _18451 = ~ _18450;
    assign _18439 = _18105[26:26];
    assign _18436 = _18431 - _17525;
    assign _18437 = _18433 ? _18436 : _18431;
    assign _18438 = _18437[62:0];
    assign _18440 = { _18438,
                      _18439 };
    assign _18441 = _18440 < _17525;
    assign _18442 = ~ _18441;
    assign _18430 = _18105[27:27];
    assign _18427 = _18422 - _17525;
    assign _18428 = _18424 ? _18427 : _18422;
    assign _18429 = _18428[62:0];
    assign _18431 = { _18429,
                      _18430 };
    assign _18432 = _18431 < _17525;
    assign _18433 = ~ _18432;
    assign _18421 = _18105[28:28];
    assign _18418 = _18413 - _17525;
    assign _18419 = _18415 ? _18418 : _18413;
    assign _18420 = _18419[62:0];
    assign _18422 = { _18420,
                      _18421 };
    assign _18423 = _18422 < _17525;
    assign _18424 = ~ _18423;
    assign _18412 = _18105[29:29];
    assign _18409 = _18404 - _17525;
    assign _18410 = _18406 ? _18409 : _18404;
    assign _18411 = _18410[62:0];
    assign _18413 = { _18411,
                      _18412 };
    assign _18414 = _18413 < _17525;
    assign _18415 = ~ _18414;
    assign _18403 = _18105[30:30];
    assign _18400 = _18395 - _17525;
    assign _18401 = _18397 ? _18400 : _18395;
    assign _18402 = _18401[62:0];
    assign _18404 = { _18402,
                      _18403 };
    assign _18405 = _18404 < _17525;
    assign _18406 = ~ _18405;
    assign _18394 = _18105[31:31];
    assign _18391 = _18386 - _17525;
    assign _18392 = _18388 ? _18391 : _18386;
    assign _18393 = _18392[62:0];
    assign _18395 = { _18393,
                      _18394 };
    assign _18396 = _18395 < _17525;
    assign _18397 = ~ _18396;
    assign _18385 = _18105[32:32];
    assign _18382 = _18377 - _17525;
    assign _18383 = _18379 ? _18382 : _18377;
    assign _18384 = _18383[62:0];
    assign _18386 = { _18384,
                      _18385 };
    assign _18387 = _18386 < _17525;
    assign _18388 = ~ _18387;
    assign _18376 = _18105[33:33];
    assign _18373 = _18368 - _17525;
    assign _18374 = _18370 ? _18373 : _18368;
    assign _18375 = _18374[62:0];
    assign _18377 = { _18375,
                      _18376 };
    assign _18378 = _18377 < _17525;
    assign _18379 = ~ _18378;
    assign _18367 = _18105[34:34];
    assign _18364 = _18359 - _17525;
    assign _18365 = _18361 ? _18364 : _18359;
    assign _18366 = _18365[62:0];
    assign _18368 = { _18366,
                      _18367 };
    assign _18369 = _18368 < _17525;
    assign _18370 = ~ _18369;
    assign _18358 = _18105[35:35];
    assign _18355 = _18350 - _17525;
    assign _18356 = _18352 ? _18355 : _18350;
    assign _18357 = _18356[62:0];
    assign _18359 = { _18357,
                      _18358 };
    assign _18360 = _18359 < _17525;
    assign _18361 = ~ _18360;
    assign _18349 = _18105[36:36];
    assign _18346 = _18341 - _17525;
    assign _18347 = _18343 ? _18346 : _18341;
    assign _18348 = _18347[62:0];
    assign _18350 = { _18348,
                      _18349 };
    assign _18351 = _18350 < _17525;
    assign _18352 = ~ _18351;
    assign _18340 = _18105[37:37];
    assign _18337 = _18332 - _17525;
    assign _18338 = _18334 ? _18337 : _18332;
    assign _18339 = _18338[62:0];
    assign _18341 = { _18339,
                      _18340 };
    assign _18342 = _18341 < _17525;
    assign _18343 = ~ _18342;
    assign _18331 = _18105[38:38];
    assign _18328 = _18323 - _17525;
    assign _18329 = _18325 ? _18328 : _18323;
    assign _18330 = _18329[62:0];
    assign _18332 = { _18330,
                      _18331 };
    assign _18333 = _18332 < _17525;
    assign _18334 = ~ _18333;
    assign _18322 = _18105[39:39];
    assign _18319 = _18314 - _17525;
    assign _18320 = _18316 ? _18319 : _18314;
    assign _18321 = _18320[62:0];
    assign _18323 = { _18321,
                      _18322 };
    assign _18324 = _18323 < _17525;
    assign _18325 = ~ _18324;
    assign _18313 = _18105[40:40];
    assign _18310 = _18305 - _17525;
    assign _18311 = _18307 ? _18310 : _18305;
    assign _18312 = _18311[62:0];
    assign _18314 = { _18312,
                      _18313 };
    assign _18315 = _18314 < _17525;
    assign _18316 = ~ _18315;
    assign _18304 = _18105[41:41];
    assign _18301 = _18296 - _17525;
    assign _18302 = _18298 ? _18301 : _18296;
    assign _18303 = _18302[62:0];
    assign _18305 = { _18303,
                      _18304 };
    assign _18306 = _18305 < _17525;
    assign _18307 = ~ _18306;
    assign _18295 = _18105[42:42];
    assign _18292 = _18287 - _17525;
    assign _18293 = _18289 ? _18292 : _18287;
    assign _18294 = _18293[62:0];
    assign _18296 = { _18294,
                      _18295 };
    assign _18297 = _18296 < _17525;
    assign _18298 = ~ _18297;
    assign _18286 = _18105[43:43];
    assign _18283 = _18278 - _17525;
    assign _18284 = _18280 ? _18283 : _18278;
    assign _18285 = _18284[62:0];
    assign _18287 = { _18285,
                      _18286 };
    assign _18288 = _18287 < _17525;
    assign _18289 = ~ _18288;
    assign _18277 = _18105[44:44];
    assign _18274 = _18269 - _17525;
    assign _18275 = _18271 ? _18274 : _18269;
    assign _18276 = _18275[62:0];
    assign _18278 = { _18276,
                      _18277 };
    assign _18279 = _18278 < _17525;
    assign _18280 = ~ _18279;
    assign _18268 = _18105[45:45];
    assign _18265 = _18260 - _17525;
    assign _18266 = _18262 ? _18265 : _18260;
    assign _18267 = _18266[62:0];
    assign _18269 = { _18267,
                      _18268 };
    assign _18270 = _18269 < _17525;
    assign _18271 = ~ _18270;
    assign _18259 = _18105[46:46];
    assign _18256 = _18251 - _17525;
    assign _18257 = _18253 ? _18256 : _18251;
    assign _18258 = _18257[62:0];
    assign _18260 = { _18258,
                      _18259 };
    assign _18261 = _18260 < _17525;
    assign _18262 = ~ _18261;
    assign _18250 = _18105[47:47];
    assign _18247 = _18242 - _17525;
    assign _18248 = _18244 ? _18247 : _18242;
    assign _18249 = _18248[62:0];
    assign _18251 = { _18249,
                      _18250 };
    assign _18252 = _18251 < _17525;
    assign _18253 = ~ _18252;
    assign _18241 = _18105[48:48];
    assign _18238 = _18233 - _17525;
    assign _18239 = _18235 ? _18238 : _18233;
    assign _18240 = _18239[62:0];
    assign _18242 = { _18240,
                      _18241 };
    assign _18243 = _18242 < _17525;
    assign _18244 = ~ _18243;
    assign _18232 = _18105[49:49];
    assign _18229 = _18224 - _17525;
    assign _18230 = _18226 ? _18229 : _18224;
    assign _18231 = _18230[62:0];
    assign _18233 = { _18231,
                      _18232 };
    assign _18234 = _18233 < _17525;
    assign _18235 = ~ _18234;
    assign _18223 = _18105[50:50];
    assign _18220 = _18215 - _17525;
    assign _18221 = _18217 ? _18220 : _18215;
    assign _18222 = _18221[62:0];
    assign _18224 = { _18222,
                      _18223 };
    assign _18225 = _18224 < _17525;
    assign _18226 = ~ _18225;
    assign _18214 = _18105[51:51];
    assign _18211 = _18206 - _17525;
    assign _18212 = _18208 ? _18211 : _18206;
    assign _18213 = _18212[62:0];
    assign _18215 = { _18213,
                      _18214 };
    assign _18216 = _18215 < _17525;
    assign _18217 = ~ _18216;
    assign _18205 = _18105[52:52];
    assign _18202 = _18197 - _17525;
    assign _18203 = _18199 ? _18202 : _18197;
    assign _18204 = _18203[62:0];
    assign _18206 = { _18204,
                      _18205 };
    assign _18207 = _18206 < _17525;
    assign _18208 = ~ _18207;
    assign _18196 = _18105[53:53];
    assign _18193 = _18188 - _17525;
    assign _18194 = _18190 ? _18193 : _18188;
    assign _18195 = _18194[62:0];
    assign _18197 = { _18195,
                      _18196 };
    assign _18198 = _18197 < _17525;
    assign _18199 = ~ _18198;
    assign _18187 = _18105[54:54];
    assign _18184 = _18179 - _17525;
    assign _18185 = _18181 ? _18184 : _18179;
    assign _18186 = _18185[62:0];
    assign _18188 = { _18186,
                      _18187 };
    assign _18189 = _18188 < _17525;
    assign _18190 = ~ _18189;
    assign _18178 = _18105[55:55];
    assign _18175 = _18170 - _17525;
    assign _18176 = _18172 ? _18175 : _18170;
    assign _18177 = _18176[62:0];
    assign _18179 = { _18177,
                      _18178 };
    assign _18180 = _18179 < _17525;
    assign _18181 = ~ _18180;
    assign _18169 = _18105[56:56];
    assign _18166 = _18161 - _17525;
    assign _18167 = _18163 ? _18166 : _18161;
    assign _18168 = _18167[62:0];
    assign _18170 = { _18168,
                      _18169 };
    assign _18171 = _18170 < _17525;
    assign _18172 = ~ _18171;
    assign _18160 = _18105[57:57];
    assign _18157 = _18152 - _17525;
    assign _18158 = _18154 ? _18157 : _18152;
    assign _18159 = _18158[62:0];
    assign _18161 = { _18159,
                      _18160 };
    assign _18162 = _18161 < _17525;
    assign _18163 = ~ _18162;
    assign _18151 = _18105[58:58];
    assign _18148 = _18143 - _17525;
    assign _18149 = _18145 ? _18148 : _18143;
    assign _18150 = _18149[62:0];
    assign _18152 = { _18150,
                      _18151 };
    assign _18153 = _18152 < _17525;
    assign _18154 = ~ _18153;
    assign _18142 = _18105[59:59];
    assign _18139 = _18134 - _17525;
    assign _18140 = _18136 ? _18139 : _18134;
    assign _18141 = _18140[62:0];
    assign _18143 = { _18141,
                      _18142 };
    assign _18144 = _18143 < _17525;
    assign _18145 = ~ _18144;
    assign _18133 = _18105[60:60];
    assign _18130 = _18125 - _17525;
    assign _18131 = _18127 ? _18130 : _18125;
    assign _18132 = _18131[62:0];
    assign _18134 = { _18132,
                      _18133 };
    assign _18135 = _18134 < _17525;
    assign _18136 = ~ _18135;
    assign _18124 = _18105[61:61];
    assign _18121 = _18116 - _17525;
    assign _18122 = _18118 ? _18121 : _18116;
    assign _18123 = _18122[62:0];
    assign _18125 = { _18123,
                      _18124 };
    assign _18126 = _18125 < _17525;
    assign _18127 = ~ _18126;
    assign _18115 = _18105[62:62];
    assign _18112 = _18107 - _17525;
    assign _18113 = _18109 ? _18112 : _18107;
    assign _18114 = _18113[62:0];
    assign _18116 = { _18114,
                      _18115 };
    assign _18117 = _18116 < _17525;
    assign _18118 = ~ _18117;
    assign _18105 = _17517 - _18099;
    assign _18106 = _18105[63:63];
    assign _18107 = { _22185,
                      _18106 };
    assign _18108 = _18107 < _17525;
    assign _18109 = ~ _18108;
    assign _18110 = { _22185,
                      _18109 };
    assign _18111 = _18110[62:0];
    assign _18119 = { _18111,
                      _18118 };
    assign _18120 = _18119[62:0];
    assign _18128 = { _18120,
                      _18127 };
    assign _18129 = _18128[62:0];
    assign _18137 = { _18129,
                      _18136 };
    assign _18138 = _18137[62:0];
    assign _18146 = { _18138,
                      _18145 };
    assign _18147 = _18146[62:0];
    assign _18155 = { _18147,
                      _18154 };
    assign _18156 = _18155[62:0];
    assign _18164 = { _18156,
                      _18163 };
    assign _18165 = _18164[62:0];
    assign _18173 = { _18165,
                      _18172 };
    assign _18174 = _18173[62:0];
    assign _18182 = { _18174,
                      _18181 };
    assign _18183 = _18182[62:0];
    assign _18191 = { _18183,
                      _18190 };
    assign _18192 = _18191[62:0];
    assign _18200 = { _18192,
                      _18199 };
    assign _18201 = _18200[62:0];
    assign _18209 = { _18201,
                      _18208 };
    assign _18210 = _18209[62:0];
    assign _18218 = { _18210,
                      _18217 };
    assign _18219 = _18218[62:0];
    assign _18227 = { _18219,
                      _18226 };
    assign _18228 = _18227[62:0];
    assign _18236 = { _18228,
                      _18235 };
    assign _18237 = _18236[62:0];
    assign _18245 = { _18237,
                      _18244 };
    assign _18246 = _18245[62:0];
    assign _18254 = { _18246,
                      _18253 };
    assign _18255 = _18254[62:0];
    assign _18263 = { _18255,
                      _18262 };
    assign _18264 = _18263[62:0];
    assign _18272 = { _18264,
                      _18271 };
    assign _18273 = _18272[62:0];
    assign _18281 = { _18273,
                      _18280 };
    assign _18282 = _18281[62:0];
    assign _18290 = { _18282,
                      _18289 };
    assign _18291 = _18290[62:0];
    assign _18299 = { _18291,
                      _18298 };
    assign _18300 = _18299[62:0];
    assign _18308 = { _18300,
                      _18307 };
    assign _18309 = _18308[62:0];
    assign _18317 = { _18309,
                      _18316 };
    assign _18318 = _18317[62:0];
    assign _18326 = { _18318,
                      _18325 };
    assign _18327 = _18326[62:0];
    assign _18335 = { _18327,
                      _18334 };
    assign _18336 = _18335[62:0];
    assign _18344 = { _18336,
                      _18343 };
    assign _18345 = _18344[62:0];
    assign _18353 = { _18345,
                      _18352 };
    assign _18354 = _18353[62:0];
    assign _18362 = { _18354,
                      _18361 };
    assign _18363 = _18362[62:0];
    assign _18371 = { _18363,
                      _18370 };
    assign _18372 = _18371[62:0];
    assign _18380 = { _18372,
                      _18379 };
    assign _18381 = _18380[62:0];
    assign _18389 = { _18381,
                      _18388 };
    assign _18390 = _18389[62:0];
    assign _18398 = { _18390,
                      _18397 };
    assign _18399 = _18398[62:0];
    assign _18407 = { _18399,
                      _18406 };
    assign _18408 = _18407[62:0];
    assign _18416 = { _18408,
                      _18415 };
    assign _18417 = _18416[62:0];
    assign _18425 = { _18417,
                      _18424 };
    assign _18426 = _18425[62:0];
    assign _18434 = { _18426,
                      _18433 };
    assign _18435 = _18434[62:0];
    assign _18443 = { _18435,
                      _18442 };
    assign _18444 = _18443[62:0];
    assign _18452 = { _18444,
                      _18451 };
    assign _18453 = _18452[62:0];
    assign _18461 = { _18453,
                      _18460 };
    assign _18462 = _18461[62:0];
    assign _18470 = { _18462,
                      _18469 };
    assign _18471 = _18470[62:0];
    assign _18479 = { _18471,
                      _18478 };
    assign _18480 = _18479[62:0];
    assign _18488 = { _18480,
                      _18487 };
    assign _18489 = _18488[62:0];
    assign _18497 = { _18489,
                      _18496 };
    assign _18498 = _18497[62:0];
    assign _18506 = { _18498,
                      _18505 };
    assign _18507 = _18506[62:0];
    assign _18515 = { _18507,
                      _18514 };
    assign _18516 = _18515[62:0];
    assign _18524 = { _18516,
                      _18523 };
    assign _18525 = _18524[62:0];
    assign _18533 = { _18525,
                      _18532 };
    assign _18534 = _18533[62:0];
    assign _18542 = { _18534,
                      _18541 };
    assign _18543 = _18542[62:0];
    assign _18551 = { _18543,
                      _18550 };
    assign _18552 = _18551[62:0];
    assign _18560 = { _18552,
                      _18559 };
    assign _18561 = _18560[62:0];
    assign _18569 = { _18561,
                      _18568 };
    assign _18570 = _18569[62:0];
    assign _18578 = { _18570,
                      _18577 };
    assign _18579 = _18578[62:0];
    assign _18587 = { _18579,
                      _18586 };
    assign _18588 = _18587[62:0];
    assign _18596 = { _18588,
                      _18595 };
    assign _18597 = _18596[62:0];
    assign _18605 = { _18597,
                      _18604 };
    assign _18606 = _18605[62:0];
    assign _18614 = { _18606,
                      _18613 };
    assign _18615 = _18614[62:0];
    assign _18623 = { _18615,
                      _18622 };
    assign _18624 = _18623[62:0];
    assign _18632 = { _18624,
                      _18631 };
    assign _18633 = _18632[62:0];
    assign _18641 = { _18633,
                      _18640 };
    assign _18642 = _18641[62:0];
    assign _18650 = { _18642,
                      _18649 };
    assign _18651 = _18650[62:0];
    assign _18659 = { _18651,
                      _18658 };
    assign _18660 = _18659[62:0];
    assign _18668 = { _18660,
                      _18667 };
    assign _18669 = _18668[62:0];
    assign _18677 = { _18669,
                      _18676 };
    assign _18679 = _18677 + _22186;
    assign _18680 = _18679 * _18099;
    assign _18681 = _18680[63:0];
    assign _19263 = _18681 + _19262;
    assign _18091 = _17522[0:0];
    assign _18088 = _18083 - _17525;
    assign _18089 = _18085 ? _18088 : _18083;
    assign _18090 = _18089[62:0];
    assign _18092 = { _18090,
                      _18091 };
    assign _18093 = _18092 < _17525;
    assign _18094 = ~ _18093;
    assign _18082 = _17522[1:1];
    assign _18079 = _18074 - _17525;
    assign _18080 = _18076 ? _18079 : _18074;
    assign _18081 = _18080[62:0];
    assign _18083 = { _18081,
                      _18082 };
    assign _18084 = _18083 < _17525;
    assign _18085 = ~ _18084;
    assign _18073 = _17522[2:2];
    assign _18070 = _18065 - _17525;
    assign _18071 = _18067 ? _18070 : _18065;
    assign _18072 = _18071[62:0];
    assign _18074 = { _18072,
                      _18073 };
    assign _18075 = _18074 < _17525;
    assign _18076 = ~ _18075;
    assign _18064 = _17522[3:3];
    assign _18061 = _18056 - _17525;
    assign _18062 = _18058 ? _18061 : _18056;
    assign _18063 = _18062[62:0];
    assign _18065 = { _18063,
                      _18064 };
    assign _18066 = _18065 < _17525;
    assign _18067 = ~ _18066;
    assign _18055 = _17522[4:4];
    assign _18052 = _18047 - _17525;
    assign _18053 = _18049 ? _18052 : _18047;
    assign _18054 = _18053[62:0];
    assign _18056 = { _18054,
                      _18055 };
    assign _18057 = _18056 < _17525;
    assign _18058 = ~ _18057;
    assign _18046 = _17522[5:5];
    assign _18043 = _18038 - _17525;
    assign _18044 = _18040 ? _18043 : _18038;
    assign _18045 = _18044[62:0];
    assign _18047 = { _18045,
                      _18046 };
    assign _18048 = _18047 < _17525;
    assign _18049 = ~ _18048;
    assign _18037 = _17522[6:6];
    assign _18034 = _18029 - _17525;
    assign _18035 = _18031 ? _18034 : _18029;
    assign _18036 = _18035[62:0];
    assign _18038 = { _18036,
                      _18037 };
    assign _18039 = _18038 < _17525;
    assign _18040 = ~ _18039;
    assign _18028 = _17522[7:7];
    assign _18025 = _18020 - _17525;
    assign _18026 = _18022 ? _18025 : _18020;
    assign _18027 = _18026[62:0];
    assign _18029 = { _18027,
                      _18028 };
    assign _18030 = _18029 < _17525;
    assign _18031 = ~ _18030;
    assign _18019 = _17522[8:8];
    assign _18016 = _18011 - _17525;
    assign _18017 = _18013 ? _18016 : _18011;
    assign _18018 = _18017[62:0];
    assign _18020 = { _18018,
                      _18019 };
    assign _18021 = _18020 < _17525;
    assign _18022 = ~ _18021;
    assign _18010 = _17522[9:9];
    assign _18007 = _18002 - _17525;
    assign _18008 = _18004 ? _18007 : _18002;
    assign _18009 = _18008[62:0];
    assign _18011 = { _18009,
                      _18010 };
    assign _18012 = _18011 < _17525;
    assign _18013 = ~ _18012;
    assign _18001 = _17522[10:10];
    assign _17998 = _17993 - _17525;
    assign _17999 = _17995 ? _17998 : _17993;
    assign _18000 = _17999[62:0];
    assign _18002 = { _18000,
                      _18001 };
    assign _18003 = _18002 < _17525;
    assign _18004 = ~ _18003;
    assign _17992 = _17522[11:11];
    assign _17989 = _17984 - _17525;
    assign _17990 = _17986 ? _17989 : _17984;
    assign _17991 = _17990[62:0];
    assign _17993 = { _17991,
                      _17992 };
    assign _17994 = _17993 < _17525;
    assign _17995 = ~ _17994;
    assign _17983 = _17522[12:12];
    assign _17980 = _17975 - _17525;
    assign _17981 = _17977 ? _17980 : _17975;
    assign _17982 = _17981[62:0];
    assign _17984 = { _17982,
                      _17983 };
    assign _17985 = _17984 < _17525;
    assign _17986 = ~ _17985;
    assign _17974 = _17522[13:13];
    assign _17971 = _17966 - _17525;
    assign _17972 = _17968 ? _17971 : _17966;
    assign _17973 = _17972[62:0];
    assign _17975 = { _17973,
                      _17974 };
    assign _17976 = _17975 < _17525;
    assign _17977 = ~ _17976;
    assign _17965 = _17522[14:14];
    assign _17962 = _17957 - _17525;
    assign _17963 = _17959 ? _17962 : _17957;
    assign _17964 = _17963[62:0];
    assign _17966 = { _17964,
                      _17965 };
    assign _17967 = _17966 < _17525;
    assign _17968 = ~ _17967;
    assign _17956 = _17522[15:15];
    assign _17953 = _17948 - _17525;
    assign _17954 = _17950 ? _17953 : _17948;
    assign _17955 = _17954[62:0];
    assign _17957 = { _17955,
                      _17956 };
    assign _17958 = _17957 < _17525;
    assign _17959 = ~ _17958;
    assign _17947 = _17522[16:16];
    assign _17944 = _17939 - _17525;
    assign _17945 = _17941 ? _17944 : _17939;
    assign _17946 = _17945[62:0];
    assign _17948 = { _17946,
                      _17947 };
    assign _17949 = _17948 < _17525;
    assign _17950 = ~ _17949;
    assign _17938 = _17522[17:17];
    assign _17935 = _17930 - _17525;
    assign _17936 = _17932 ? _17935 : _17930;
    assign _17937 = _17936[62:0];
    assign _17939 = { _17937,
                      _17938 };
    assign _17940 = _17939 < _17525;
    assign _17941 = ~ _17940;
    assign _17929 = _17522[18:18];
    assign _17926 = _17921 - _17525;
    assign _17927 = _17923 ? _17926 : _17921;
    assign _17928 = _17927[62:0];
    assign _17930 = { _17928,
                      _17929 };
    assign _17931 = _17930 < _17525;
    assign _17932 = ~ _17931;
    assign _17920 = _17522[19:19];
    assign _17917 = _17912 - _17525;
    assign _17918 = _17914 ? _17917 : _17912;
    assign _17919 = _17918[62:0];
    assign _17921 = { _17919,
                      _17920 };
    assign _17922 = _17921 < _17525;
    assign _17923 = ~ _17922;
    assign _17911 = _17522[20:20];
    assign _17908 = _17903 - _17525;
    assign _17909 = _17905 ? _17908 : _17903;
    assign _17910 = _17909[62:0];
    assign _17912 = { _17910,
                      _17911 };
    assign _17913 = _17912 < _17525;
    assign _17914 = ~ _17913;
    assign _17902 = _17522[21:21];
    assign _17899 = _17894 - _17525;
    assign _17900 = _17896 ? _17899 : _17894;
    assign _17901 = _17900[62:0];
    assign _17903 = { _17901,
                      _17902 };
    assign _17904 = _17903 < _17525;
    assign _17905 = ~ _17904;
    assign _17893 = _17522[22:22];
    assign _17890 = _17885 - _17525;
    assign _17891 = _17887 ? _17890 : _17885;
    assign _17892 = _17891[62:0];
    assign _17894 = { _17892,
                      _17893 };
    assign _17895 = _17894 < _17525;
    assign _17896 = ~ _17895;
    assign _17884 = _17522[23:23];
    assign _17881 = _17876 - _17525;
    assign _17882 = _17878 ? _17881 : _17876;
    assign _17883 = _17882[62:0];
    assign _17885 = { _17883,
                      _17884 };
    assign _17886 = _17885 < _17525;
    assign _17887 = ~ _17886;
    assign _17875 = _17522[24:24];
    assign _17872 = _17867 - _17525;
    assign _17873 = _17869 ? _17872 : _17867;
    assign _17874 = _17873[62:0];
    assign _17876 = { _17874,
                      _17875 };
    assign _17877 = _17876 < _17525;
    assign _17878 = ~ _17877;
    assign _17866 = _17522[25:25];
    assign _17863 = _17858 - _17525;
    assign _17864 = _17860 ? _17863 : _17858;
    assign _17865 = _17864[62:0];
    assign _17867 = { _17865,
                      _17866 };
    assign _17868 = _17867 < _17525;
    assign _17869 = ~ _17868;
    assign _17857 = _17522[26:26];
    assign _17854 = _17849 - _17525;
    assign _17855 = _17851 ? _17854 : _17849;
    assign _17856 = _17855[62:0];
    assign _17858 = { _17856,
                      _17857 };
    assign _17859 = _17858 < _17525;
    assign _17860 = ~ _17859;
    assign _17848 = _17522[27:27];
    assign _17845 = _17840 - _17525;
    assign _17846 = _17842 ? _17845 : _17840;
    assign _17847 = _17846[62:0];
    assign _17849 = { _17847,
                      _17848 };
    assign _17850 = _17849 < _17525;
    assign _17851 = ~ _17850;
    assign _17839 = _17522[28:28];
    assign _17836 = _17831 - _17525;
    assign _17837 = _17833 ? _17836 : _17831;
    assign _17838 = _17837[62:0];
    assign _17840 = { _17838,
                      _17839 };
    assign _17841 = _17840 < _17525;
    assign _17842 = ~ _17841;
    assign _17830 = _17522[29:29];
    assign _17827 = _17822 - _17525;
    assign _17828 = _17824 ? _17827 : _17822;
    assign _17829 = _17828[62:0];
    assign _17831 = { _17829,
                      _17830 };
    assign _17832 = _17831 < _17525;
    assign _17833 = ~ _17832;
    assign _17821 = _17522[30:30];
    assign _17818 = _17813 - _17525;
    assign _17819 = _17815 ? _17818 : _17813;
    assign _17820 = _17819[62:0];
    assign _17822 = { _17820,
                      _17821 };
    assign _17823 = _17822 < _17525;
    assign _17824 = ~ _17823;
    assign _17812 = _17522[31:31];
    assign _17809 = _17804 - _17525;
    assign _17810 = _17806 ? _17809 : _17804;
    assign _17811 = _17810[62:0];
    assign _17813 = { _17811,
                      _17812 };
    assign _17814 = _17813 < _17525;
    assign _17815 = ~ _17814;
    assign _17803 = _17522[32:32];
    assign _17800 = _17795 - _17525;
    assign _17801 = _17797 ? _17800 : _17795;
    assign _17802 = _17801[62:0];
    assign _17804 = { _17802,
                      _17803 };
    assign _17805 = _17804 < _17525;
    assign _17806 = ~ _17805;
    assign _17794 = _17522[33:33];
    assign _17791 = _17786 - _17525;
    assign _17792 = _17788 ? _17791 : _17786;
    assign _17793 = _17792[62:0];
    assign _17795 = { _17793,
                      _17794 };
    assign _17796 = _17795 < _17525;
    assign _17797 = ~ _17796;
    assign _17785 = _17522[34:34];
    assign _17782 = _17777 - _17525;
    assign _17783 = _17779 ? _17782 : _17777;
    assign _17784 = _17783[62:0];
    assign _17786 = { _17784,
                      _17785 };
    assign _17787 = _17786 < _17525;
    assign _17788 = ~ _17787;
    assign _17776 = _17522[35:35];
    assign _17773 = _17768 - _17525;
    assign _17774 = _17770 ? _17773 : _17768;
    assign _17775 = _17774[62:0];
    assign _17777 = { _17775,
                      _17776 };
    assign _17778 = _17777 < _17525;
    assign _17779 = ~ _17778;
    assign _17767 = _17522[36:36];
    assign _17764 = _17759 - _17525;
    assign _17765 = _17761 ? _17764 : _17759;
    assign _17766 = _17765[62:0];
    assign _17768 = { _17766,
                      _17767 };
    assign _17769 = _17768 < _17525;
    assign _17770 = ~ _17769;
    assign _17758 = _17522[37:37];
    assign _17755 = _17750 - _17525;
    assign _17756 = _17752 ? _17755 : _17750;
    assign _17757 = _17756[62:0];
    assign _17759 = { _17757,
                      _17758 };
    assign _17760 = _17759 < _17525;
    assign _17761 = ~ _17760;
    assign _17749 = _17522[38:38];
    assign _17746 = _17741 - _17525;
    assign _17747 = _17743 ? _17746 : _17741;
    assign _17748 = _17747[62:0];
    assign _17750 = { _17748,
                      _17749 };
    assign _17751 = _17750 < _17525;
    assign _17752 = ~ _17751;
    assign _17740 = _17522[39:39];
    assign _17737 = _17732 - _17525;
    assign _17738 = _17734 ? _17737 : _17732;
    assign _17739 = _17738[62:0];
    assign _17741 = { _17739,
                      _17740 };
    assign _17742 = _17741 < _17525;
    assign _17743 = ~ _17742;
    assign _17731 = _17522[40:40];
    assign _17728 = _17723 - _17525;
    assign _17729 = _17725 ? _17728 : _17723;
    assign _17730 = _17729[62:0];
    assign _17732 = { _17730,
                      _17731 };
    assign _17733 = _17732 < _17525;
    assign _17734 = ~ _17733;
    assign _17722 = _17522[41:41];
    assign _17719 = _17714 - _17525;
    assign _17720 = _17716 ? _17719 : _17714;
    assign _17721 = _17720[62:0];
    assign _17723 = { _17721,
                      _17722 };
    assign _17724 = _17723 < _17525;
    assign _17725 = ~ _17724;
    assign _17713 = _17522[42:42];
    assign _17710 = _17705 - _17525;
    assign _17711 = _17707 ? _17710 : _17705;
    assign _17712 = _17711[62:0];
    assign _17714 = { _17712,
                      _17713 };
    assign _17715 = _17714 < _17525;
    assign _17716 = ~ _17715;
    assign _17704 = _17522[43:43];
    assign _17701 = _17696 - _17525;
    assign _17702 = _17698 ? _17701 : _17696;
    assign _17703 = _17702[62:0];
    assign _17705 = { _17703,
                      _17704 };
    assign _17706 = _17705 < _17525;
    assign _17707 = ~ _17706;
    assign _17695 = _17522[44:44];
    assign _17692 = _17687 - _17525;
    assign _17693 = _17689 ? _17692 : _17687;
    assign _17694 = _17693[62:0];
    assign _17696 = { _17694,
                      _17695 };
    assign _17697 = _17696 < _17525;
    assign _17698 = ~ _17697;
    assign _17686 = _17522[45:45];
    assign _17683 = _17678 - _17525;
    assign _17684 = _17680 ? _17683 : _17678;
    assign _17685 = _17684[62:0];
    assign _17687 = { _17685,
                      _17686 };
    assign _17688 = _17687 < _17525;
    assign _17689 = ~ _17688;
    assign _17677 = _17522[46:46];
    assign _17674 = _17669 - _17525;
    assign _17675 = _17671 ? _17674 : _17669;
    assign _17676 = _17675[62:0];
    assign _17678 = { _17676,
                      _17677 };
    assign _17679 = _17678 < _17525;
    assign _17680 = ~ _17679;
    assign _17668 = _17522[47:47];
    assign _17665 = _17660 - _17525;
    assign _17666 = _17662 ? _17665 : _17660;
    assign _17667 = _17666[62:0];
    assign _17669 = { _17667,
                      _17668 };
    assign _17670 = _17669 < _17525;
    assign _17671 = ~ _17670;
    assign _17659 = _17522[48:48];
    assign _17656 = _17651 - _17525;
    assign _17657 = _17653 ? _17656 : _17651;
    assign _17658 = _17657[62:0];
    assign _17660 = { _17658,
                      _17659 };
    assign _17661 = _17660 < _17525;
    assign _17662 = ~ _17661;
    assign _17650 = _17522[49:49];
    assign _17647 = _17642 - _17525;
    assign _17648 = _17644 ? _17647 : _17642;
    assign _17649 = _17648[62:0];
    assign _17651 = { _17649,
                      _17650 };
    assign _17652 = _17651 < _17525;
    assign _17653 = ~ _17652;
    assign _17641 = _17522[50:50];
    assign _17638 = _17633 - _17525;
    assign _17639 = _17635 ? _17638 : _17633;
    assign _17640 = _17639[62:0];
    assign _17642 = { _17640,
                      _17641 };
    assign _17643 = _17642 < _17525;
    assign _17644 = ~ _17643;
    assign _17632 = _17522[51:51];
    assign _17629 = _17624 - _17525;
    assign _17630 = _17626 ? _17629 : _17624;
    assign _17631 = _17630[62:0];
    assign _17633 = { _17631,
                      _17632 };
    assign _17634 = _17633 < _17525;
    assign _17635 = ~ _17634;
    assign _17623 = _17522[52:52];
    assign _17620 = _17615 - _17525;
    assign _17621 = _17617 ? _17620 : _17615;
    assign _17622 = _17621[62:0];
    assign _17624 = { _17622,
                      _17623 };
    assign _17625 = _17624 < _17525;
    assign _17626 = ~ _17625;
    assign _17614 = _17522[53:53];
    assign _17611 = _17606 - _17525;
    assign _17612 = _17608 ? _17611 : _17606;
    assign _17613 = _17612[62:0];
    assign _17615 = { _17613,
                      _17614 };
    assign _17616 = _17615 < _17525;
    assign _17617 = ~ _17616;
    assign _17605 = _17522[54:54];
    assign _17602 = _17597 - _17525;
    assign _17603 = _17599 ? _17602 : _17597;
    assign _17604 = _17603[62:0];
    assign _17606 = { _17604,
                      _17605 };
    assign _17607 = _17606 < _17525;
    assign _17608 = ~ _17607;
    assign _17596 = _17522[55:55];
    assign _17593 = _17588 - _17525;
    assign _17594 = _17590 ? _17593 : _17588;
    assign _17595 = _17594[62:0];
    assign _17597 = { _17595,
                      _17596 };
    assign _17598 = _17597 < _17525;
    assign _17599 = ~ _17598;
    assign _17587 = _17522[56:56];
    assign _17584 = _17579 - _17525;
    assign _17585 = _17581 ? _17584 : _17579;
    assign _17586 = _17585[62:0];
    assign _17588 = { _17586,
                      _17587 };
    assign _17589 = _17588 < _17525;
    assign _17590 = ~ _17589;
    assign _17578 = _17522[57:57];
    assign _17575 = _17570 - _17525;
    assign _17576 = _17572 ? _17575 : _17570;
    assign _17577 = _17576[62:0];
    assign _17579 = { _17577,
                      _17578 };
    assign _17580 = _17579 < _17525;
    assign _17581 = ~ _17580;
    assign _17569 = _17522[58:58];
    assign _17566 = _17561 - _17525;
    assign _17567 = _17563 ? _17566 : _17561;
    assign _17568 = _17567[62:0];
    assign _17570 = { _17568,
                      _17569 };
    assign _17571 = _17570 < _17525;
    assign _17572 = ~ _17571;
    assign _17560 = _17522[59:59];
    assign _17557 = _17552 - _17525;
    assign _17558 = _17554 ? _17557 : _17552;
    assign _17559 = _17558[62:0];
    assign _17561 = { _17559,
                      _17560 };
    assign _17562 = _17561 < _17525;
    assign _17563 = ~ _17562;
    assign _17551 = _17522[60:60];
    assign _17548 = _17543 - _17525;
    assign _17549 = _17545 ? _17548 : _17543;
    assign _17550 = _17549[62:0];
    assign _17552 = { _17550,
                      _17551 };
    assign _17553 = _17552 < _17525;
    assign _17554 = ~ _17553;
    assign _17542 = _17522[61:61];
    assign _17539 = _17534 - _17525;
    assign _17540 = _17536 ? _17539 : _17534;
    assign _17541 = _17540[62:0];
    assign _17543 = { _17541,
                      _17542 };
    assign _17544 = _17543 < _17525;
    assign _17545 = ~ _17544;
    assign _17533 = _17522[62:62];
    assign _17530 = _17524 - _17525;
    assign _17531 = _17527 ? _17530 : _17524;
    assign _17532 = _17531[62:0];
    assign _17534 = { _17532,
                      _17533 };
    assign _17535 = _17534 < _17525;
    assign _17536 = ~ _17535;
    assign _17525 = 64'b0000000000000000000000000000000000000110000001010100101010110101;
    assign _17521 = 64'b0000000000000000000000000000000000000110000001010100101010110100;
    assign _17522 = _3 + _17521;
    assign _17523 = _17522[63:63];
    assign _17524 = { _22185,
                      _17523 };
    assign _17526 = _17524 < _17525;
    assign _17527 = ~ _17526;
    assign _17528 = { _22185,
                      _17527 };
    assign _17529 = _17528[62:0];
    assign _17537 = { _17529,
                      _17536 };
    assign _17538 = _17537[62:0];
    assign _17546 = { _17538,
                      _17545 };
    assign _17547 = _17546[62:0];
    assign _17555 = { _17547,
                      _17554 };
    assign _17556 = _17555[62:0];
    assign _17564 = { _17556,
                      _17563 };
    assign _17565 = _17564[62:0];
    assign _17573 = { _17565,
                      _17572 };
    assign _17574 = _17573[62:0];
    assign _17582 = { _17574,
                      _17581 };
    assign _17583 = _17582[62:0];
    assign _17591 = { _17583,
                      _17590 };
    assign _17592 = _17591[62:0];
    assign _17600 = { _17592,
                      _17599 };
    assign _17601 = _17600[62:0];
    assign _17609 = { _17601,
                      _17608 };
    assign _17610 = _17609[62:0];
    assign _17618 = { _17610,
                      _17617 };
    assign _17619 = _17618[62:0];
    assign _17627 = { _17619,
                      _17626 };
    assign _17628 = _17627[62:0];
    assign _17636 = { _17628,
                      _17635 };
    assign _17637 = _17636[62:0];
    assign _17645 = { _17637,
                      _17644 };
    assign _17646 = _17645[62:0];
    assign _17654 = { _17646,
                      _17653 };
    assign _17655 = _17654[62:0];
    assign _17663 = { _17655,
                      _17662 };
    assign _17664 = _17663[62:0];
    assign _17672 = { _17664,
                      _17671 };
    assign _17673 = _17672[62:0];
    assign _17681 = { _17673,
                      _17680 };
    assign _17682 = _17681[62:0];
    assign _17690 = { _17682,
                      _17689 };
    assign _17691 = _17690[62:0];
    assign _17699 = { _17691,
                      _17698 };
    assign _17700 = _17699[62:0];
    assign _17708 = { _17700,
                      _17707 };
    assign _17709 = _17708[62:0];
    assign _17717 = { _17709,
                      _17716 };
    assign _17718 = _17717[62:0];
    assign _17726 = { _17718,
                      _17725 };
    assign _17727 = _17726[62:0];
    assign _17735 = { _17727,
                      _17734 };
    assign _17736 = _17735[62:0];
    assign _17744 = { _17736,
                      _17743 };
    assign _17745 = _17744[62:0];
    assign _17753 = { _17745,
                      _17752 };
    assign _17754 = _17753[62:0];
    assign _17762 = { _17754,
                      _17761 };
    assign _17763 = _17762[62:0];
    assign _17771 = { _17763,
                      _17770 };
    assign _17772 = _17771[62:0];
    assign _17780 = { _17772,
                      _17779 };
    assign _17781 = _17780[62:0];
    assign _17789 = { _17781,
                      _17788 };
    assign _17790 = _17789[62:0];
    assign _17798 = { _17790,
                      _17797 };
    assign _17799 = _17798[62:0];
    assign _17807 = { _17799,
                      _17806 };
    assign _17808 = _17807[62:0];
    assign _17816 = { _17808,
                      _17815 };
    assign _17817 = _17816[62:0];
    assign _17825 = { _17817,
                      _17824 };
    assign _17826 = _17825[62:0];
    assign _17834 = { _17826,
                      _17833 };
    assign _17835 = _17834[62:0];
    assign _17843 = { _17835,
                      _17842 };
    assign _17844 = _17843[62:0];
    assign _17852 = { _17844,
                      _17851 };
    assign _17853 = _17852[62:0];
    assign _17861 = { _17853,
                      _17860 };
    assign _17862 = _17861[62:0];
    assign _17870 = { _17862,
                      _17869 };
    assign _17871 = _17870[62:0];
    assign _17879 = { _17871,
                      _17878 };
    assign _17880 = _17879[62:0];
    assign _17888 = { _17880,
                      _17887 };
    assign _17889 = _17888[62:0];
    assign _17897 = { _17889,
                      _17896 };
    assign _17898 = _17897[62:0];
    assign _17906 = { _17898,
                      _17905 };
    assign _17907 = _17906[62:0];
    assign _17915 = { _17907,
                      _17914 };
    assign _17916 = _17915[62:0];
    assign _17924 = { _17916,
                      _17923 };
    assign _17925 = _17924[62:0];
    assign _17933 = { _17925,
                      _17932 };
    assign _17934 = _17933[62:0];
    assign _17942 = { _17934,
                      _17941 };
    assign _17943 = _17942[62:0];
    assign _17951 = { _17943,
                      _17950 };
    assign _17952 = _17951[62:0];
    assign _17960 = { _17952,
                      _17959 };
    assign _17961 = _17960[62:0];
    assign _17969 = { _17961,
                      _17968 };
    assign _17970 = _17969[62:0];
    assign _17978 = { _17970,
                      _17977 };
    assign _17979 = _17978[62:0];
    assign _17987 = { _17979,
                      _17986 };
    assign _17988 = _17987[62:0];
    assign _17996 = { _17988,
                      _17995 };
    assign _17997 = _17996[62:0];
    assign _18005 = { _17997,
                      _18004 };
    assign _18006 = _18005[62:0];
    assign _18014 = { _18006,
                      _18013 };
    assign _18015 = _18014[62:0];
    assign _18023 = { _18015,
                      _18022 };
    assign _18024 = _18023[62:0];
    assign _18032 = { _18024,
                      _18031 };
    assign _18033 = _18032[62:0];
    assign _18041 = { _18033,
                      _18040 };
    assign _18042 = _18041[62:0];
    assign _18050 = { _18042,
                      _18049 };
    assign _18051 = _18050[62:0];
    assign _18059 = { _18051,
                      _18058 };
    assign _18060 = _18059[62:0];
    assign _18068 = { _18060,
                      _18067 };
    assign _18069 = _18068[62:0];
    assign _18077 = { _18069,
                      _18076 };
    assign _18078 = _18077[62:0];
    assign _18086 = { _18078,
                      _18085 };
    assign _18087 = _18086[62:0];
    assign _18095 = { _18087,
                      _18094 };
    assign _18096 = _18095 * _17525;
    assign _18097 = _18096[63:0];
    assign _17518 = 64'b0000000000000000000000000000000000111100001101001110101100010010;
    assign _18098 = _17518 < _18097;
    assign _18099 = _18098 ? _18097 : _17518;
    assign _17516 = _5 < _21017;
    assign _17517 = _17516 ? _5 : _21017;
    assign _18100 = _17517 < _18099;
    assign _18101 = ~ _18100;
    assign _19264 = _18101 ? _19263 : _21604;
    assign _17505 = _16936[0:0];
    assign _17502 = _17497 - _22192;
    assign _17503 = _17499 ? _17502 : _17497;
    assign _17504 = _17503[62:0];
    assign _17506 = { _17504,
                      _17505 };
    assign _17507 = _17506 < _22192;
    assign _17508 = ~ _17507;
    assign _17496 = _16936[1:1];
    assign _17493 = _17488 - _22192;
    assign _17494 = _17490 ? _17493 : _17488;
    assign _17495 = _17494[62:0];
    assign _17497 = { _17495,
                      _17496 };
    assign _17498 = _17497 < _22192;
    assign _17499 = ~ _17498;
    assign _17487 = _16936[2:2];
    assign _17484 = _17479 - _22192;
    assign _17485 = _17481 ? _17484 : _17479;
    assign _17486 = _17485[62:0];
    assign _17488 = { _17486,
                      _17487 };
    assign _17489 = _17488 < _22192;
    assign _17490 = ~ _17489;
    assign _17478 = _16936[3:3];
    assign _17475 = _17470 - _22192;
    assign _17476 = _17472 ? _17475 : _17470;
    assign _17477 = _17476[62:0];
    assign _17479 = { _17477,
                      _17478 };
    assign _17480 = _17479 < _22192;
    assign _17481 = ~ _17480;
    assign _17469 = _16936[4:4];
    assign _17466 = _17461 - _22192;
    assign _17467 = _17463 ? _17466 : _17461;
    assign _17468 = _17467[62:0];
    assign _17470 = { _17468,
                      _17469 };
    assign _17471 = _17470 < _22192;
    assign _17472 = ~ _17471;
    assign _17460 = _16936[5:5];
    assign _17457 = _17452 - _22192;
    assign _17458 = _17454 ? _17457 : _17452;
    assign _17459 = _17458[62:0];
    assign _17461 = { _17459,
                      _17460 };
    assign _17462 = _17461 < _22192;
    assign _17463 = ~ _17462;
    assign _17451 = _16936[6:6];
    assign _17448 = _17443 - _22192;
    assign _17449 = _17445 ? _17448 : _17443;
    assign _17450 = _17449[62:0];
    assign _17452 = { _17450,
                      _17451 };
    assign _17453 = _17452 < _22192;
    assign _17454 = ~ _17453;
    assign _17442 = _16936[7:7];
    assign _17439 = _17434 - _22192;
    assign _17440 = _17436 ? _17439 : _17434;
    assign _17441 = _17440[62:0];
    assign _17443 = { _17441,
                      _17442 };
    assign _17444 = _17443 < _22192;
    assign _17445 = ~ _17444;
    assign _17433 = _16936[8:8];
    assign _17430 = _17425 - _22192;
    assign _17431 = _17427 ? _17430 : _17425;
    assign _17432 = _17431[62:0];
    assign _17434 = { _17432,
                      _17433 };
    assign _17435 = _17434 < _22192;
    assign _17436 = ~ _17435;
    assign _17424 = _16936[9:9];
    assign _17421 = _17416 - _22192;
    assign _17422 = _17418 ? _17421 : _17416;
    assign _17423 = _17422[62:0];
    assign _17425 = { _17423,
                      _17424 };
    assign _17426 = _17425 < _22192;
    assign _17427 = ~ _17426;
    assign _17415 = _16936[10:10];
    assign _17412 = _17407 - _22192;
    assign _17413 = _17409 ? _17412 : _17407;
    assign _17414 = _17413[62:0];
    assign _17416 = { _17414,
                      _17415 };
    assign _17417 = _17416 < _22192;
    assign _17418 = ~ _17417;
    assign _17406 = _16936[11:11];
    assign _17403 = _17398 - _22192;
    assign _17404 = _17400 ? _17403 : _17398;
    assign _17405 = _17404[62:0];
    assign _17407 = { _17405,
                      _17406 };
    assign _17408 = _17407 < _22192;
    assign _17409 = ~ _17408;
    assign _17397 = _16936[12:12];
    assign _17394 = _17389 - _22192;
    assign _17395 = _17391 ? _17394 : _17389;
    assign _17396 = _17395[62:0];
    assign _17398 = { _17396,
                      _17397 };
    assign _17399 = _17398 < _22192;
    assign _17400 = ~ _17399;
    assign _17388 = _16936[13:13];
    assign _17385 = _17380 - _22192;
    assign _17386 = _17382 ? _17385 : _17380;
    assign _17387 = _17386[62:0];
    assign _17389 = { _17387,
                      _17388 };
    assign _17390 = _17389 < _22192;
    assign _17391 = ~ _17390;
    assign _17379 = _16936[14:14];
    assign _17376 = _17371 - _22192;
    assign _17377 = _17373 ? _17376 : _17371;
    assign _17378 = _17377[62:0];
    assign _17380 = { _17378,
                      _17379 };
    assign _17381 = _17380 < _22192;
    assign _17382 = ~ _17381;
    assign _17370 = _16936[15:15];
    assign _17367 = _17362 - _22192;
    assign _17368 = _17364 ? _17367 : _17362;
    assign _17369 = _17368[62:0];
    assign _17371 = { _17369,
                      _17370 };
    assign _17372 = _17371 < _22192;
    assign _17373 = ~ _17372;
    assign _17361 = _16936[16:16];
    assign _17358 = _17353 - _22192;
    assign _17359 = _17355 ? _17358 : _17353;
    assign _17360 = _17359[62:0];
    assign _17362 = { _17360,
                      _17361 };
    assign _17363 = _17362 < _22192;
    assign _17364 = ~ _17363;
    assign _17352 = _16936[17:17];
    assign _17349 = _17344 - _22192;
    assign _17350 = _17346 ? _17349 : _17344;
    assign _17351 = _17350[62:0];
    assign _17353 = { _17351,
                      _17352 };
    assign _17354 = _17353 < _22192;
    assign _17355 = ~ _17354;
    assign _17343 = _16936[18:18];
    assign _17340 = _17335 - _22192;
    assign _17341 = _17337 ? _17340 : _17335;
    assign _17342 = _17341[62:0];
    assign _17344 = { _17342,
                      _17343 };
    assign _17345 = _17344 < _22192;
    assign _17346 = ~ _17345;
    assign _17334 = _16936[19:19];
    assign _17331 = _17326 - _22192;
    assign _17332 = _17328 ? _17331 : _17326;
    assign _17333 = _17332[62:0];
    assign _17335 = { _17333,
                      _17334 };
    assign _17336 = _17335 < _22192;
    assign _17337 = ~ _17336;
    assign _17325 = _16936[20:20];
    assign _17322 = _17317 - _22192;
    assign _17323 = _17319 ? _17322 : _17317;
    assign _17324 = _17323[62:0];
    assign _17326 = { _17324,
                      _17325 };
    assign _17327 = _17326 < _22192;
    assign _17328 = ~ _17327;
    assign _17316 = _16936[21:21];
    assign _17313 = _17308 - _22192;
    assign _17314 = _17310 ? _17313 : _17308;
    assign _17315 = _17314[62:0];
    assign _17317 = { _17315,
                      _17316 };
    assign _17318 = _17317 < _22192;
    assign _17319 = ~ _17318;
    assign _17307 = _16936[22:22];
    assign _17304 = _17299 - _22192;
    assign _17305 = _17301 ? _17304 : _17299;
    assign _17306 = _17305[62:0];
    assign _17308 = { _17306,
                      _17307 };
    assign _17309 = _17308 < _22192;
    assign _17310 = ~ _17309;
    assign _17298 = _16936[23:23];
    assign _17295 = _17290 - _22192;
    assign _17296 = _17292 ? _17295 : _17290;
    assign _17297 = _17296[62:0];
    assign _17299 = { _17297,
                      _17298 };
    assign _17300 = _17299 < _22192;
    assign _17301 = ~ _17300;
    assign _17289 = _16936[24:24];
    assign _17286 = _17281 - _22192;
    assign _17287 = _17283 ? _17286 : _17281;
    assign _17288 = _17287[62:0];
    assign _17290 = { _17288,
                      _17289 };
    assign _17291 = _17290 < _22192;
    assign _17292 = ~ _17291;
    assign _17280 = _16936[25:25];
    assign _17277 = _17272 - _22192;
    assign _17278 = _17274 ? _17277 : _17272;
    assign _17279 = _17278[62:0];
    assign _17281 = { _17279,
                      _17280 };
    assign _17282 = _17281 < _22192;
    assign _17283 = ~ _17282;
    assign _17271 = _16936[26:26];
    assign _17268 = _17263 - _22192;
    assign _17269 = _17265 ? _17268 : _17263;
    assign _17270 = _17269[62:0];
    assign _17272 = { _17270,
                      _17271 };
    assign _17273 = _17272 < _22192;
    assign _17274 = ~ _17273;
    assign _17262 = _16936[27:27];
    assign _17259 = _17254 - _22192;
    assign _17260 = _17256 ? _17259 : _17254;
    assign _17261 = _17260[62:0];
    assign _17263 = { _17261,
                      _17262 };
    assign _17264 = _17263 < _22192;
    assign _17265 = ~ _17264;
    assign _17253 = _16936[28:28];
    assign _17250 = _17245 - _22192;
    assign _17251 = _17247 ? _17250 : _17245;
    assign _17252 = _17251[62:0];
    assign _17254 = { _17252,
                      _17253 };
    assign _17255 = _17254 < _22192;
    assign _17256 = ~ _17255;
    assign _17244 = _16936[29:29];
    assign _17241 = _17236 - _22192;
    assign _17242 = _17238 ? _17241 : _17236;
    assign _17243 = _17242[62:0];
    assign _17245 = { _17243,
                      _17244 };
    assign _17246 = _17245 < _22192;
    assign _17247 = ~ _17246;
    assign _17235 = _16936[30:30];
    assign _17232 = _17227 - _22192;
    assign _17233 = _17229 ? _17232 : _17227;
    assign _17234 = _17233[62:0];
    assign _17236 = { _17234,
                      _17235 };
    assign _17237 = _17236 < _22192;
    assign _17238 = ~ _17237;
    assign _17226 = _16936[31:31];
    assign _17223 = _17218 - _22192;
    assign _17224 = _17220 ? _17223 : _17218;
    assign _17225 = _17224[62:0];
    assign _17227 = { _17225,
                      _17226 };
    assign _17228 = _17227 < _22192;
    assign _17229 = ~ _17228;
    assign _17217 = _16936[32:32];
    assign _17214 = _17209 - _22192;
    assign _17215 = _17211 ? _17214 : _17209;
    assign _17216 = _17215[62:0];
    assign _17218 = { _17216,
                      _17217 };
    assign _17219 = _17218 < _22192;
    assign _17220 = ~ _17219;
    assign _17208 = _16936[33:33];
    assign _17205 = _17200 - _22192;
    assign _17206 = _17202 ? _17205 : _17200;
    assign _17207 = _17206[62:0];
    assign _17209 = { _17207,
                      _17208 };
    assign _17210 = _17209 < _22192;
    assign _17211 = ~ _17210;
    assign _17199 = _16936[34:34];
    assign _17196 = _17191 - _22192;
    assign _17197 = _17193 ? _17196 : _17191;
    assign _17198 = _17197[62:0];
    assign _17200 = { _17198,
                      _17199 };
    assign _17201 = _17200 < _22192;
    assign _17202 = ~ _17201;
    assign _17190 = _16936[35:35];
    assign _17187 = _17182 - _22192;
    assign _17188 = _17184 ? _17187 : _17182;
    assign _17189 = _17188[62:0];
    assign _17191 = { _17189,
                      _17190 };
    assign _17192 = _17191 < _22192;
    assign _17193 = ~ _17192;
    assign _17181 = _16936[36:36];
    assign _17178 = _17173 - _22192;
    assign _17179 = _17175 ? _17178 : _17173;
    assign _17180 = _17179[62:0];
    assign _17182 = { _17180,
                      _17181 };
    assign _17183 = _17182 < _22192;
    assign _17184 = ~ _17183;
    assign _17172 = _16936[37:37];
    assign _17169 = _17164 - _22192;
    assign _17170 = _17166 ? _17169 : _17164;
    assign _17171 = _17170[62:0];
    assign _17173 = { _17171,
                      _17172 };
    assign _17174 = _17173 < _22192;
    assign _17175 = ~ _17174;
    assign _17163 = _16936[38:38];
    assign _17160 = _17155 - _22192;
    assign _17161 = _17157 ? _17160 : _17155;
    assign _17162 = _17161[62:0];
    assign _17164 = { _17162,
                      _17163 };
    assign _17165 = _17164 < _22192;
    assign _17166 = ~ _17165;
    assign _17154 = _16936[39:39];
    assign _17151 = _17146 - _22192;
    assign _17152 = _17148 ? _17151 : _17146;
    assign _17153 = _17152[62:0];
    assign _17155 = { _17153,
                      _17154 };
    assign _17156 = _17155 < _22192;
    assign _17157 = ~ _17156;
    assign _17145 = _16936[40:40];
    assign _17142 = _17137 - _22192;
    assign _17143 = _17139 ? _17142 : _17137;
    assign _17144 = _17143[62:0];
    assign _17146 = { _17144,
                      _17145 };
    assign _17147 = _17146 < _22192;
    assign _17148 = ~ _17147;
    assign _17136 = _16936[41:41];
    assign _17133 = _17128 - _22192;
    assign _17134 = _17130 ? _17133 : _17128;
    assign _17135 = _17134[62:0];
    assign _17137 = { _17135,
                      _17136 };
    assign _17138 = _17137 < _22192;
    assign _17139 = ~ _17138;
    assign _17127 = _16936[42:42];
    assign _17124 = _17119 - _22192;
    assign _17125 = _17121 ? _17124 : _17119;
    assign _17126 = _17125[62:0];
    assign _17128 = { _17126,
                      _17127 };
    assign _17129 = _17128 < _22192;
    assign _17130 = ~ _17129;
    assign _17118 = _16936[43:43];
    assign _17115 = _17110 - _22192;
    assign _17116 = _17112 ? _17115 : _17110;
    assign _17117 = _17116[62:0];
    assign _17119 = { _17117,
                      _17118 };
    assign _17120 = _17119 < _22192;
    assign _17121 = ~ _17120;
    assign _17109 = _16936[44:44];
    assign _17106 = _17101 - _22192;
    assign _17107 = _17103 ? _17106 : _17101;
    assign _17108 = _17107[62:0];
    assign _17110 = { _17108,
                      _17109 };
    assign _17111 = _17110 < _22192;
    assign _17112 = ~ _17111;
    assign _17100 = _16936[45:45];
    assign _17097 = _17092 - _22192;
    assign _17098 = _17094 ? _17097 : _17092;
    assign _17099 = _17098[62:0];
    assign _17101 = { _17099,
                      _17100 };
    assign _17102 = _17101 < _22192;
    assign _17103 = ~ _17102;
    assign _17091 = _16936[46:46];
    assign _17088 = _17083 - _22192;
    assign _17089 = _17085 ? _17088 : _17083;
    assign _17090 = _17089[62:0];
    assign _17092 = { _17090,
                      _17091 };
    assign _17093 = _17092 < _22192;
    assign _17094 = ~ _17093;
    assign _17082 = _16936[47:47];
    assign _17079 = _17074 - _22192;
    assign _17080 = _17076 ? _17079 : _17074;
    assign _17081 = _17080[62:0];
    assign _17083 = { _17081,
                      _17082 };
    assign _17084 = _17083 < _22192;
    assign _17085 = ~ _17084;
    assign _17073 = _16936[48:48];
    assign _17070 = _17065 - _22192;
    assign _17071 = _17067 ? _17070 : _17065;
    assign _17072 = _17071[62:0];
    assign _17074 = { _17072,
                      _17073 };
    assign _17075 = _17074 < _22192;
    assign _17076 = ~ _17075;
    assign _17064 = _16936[49:49];
    assign _17061 = _17056 - _22192;
    assign _17062 = _17058 ? _17061 : _17056;
    assign _17063 = _17062[62:0];
    assign _17065 = { _17063,
                      _17064 };
    assign _17066 = _17065 < _22192;
    assign _17067 = ~ _17066;
    assign _17055 = _16936[50:50];
    assign _17052 = _17047 - _22192;
    assign _17053 = _17049 ? _17052 : _17047;
    assign _17054 = _17053[62:0];
    assign _17056 = { _17054,
                      _17055 };
    assign _17057 = _17056 < _22192;
    assign _17058 = ~ _17057;
    assign _17046 = _16936[51:51];
    assign _17043 = _17038 - _22192;
    assign _17044 = _17040 ? _17043 : _17038;
    assign _17045 = _17044[62:0];
    assign _17047 = { _17045,
                      _17046 };
    assign _17048 = _17047 < _22192;
    assign _17049 = ~ _17048;
    assign _17037 = _16936[52:52];
    assign _17034 = _17029 - _22192;
    assign _17035 = _17031 ? _17034 : _17029;
    assign _17036 = _17035[62:0];
    assign _17038 = { _17036,
                      _17037 };
    assign _17039 = _17038 < _22192;
    assign _17040 = ~ _17039;
    assign _17028 = _16936[53:53];
    assign _17025 = _17020 - _22192;
    assign _17026 = _17022 ? _17025 : _17020;
    assign _17027 = _17026[62:0];
    assign _17029 = { _17027,
                      _17028 };
    assign _17030 = _17029 < _22192;
    assign _17031 = ~ _17030;
    assign _17019 = _16936[54:54];
    assign _17016 = _17011 - _22192;
    assign _17017 = _17013 ? _17016 : _17011;
    assign _17018 = _17017[62:0];
    assign _17020 = { _17018,
                      _17019 };
    assign _17021 = _17020 < _22192;
    assign _17022 = ~ _17021;
    assign _17010 = _16936[55:55];
    assign _17007 = _17002 - _22192;
    assign _17008 = _17004 ? _17007 : _17002;
    assign _17009 = _17008[62:0];
    assign _17011 = { _17009,
                      _17010 };
    assign _17012 = _17011 < _22192;
    assign _17013 = ~ _17012;
    assign _17001 = _16936[56:56];
    assign _16998 = _16993 - _22192;
    assign _16999 = _16995 ? _16998 : _16993;
    assign _17000 = _16999[62:0];
    assign _17002 = { _17000,
                      _17001 };
    assign _17003 = _17002 < _22192;
    assign _17004 = ~ _17003;
    assign _16992 = _16936[57:57];
    assign _16989 = _16984 - _22192;
    assign _16990 = _16986 ? _16989 : _16984;
    assign _16991 = _16990[62:0];
    assign _16993 = { _16991,
                      _16992 };
    assign _16994 = _16993 < _22192;
    assign _16995 = ~ _16994;
    assign _16983 = _16936[58:58];
    assign _16980 = _16975 - _22192;
    assign _16981 = _16977 ? _16980 : _16975;
    assign _16982 = _16981[62:0];
    assign _16984 = { _16982,
                      _16983 };
    assign _16985 = _16984 < _22192;
    assign _16986 = ~ _16985;
    assign _16974 = _16936[59:59];
    assign _16971 = _16966 - _22192;
    assign _16972 = _16968 ? _16971 : _16966;
    assign _16973 = _16972[62:0];
    assign _16975 = { _16973,
                      _16974 };
    assign _16976 = _16975 < _22192;
    assign _16977 = ~ _16976;
    assign _16965 = _16936[60:60];
    assign _16962 = _16957 - _22192;
    assign _16963 = _16959 ? _16962 : _16957;
    assign _16964 = _16963[62:0];
    assign _16966 = { _16964,
                      _16965 };
    assign _16967 = _16966 < _22192;
    assign _16968 = ~ _16967;
    assign _16956 = _16936[61:61];
    assign _16953 = _16948 - _22192;
    assign _16954 = _16950 ? _16953 : _16948;
    assign _16955 = _16954[62:0];
    assign _16957 = { _16955,
                      _16956 };
    assign _16958 = _16957 < _22192;
    assign _16959 = ~ _16958;
    assign _16947 = _16936[62:62];
    assign _16944 = _16938 - _22192;
    assign _16945 = _16941 ? _16944 : _16938;
    assign _16946 = _16945[62:0];
    assign _16948 = { _16946,
                      _16947 };
    assign _16949 = _16948 < _22192;
    assign _16950 = ~ _16949;
    assign _16934 = _16926 + _22186;
    assign _16935 = _16926 * _16934;
    assign _16936 = _16935[63:0];
    assign _16937 = _16936[63:63];
    assign _16938 = { _22185,
                      _16937 };
    assign _16940 = _16938 < _22192;
    assign _16941 = ~ _16940;
    assign _16942 = { _22185,
                      _16941 };
    assign _16943 = _16942[62:0];
    assign _16951 = { _16943,
                      _16950 };
    assign _16952 = _16951[62:0];
    assign _16960 = { _16952,
                      _16959 };
    assign _16961 = _16960[62:0];
    assign _16969 = { _16961,
                      _16968 };
    assign _16970 = _16969[62:0];
    assign _16978 = { _16970,
                      _16977 };
    assign _16979 = _16978[62:0];
    assign _16987 = { _16979,
                      _16986 };
    assign _16988 = _16987[62:0];
    assign _16996 = { _16988,
                      _16995 };
    assign _16997 = _16996[62:0];
    assign _17005 = { _16997,
                      _17004 };
    assign _17006 = _17005[62:0];
    assign _17014 = { _17006,
                      _17013 };
    assign _17015 = _17014[62:0];
    assign _17023 = { _17015,
                      _17022 };
    assign _17024 = _17023[62:0];
    assign _17032 = { _17024,
                      _17031 };
    assign _17033 = _17032[62:0];
    assign _17041 = { _17033,
                      _17040 };
    assign _17042 = _17041[62:0];
    assign _17050 = { _17042,
                      _17049 };
    assign _17051 = _17050[62:0];
    assign _17059 = { _17051,
                      _17058 };
    assign _17060 = _17059[62:0];
    assign _17068 = { _17060,
                      _17067 };
    assign _17069 = _17068[62:0];
    assign _17077 = { _17069,
                      _17076 };
    assign _17078 = _17077[62:0];
    assign _17086 = { _17078,
                      _17085 };
    assign _17087 = _17086[62:0];
    assign _17095 = { _17087,
                      _17094 };
    assign _17096 = _17095[62:0];
    assign _17104 = { _17096,
                      _17103 };
    assign _17105 = _17104[62:0];
    assign _17113 = { _17105,
                      _17112 };
    assign _17114 = _17113[62:0];
    assign _17122 = { _17114,
                      _17121 };
    assign _17123 = _17122[62:0];
    assign _17131 = { _17123,
                      _17130 };
    assign _17132 = _17131[62:0];
    assign _17140 = { _17132,
                      _17139 };
    assign _17141 = _17140[62:0];
    assign _17149 = { _17141,
                      _17148 };
    assign _17150 = _17149[62:0];
    assign _17158 = { _17150,
                      _17157 };
    assign _17159 = _17158[62:0];
    assign _17167 = { _17159,
                      _17166 };
    assign _17168 = _17167[62:0];
    assign _17176 = { _17168,
                      _17175 };
    assign _17177 = _17176[62:0];
    assign _17185 = { _17177,
                      _17184 };
    assign _17186 = _17185[62:0];
    assign _17194 = { _17186,
                      _17193 };
    assign _17195 = _17194[62:0];
    assign _17203 = { _17195,
                      _17202 };
    assign _17204 = _17203[62:0];
    assign _17212 = { _17204,
                      _17211 };
    assign _17213 = _17212[62:0];
    assign _17221 = { _17213,
                      _17220 };
    assign _17222 = _17221[62:0];
    assign _17230 = { _17222,
                      _17229 };
    assign _17231 = _17230[62:0];
    assign _17239 = { _17231,
                      _17238 };
    assign _17240 = _17239[62:0];
    assign _17248 = { _17240,
                      _17247 };
    assign _17249 = _17248[62:0];
    assign _17257 = { _17249,
                      _17256 };
    assign _17258 = _17257[62:0];
    assign _17266 = { _17258,
                      _17265 };
    assign _17267 = _17266[62:0];
    assign _17275 = { _17267,
                      _17274 };
    assign _17276 = _17275[62:0];
    assign _17284 = { _17276,
                      _17283 };
    assign _17285 = _17284[62:0];
    assign _17293 = { _17285,
                      _17292 };
    assign _17294 = _17293[62:0];
    assign _17302 = { _17294,
                      _17301 };
    assign _17303 = _17302[62:0];
    assign _17311 = { _17303,
                      _17310 };
    assign _17312 = _17311[62:0];
    assign _17320 = { _17312,
                      _17319 };
    assign _17321 = _17320[62:0];
    assign _17329 = { _17321,
                      _17328 };
    assign _17330 = _17329[62:0];
    assign _17338 = { _17330,
                      _17337 };
    assign _17339 = _17338[62:0];
    assign _17347 = { _17339,
                      _17346 };
    assign _17348 = _17347[62:0];
    assign _17356 = { _17348,
                      _17355 };
    assign _17357 = _17356[62:0];
    assign _17365 = { _17357,
                      _17364 };
    assign _17366 = _17365[62:0];
    assign _17374 = { _17366,
                      _17373 };
    assign _17375 = _17374[62:0];
    assign _17383 = { _17375,
                      _17382 };
    assign _17384 = _17383[62:0];
    assign _17392 = { _17384,
                      _17391 };
    assign _17393 = _17392[62:0];
    assign _17401 = { _17393,
                      _17400 };
    assign _17402 = _17401[62:0];
    assign _17410 = { _17402,
                      _17409 };
    assign _17411 = _17410[62:0];
    assign _17419 = { _17411,
                      _17418 };
    assign _17420 = _17419[62:0];
    assign _17428 = { _17420,
                      _17427 };
    assign _17429 = _17428[62:0];
    assign _17437 = { _17429,
                      _17436 };
    assign _17438 = _17437[62:0];
    assign _17446 = { _17438,
                      _17445 };
    assign _17447 = _17446[62:0];
    assign _17455 = { _17447,
                      _17454 };
    assign _17456 = _17455[62:0];
    assign _17464 = { _17456,
                      _17463 };
    assign _17465 = _17464[62:0];
    assign _17473 = { _17465,
                      _17472 };
    assign _17474 = _17473[62:0];
    assign _17482 = { _17474,
                      _17481 };
    assign _17483 = _17482[62:0];
    assign _17491 = { _17483,
                      _17490 };
    assign _17492 = _17491[62:0];
    assign _17500 = { _17492,
                      _17499 };
    assign _17501 = _17500[62:0];
    assign _17509 = { _17501,
                      _17508 };
    assign _17510 = _15774 * _17509;
    assign _17511 = _17510[63:0];
    assign _16922 = _16354[0:0];
    assign _16919 = _16914 - _15774;
    assign _16920 = _16916 ? _16919 : _16914;
    assign _16921 = _16920[62:0];
    assign _16923 = { _16921,
                      _16922 };
    assign _16924 = _16923 < _15774;
    assign _16925 = ~ _16924;
    assign _16913 = _16354[1:1];
    assign _16910 = _16905 - _15774;
    assign _16911 = _16907 ? _16910 : _16905;
    assign _16912 = _16911[62:0];
    assign _16914 = { _16912,
                      _16913 };
    assign _16915 = _16914 < _15774;
    assign _16916 = ~ _16915;
    assign _16904 = _16354[2:2];
    assign _16901 = _16896 - _15774;
    assign _16902 = _16898 ? _16901 : _16896;
    assign _16903 = _16902[62:0];
    assign _16905 = { _16903,
                      _16904 };
    assign _16906 = _16905 < _15774;
    assign _16907 = ~ _16906;
    assign _16895 = _16354[3:3];
    assign _16892 = _16887 - _15774;
    assign _16893 = _16889 ? _16892 : _16887;
    assign _16894 = _16893[62:0];
    assign _16896 = { _16894,
                      _16895 };
    assign _16897 = _16896 < _15774;
    assign _16898 = ~ _16897;
    assign _16886 = _16354[4:4];
    assign _16883 = _16878 - _15774;
    assign _16884 = _16880 ? _16883 : _16878;
    assign _16885 = _16884[62:0];
    assign _16887 = { _16885,
                      _16886 };
    assign _16888 = _16887 < _15774;
    assign _16889 = ~ _16888;
    assign _16877 = _16354[5:5];
    assign _16874 = _16869 - _15774;
    assign _16875 = _16871 ? _16874 : _16869;
    assign _16876 = _16875[62:0];
    assign _16878 = { _16876,
                      _16877 };
    assign _16879 = _16878 < _15774;
    assign _16880 = ~ _16879;
    assign _16868 = _16354[6:6];
    assign _16865 = _16860 - _15774;
    assign _16866 = _16862 ? _16865 : _16860;
    assign _16867 = _16866[62:0];
    assign _16869 = { _16867,
                      _16868 };
    assign _16870 = _16869 < _15774;
    assign _16871 = ~ _16870;
    assign _16859 = _16354[7:7];
    assign _16856 = _16851 - _15774;
    assign _16857 = _16853 ? _16856 : _16851;
    assign _16858 = _16857[62:0];
    assign _16860 = { _16858,
                      _16859 };
    assign _16861 = _16860 < _15774;
    assign _16862 = ~ _16861;
    assign _16850 = _16354[8:8];
    assign _16847 = _16842 - _15774;
    assign _16848 = _16844 ? _16847 : _16842;
    assign _16849 = _16848[62:0];
    assign _16851 = { _16849,
                      _16850 };
    assign _16852 = _16851 < _15774;
    assign _16853 = ~ _16852;
    assign _16841 = _16354[9:9];
    assign _16838 = _16833 - _15774;
    assign _16839 = _16835 ? _16838 : _16833;
    assign _16840 = _16839[62:0];
    assign _16842 = { _16840,
                      _16841 };
    assign _16843 = _16842 < _15774;
    assign _16844 = ~ _16843;
    assign _16832 = _16354[10:10];
    assign _16829 = _16824 - _15774;
    assign _16830 = _16826 ? _16829 : _16824;
    assign _16831 = _16830[62:0];
    assign _16833 = { _16831,
                      _16832 };
    assign _16834 = _16833 < _15774;
    assign _16835 = ~ _16834;
    assign _16823 = _16354[11:11];
    assign _16820 = _16815 - _15774;
    assign _16821 = _16817 ? _16820 : _16815;
    assign _16822 = _16821[62:0];
    assign _16824 = { _16822,
                      _16823 };
    assign _16825 = _16824 < _15774;
    assign _16826 = ~ _16825;
    assign _16814 = _16354[12:12];
    assign _16811 = _16806 - _15774;
    assign _16812 = _16808 ? _16811 : _16806;
    assign _16813 = _16812[62:0];
    assign _16815 = { _16813,
                      _16814 };
    assign _16816 = _16815 < _15774;
    assign _16817 = ~ _16816;
    assign _16805 = _16354[13:13];
    assign _16802 = _16797 - _15774;
    assign _16803 = _16799 ? _16802 : _16797;
    assign _16804 = _16803[62:0];
    assign _16806 = { _16804,
                      _16805 };
    assign _16807 = _16806 < _15774;
    assign _16808 = ~ _16807;
    assign _16796 = _16354[14:14];
    assign _16793 = _16788 - _15774;
    assign _16794 = _16790 ? _16793 : _16788;
    assign _16795 = _16794[62:0];
    assign _16797 = { _16795,
                      _16796 };
    assign _16798 = _16797 < _15774;
    assign _16799 = ~ _16798;
    assign _16787 = _16354[15:15];
    assign _16784 = _16779 - _15774;
    assign _16785 = _16781 ? _16784 : _16779;
    assign _16786 = _16785[62:0];
    assign _16788 = { _16786,
                      _16787 };
    assign _16789 = _16788 < _15774;
    assign _16790 = ~ _16789;
    assign _16778 = _16354[16:16];
    assign _16775 = _16770 - _15774;
    assign _16776 = _16772 ? _16775 : _16770;
    assign _16777 = _16776[62:0];
    assign _16779 = { _16777,
                      _16778 };
    assign _16780 = _16779 < _15774;
    assign _16781 = ~ _16780;
    assign _16769 = _16354[17:17];
    assign _16766 = _16761 - _15774;
    assign _16767 = _16763 ? _16766 : _16761;
    assign _16768 = _16767[62:0];
    assign _16770 = { _16768,
                      _16769 };
    assign _16771 = _16770 < _15774;
    assign _16772 = ~ _16771;
    assign _16760 = _16354[18:18];
    assign _16757 = _16752 - _15774;
    assign _16758 = _16754 ? _16757 : _16752;
    assign _16759 = _16758[62:0];
    assign _16761 = { _16759,
                      _16760 };
    assign _16762 = _16761 < _15774;
    assign _16763 = ~ _16762;
    assign _16751 = _16354[19:19];
    assign _16748 = _16743 - _15774;
    assign _16749 = _16745 ? _16748 : _16743;
    assign _16750 = _16749[62:0];
    assign _16752 = { _16750,
                      _16751 };
    assign _16753 = _16752 < _15774;
    assign _16754 = ~ _16753;
    assign _16742 = _16354[20:20];
    assign _16739 = _16734 - _15774;
    assign _16740 = _16736 ? _16739 : _16734;
    assign _16741 = _16740[62:0];
    assign _16743 = { _16741,
                      _16742 };
    assign _16744 = _16743 < _15774;
    assign _16745 = ~ _16744;
    assign _16733 = _16354[21:21];
    assign _16730 = _16725 - _15774;
    assign _16731 = _16727 ? _16730 : _16725;
    assign _16732 = _16731[62:0];
    assign _16734 = { _16732,
                      _16733 };
    assign _16735 = _16734 < _15774;
    assign _16736 = ~ _16735;
    assign _16724 = _16354[22:22];
    assign _16721 = _16716 - _15774;
    assign _16722 = _16718 ? _16721 : _16716;
    assign _16723 = _16722[62:0];
    assign _16725 = { _16723,
                      _16724 };
    assign _16726 = _16725 < _15774;
    assign _16727 = ~ _16726;
    assign _16715 = _16354[23:23];
    assign _16712 = _16707 - _15774;
    assign _16713 = _16709 ? _16712 : _16707;
    assign _16714 = _16713[62:0];
    assign _16716 = { _16714,
                      _16715 };
    assign _16717 = _16716 < _15774;
    assign _16718 = ~ _16717;
    assign _16706 = _16354[24:24];
    assign _16703 = _16698 - _15774;
    assign _16704 = _16700 ? _16703 : _16698;
    assign _16705 = _16704[62:0];
    assign _16707 = { _16705,
                      _16706 };
    assign _16708 = _16707 < _15774;
    assign _16709 = ~ _16708;
    assign _16697 = _16354[25:25];
    assign _16694 = _16689 - _15774;
    assign _16695 = _16691 ? _16694 : _16689;
    assign _16696 = _16695[62:0];
    assign _16698 = { _16696,
                      _16697 };
    assign _16699 = _16698 < _15774;
    assign _16700 = ~ _16699;
    assign _16688 = _16354[26:26];
    assign _16685 = _16680 - _15774;
    assign _16686 = _16682 ? _16685 : _16680;
    assign _16687 = _16686[62:0];
    assign _16689 = { _16687,
                      _16688 };
    assign _16690 = _16689 < _15774;
    assign _16691 = ~ _16690;
    assign _16679 = _16354[27:27];
    assign _16676 = _16671 - _15774;
    assign _16677 = _16673 ? _16676 : _16671;
    assign _16678 = _16677[62:0];
    assign _16680 = { _16678,
                      _16679 };
    assign _16681 = _16680 < _15774;
    assign _16682 = ~ _16681;
    assign _16670 = _16354[28:28];
    assign _16667 = _16662 - _15774;
    assign _16668 = _16664 ? _16667 : _16662;
    assign _16669 = _16668[62:0];
    assign _16671 = { _16669,
                      _16670 };
    assign _16672 = _16671 < _15774;
    assign _16673 = ~ _16672;
    assign _16661 = _16354[29:29];
    assign _16658 = _16653 - _15774;
    assign _16659 = _16655 ? _16658 : _16653;
    assign _16660 = _16659[62:0];
    assign _16662 = { _16660,
                      _16661 };
    assign _16663 = _16662 < _15774;
    assign _16664 = ~ _16663;
    assign _16652 = _16354[30:30];
    assign _16649 = _16644 - _15774;
    assign _16650 = _16646 ? _16649 : _16644;
    assign _16651 = _16650[62:0];
    assign _16653 = { _16651,
                      _16652 };
    assign _16654 = _16653 < _15774;
    assign _16655 = ~ _16654;
    assign _16643 = _16354[31:31];
    assign _16640 = _16635 - _15774;
    assign _16641 = _16637 ? _16640 : _16635;
    assign _16642 = _16641[62:0];
    assign _16644 = { _16642,
                      _16643 };
    assign _16645 = _16644 < _15774;
    assign _16646 = ~ _16645;
    assign _16634 = _16354[32:32];
    assign _16631 = _16626 - _15774;
    assign _16632 = _16628 ? _16631 : _16626;
    assign _16633 = _16632[62:0];
    assign _16635 = { _16633,
                      _16634 };
    assign _16636 = _16635 < _15774;
    assign _16637 = ~ _16636;
    assign _16625 = _16354[33:33];
    assign _16622 = _16617 - _15774;
    assign _16623 = _16619 ? _16622 : _16617;
    assign _16624 = _16623[62:0];
    assign _16626 = { _16624,
                      _16625 };
    assign _16627 = _16626 < _15774;
    assign _16628 = ~ _16627;
    assign _16616 = _16354[34:34];
    assign _16613 = _16608 - _15774;
    assign _16614 = _16610 ? _16613 : _16608;
    assign _16615 = _16614[62:0];
    assign _16617 = { _16615,
                      _16616 };
    assign _16618 = _16617 < _15774;
    assign _16619 = ~ _16618;
    assign _16607 = _16354[35:35];
    assign _16604 = _16599 - _15774;
    assign _16605 = _16601 ? _16604 : _16599;
    assign _16606 = _16605[62:0];
    assign _16608 = { _16606,
                      _16607 };
    assign _16609 = _16608 < _15774;
    assign _16610 = ~ _16609;
    assign _16598 = _16354[36:36];
    assign _16595 = _16590 - _15774;
    assign _16596 = _16592 ? _16595 : _16590;
    assign _16597 = _16596[62:0];
    assign _16599 = { _16597,
                      _16598 };
    assign _16600 = _16599 < _15774;
    assign _16601 = ~ _16600;
    assign _16589 = _16354[37:37];
    assign _16586 = _16581 - _15774;
    assign _16587 = _16583 ? _16586 : _16581;
    assign _16588 = _16587[62:0];
    assign _16590 = { _16588,
                      _16589 };
    assign _16591 = _16590 < _15774;
    assign _16592 = ~ _16591;
    assign _16580 = _16354[38:38];
    assign _16577 = _16572 - _15774;
    assign _16578 = _16574 ? _16577 : _16572;
    assign _16579 = _16578[62:0];
    assign _16581 = { _16579,
                      _16580 };
    assign _16582 = _16581 < _15774;
    assign _16583 = ~ _16582;
    assign _16571 = _16354[39:39];
    assign _16568 = _16563 - _15774;
    assign _16569 = _16565 ? _16568 : _16563;
    assign _16570 = _16569[62:0];
    assign _16572 = { _16570,
                      _16571 };
    assign _16573 = _16572 < _15774;
    assign _16574 = ~ _16573;
    assign _16562 = _16354[40:40];
    assign _16559 = _16554 - _15774;
    assign _16560 = _16556 ? _16559 : _16554;
    assign _16561 = _16560[62:0];
    assign _16563 = { _16561,
                      _16562 };
    assign _16564 = _16563 < _15774;
    assign _16565 = ~ _16564;
    assign _16553 = _16354[41:41];
    assign _16550 = _16545 - _15774;
    assign _16551 = _16547 ? _16550 : _16545;
    assign _16552 = _16551[62:0];
    assign _16554 = { _16552,
                      _16553 };
    assign _16555 = _16554 < _15774;
    assign _16556 = ~ _16555;
    assign _16544 = _16354[42:42];
    assign _16541 = _16536 - _15774;
    assign _16542 = _16538 ? _16541 : _16536;
    assign _16543 = _16542[62:0];
    assign _16545 = { _16543,
                      _16544 };
    assign _16546 = _16545 < _15774;
    assign _16547 = ~ _16546;
    assign _16535 = _16354[43:43];
    assign _16532 = _16527 - _15774;
    assign _16533 = _16529 ? _16532 : _16527;
    assign _16534 = _16533[62:0];
    assign _16536 = { _16534,
                      _16535 };
    assign _16537 = _16536 < _15774;
    assign _16538 = ~ _16537;
    assign _16526 = _16354[44:44];
    assign _16523 = _16518 - _15774;
    assign _16524 = _16520 ? _16523 : _16518;
    assign _16525 = _16524[62:0];
    assign _16527 = { _16525,
                      _16526 };
    assign _16528 = _16527 < _15774;
    assign _16529 = ~ _16528;
    assign _16517 = _16354[45:45];
    assign _16514 = _16509 - _15774;
    assign _16515 = _16511 ? _16514 : _16509;
    assign _16516 = _16515[62:0];
    assign _16518 = { _16516,
                      _16517 };
    assign _16519 = _16518 < _15774;
    assign _16520 = ~ _16519;
    assign _16508 = _16354[46:46];
    assign _16505 = _16500 - _15774;
    assign _16506 = _16502 ? _16505 : _16500;
    assign _16507 = _16506[62:0];
    assign _16509 = { _16507,
                      _16508 };
    assign _16510 = _16509 < _15774;
    assign _16511 = ~ _16510;
    assign _16499 = _16354[47:47];
    assign _16496 = _16491 - _15774;
    assign _16497 = _16493 ? _16496 : _16491;
    assign _16498 = _16497[62:0];
    assign _16500 = { _16498,
                      _16499 };
    assign _16501 = _16500 < _15774;
    assign _16502 = ~ _16501;
    assign _16490 = _16354[48:48];
    assign _16487 = _16482 - _15774;
    assign _16488 = _16484 ? _16487 : _16482;
    assign _16489 = _16488[62:0];
    assign _16491 = { _16489,
                      _16490 };
    assign _16492 = _16491 < _15774;
    assign _16493 = ~ _16492;
    assign _16481 = _16354[49:49];
    assign _16478 = _16473 - _15774;
    assign _16479 = _16475 ? _16478 : _16473;
    assign _16480 = _16479[62:0];
    assign _16482 = { _16480,
                      _16481 };
    assign _16483 = _16482 < _15774;
    assign _16484 = ~ _16483;
    assign _16472 = _16354[50:50];
    assign _16469 = _16464 - _15774;
    assign _16470 = _16466 ? _16469 : _16464;
    assign _16471 = _16470[62:0];
    assign _16473 = { _16471,
                      _16472 };
    assign _16474 = _16473 < _15774;
    assign _16475 = ~ _16474;
    assign _16463 = _16354[51:51];
    assign _16460 = _16455 - _15774;
    assign _16461 = _16457 ? _16460 : _16455;
    assign _16462 = _16461[62:0];
    assign _16464 = { _16462,
                      _16463 };
    assign _16465 = _16464 < _15774;
    assign _16466 = ~ _16465;
    assign _16454 = _16354[52:52];
    assign _16451 = _16446 - _15774;
    assign _16452 = _16448 ? _16451 : _16446;
    assign _16453 = _16452[62:0];
    assign _16455 = { _16453,
                      _16454 };
    assign _16456 = _16455 < _15774;
    assign _16457 = ~ _16456;
    assign _16445 = _16354[53:53];
    assign _16442 = _16437 - _15774;
    assign _16443 = _16439 ? _16442 : _16437;
    assign _16444 = _16443[62:0];
    assign _16446 = { _16444,
                      _16445 };
    assign _16447 = _16446 < _15774;
    assign _16448 = ~ _16447;
    assign _16436 = _16354[54:54];
    assign _16433 = _16428 - _15774;
    assign _16434 = _16430 ? _16433 : _16428;
    assign _16435 = _16434[62:0];
    assign _16437 = { _16435,
                      _16436 };
    assign _16438 = _16437 < _15774;
    assign _16439 = ~ _16438;
    assign _16427 = _16354[55:55];
    assign _16424 = _16419 - _15774;
    assign _16425 = _16421 ? _16424 : _16419;
    assign _16426 = _16425[62:0];
    assign _16428 = { _16426,
                      _16427 };
    assign _16429 = _16428 < _15774;
    assign _16430 = ~ _16429;
    assign _16418 = _16354[56:56];
    assign _16415 = _16410 - _15774;
    assign _16416 = _16412 ? _16415 : _16410;
    assign _16417 = _16416[62:0];
    assign _16419 = { _16417,
                      _16418 };
    assign _16420 = _16419 < _15774;
    assign _16421 = ~ _16420;
    assign _16409 = _16354[57:57];
    assign _16406 = _16401 - _15774;
    assign _16407 = _16403 ? _16406 : _16401;
    assign _16408 = _16407[62:0];
    assign _16410 = { _16408,
                      _16409 };
    assign _16411 = _16410 < _15774;
    assign _16412 = ~ _16411;
    assign _16400 = _16354[58:58];
    assign _16397 = _16392 - _15774;
    assign _16398 = _16394 ? _16397 : _16392;
    assign _16399 = _16398[62:0];
    assign _16401 = { _16399,
                      _16400 };
    assign _16402 = _16401 < _15774;
    assign _16403 = ~ _16402;
    assign _16391 = _16354[59:59];
    assign _16388 = _16383 - _15774;
    assign _16389 = _16385 ? _16388 : _16383;
    assign _16390 = _16389[62:0];
    assign _16392 = { _16390,
                      _16391 };
    assign _16393 = _16392 < _15774;
    assign _16394 = ~ _16393;
    assign _16382 = _16354[60:60];
    assign _16379 = _16374 - _15774;
    assign _16380 = _16376 ? _16379 : _16374;
    assign _16381 = _16380[62:0];
    assign _16383 = { _16381,
                      _16382 };
    assign _16384 = _16383 < _15774;
    assign _16385 = ~ _16384;
    assign _16373 = _16354[61:61];
    assign _16370 = _16365 - _15774;
    assign _16371 = _16367 ? _16370 : _16365;
    assign _16372 = _16371[62:0];
    assign _16374 = { _16372,
                      _16373 };
    assign _16375 = _16374 < _15774;
    assign _16376 = ~ _16375;
    assign _16364 = _16354[62:62];
    assign _16361 = _16356 - _15774;
    assign _16362 = _16358 ? _16361 : _16356;
    assign _16363 = _16362[62:0];
    assign _16365 = { _16363,
                      _16364 };
    assign _16366 = _16365 < _15774;
    assign _16367 = ~ _16366;
    assign _16354 = _15766 - _16348;
    assign _16355 = _16354[63:63];
    assign _16356 = { _22185,
                      _16355 };
    assign _16357 = _16356 < _15774;
    assign _16358 = ~ _16357;
    assign _16359 = { _22185,
                      _16358 };
    assign _16360 = _16359[62:0];
    assign _16368 = { _16360,
                      _16367 };
    assign _16369 = _16368[62:0];
    assign _16377 = { _16369,
                      _16376 };
    assign _16378 = _16377[62:0];
    assign _16386 = { _16378,
                      _16385 };
    assign _16387 = _16386[62:0];
    assign _16395 = { _16387,
                      _16394 };
    assign _16396 = _16395[62:0];
    assign _16404 = { _16396,
                      _16403 };
    assign _16405 = _16404[62:0];
    assign _16413 = { _16405,
                      _16412 };
    assign _16414 = _16413[62:0];
    assign _16422 = { _16414,
                      _16421 };
    assign _16423 = _16422[62:0];
    assign _16431 = { _16423,
                      _16430 };
    assign _16432 = _16431[62:0];
    assign _16440 = { _16432,
                      _16439 };
    assign _16441 = _16440[62:0];
    assign _16449 = { _16441,
                      _16448 };
    assign _16450 = _16449[62:0];
    assign _16458 = { _16450,
                      _16457 };
    assign _16459 = _16458[62:0];
    assign _16467 = { _16459,
                      _16466 };
    assign _16468 = _16467[62:0];
    assign _16476 = { _16468,
                      _16475 };
    assign _16477 = _16476[62:0];
    assign _16485 = { _16477,
                      _16484 };
    assign _16486 = _16485[62:0];
    assign _16494 = { _16486,
                      _16493 };
    assign _16495 = _16494[62:0];
    assign _16503 = { _16495,
                      _16502 };
    assign _16504 = _16503[62:0];
    assign _16512 = { _16504,
                      _16511 };
    assign _16513 = _16512[62:0];
    assign _16521 = { _16513,
                      _16520 };
    assign _16522 = _16521[62:0];
    assign _16530 = { _16522,
                      _16529 };
    assign _16531 = _16530[62:0];
    assign _16539 = { _16531,
                      _16538 };
    assign _16540 = _16539[62:0];
    assign _16548 = { _16540,
                      _16547 };
    assign _16549 = _16548[62:0];
    assign _16557 = { _16549,
                      _16556 };
    assign _16558 = _16557[62:0];
    assign _16566 = { _16558,
                      _16565 };
    assign _16567 = _16566[62:0];
    assign _16575 = { _16567,
                      _16574 };
    assign _16576 = _16575[62:0];
    assign _16584 = { _16576,
                      _16583 };
    assign _16585 = _16584[62:0];
    assign _16593 = { _16585,
                      _16592 };
    assign _16594 = _16593[62:0];
    assign _16602 = { _16594,
                      _16601 };
    assign _16603 = _16602[62:0];
    assign _16611 = { _16603,
                      _16610 };
    assign _16612 = _16611[62:0];
    assign _16620 = { _16612,
                      _16619 };
    assign _16621 = _16620[62:0];
    assign _16629 = { _16621,
                      _16628 };
    assign _16630 = _16629[62:0];
    assign _16638 = { _16630,
                      _16637 };
    assign _16639 = _16638[62:0];
    assign _16647 = { _16639,
                      _16646 };
    assign _16648 = _16647[62:0];
    assign _16656 = { _16648,
                      _16655 };
    assign _16657 = _16656[62:0];
    assign _16665 = { _16657,
                      _16664 };
    assign _16666 = _16665[62:0];
    assign _16674 = { _16666,
                      _16673 };
    assign _16675 = _16674[62:0];
    assign _16683 = { _16675,
                      _16682 };
    assign _16684 = _16683[62:0];
    assign _16692 = { _16684,
                      _16691 };
    assign _16693 = _16692[62:0];
    assign _16701 = { _16693,
                      _16700 };
    assign _16702 = _16701[62:0];
    assign _16710 = { _16702,
                      _16709 };
    assign _16711 = _16710[62:0];
    assign _16719 = { _16711,
                      _16718 };
    assign _16720 = _16719[62:0];
    assign _16728 = { _16720,
                      _16727 };
    assign _16729 = _16728[62:0];
    assign _16737 = { _16729,
                      _16736 };
    assign _16738 = _16737[62:0];
    assign _16746 = { _16738,
                      _16745 };
    assign _16747 = _16746[62:0];
    assign _16755 = { _16747,
                      _16754 };
    assign _16756 = _16755[62:0];
    assign _16764 = { _16756,
                      _16763 };
    assign _16765 = _16764[62:0];
    assign _16773 = { _16765,
                      _16772 };
    assign _16774 = _16773[62:0];
    assign _16782 = { _16774,
                      _16781 };
    assign _16783 = _16782[62:0];
    assign _16791 = { _16783,
                      _16790 };
    assign _16792 = _16791[62:0];
    assign _16800 = { _16792,
                      _16799 };
    assign _16801 = _16800[62:0];
    assign _16809 = { _16801,
                      _16808 };
    assign _16810 = _16809[62:0];
    assign _16818 = { _16810,
                      _16817 };
    assign _16819 = _16818[62:0];
    assign _16827 = { _16819,
                      _16826 };
    assign _16828 = _16827[62:0];
    assign _16836 = { _16828,
                      _16835 };
    assign _16837 = _16836[62:0];
    assign _16845 = { _16837,
                      _16844 };
    assign _16846 = _16845[62:0];
    assign _16854 = { _16846,
                      _16853 };
    assign _16855 = _16854[62:0];
    assign _16863 = { _16855,
                      _16862 };
    assign _16864 = _16863[62:0];
    assign _16872 = { _16864,
                      _16871 };
    assign _16873 = _16872[62:0];
    assign _16881 = { _16873,
                      _16880 };
    assign _16882 = _16881[62:0];
    assign _16890 = { _16882,
                      _16889 };
    assign _16891 = _16890[62:0];
    assign _16899 = { _16891,
                      _16898 };
    assign _16900 = _16899[62:0];
    assign _16908 = { _16900,
                      _16907 };
    assign _16909 = _16908[62:0];
    assign _16917 = { _16909,
                      _16916 };
    assign _16918 = _16917[62:0];
    assign _16926 = { _16918,
                      _16925 };
    assign _16928 = _16926 + _22186;
    assign _16929 = _16928 * _16348;
    assign _16930 = _16929[63:0];
    assign _17512 = _16930 + _17511;
    assign _16340 = _15771[0:0];
    assign _16337 = _16332 - _15774;
    assign _16338 = _16334 ? _16337 : _16332;
    assign _16339 = _16338[62:0];
    assign _16341 = { _16339,
                      _16340 };
    assign _16342 = _16341 < _15774;
    assign _16343 = ~ _16342;
    assign _16331 = _15771[1:1];
    assign _16328 = _16323 - _15774;
    assign _16329 = _16325 ? _16328 : _16323;
    assign _16330 = _16329[62:0];
    assign _16332 = { _16330,
                      _16331 };
    assign _16333 = _16332 < _15774;
    assign _16334 = ~ _16333;
    assign _16322 = _15771[2:2];
    assign _16319 = _16314 - _15774;
    assign _16320 = _16316 ? _16319 : _16314;
    assign _16321 = _16320[62:0];
    assign _16323 = { _16321,
                      _16322 };
    assign _16324 = _16323 < _15774;
    assign _16325 = ~ _16324;
    assign _16313 = _15771[3:3];
    assign _16310 = _16305 - _15774;
    assign _16311 = _16307 ? _16310 : _16305;
    assign _16312 = _16311[62:0];
    assign _16314 = { _16312,
                      _16313 };
    assign _16315 = _16314 < _15774;
    assign _16316 = ~ _16315;
    assign _16304 = _15771[4:4];
    assign _16301 = _16296 - _15774;
    assign _16302 = _16298 ? _16301 : _16296;
    assign _16303 = _16302[62:0];
    assign _16305 = { _16303,
                      _16304 };
    assign _16306 = _16305 < _15774;
    assign _16307 = ~ _16306;
    assign _16295 = _15771[5:5];
    assign _16292 = _16287 - _15774;
    assign _16293 = _16289 ? _16292 : _16287;
    assign _16294 = _16293[62:0];
    assign _16296 = { _16294,
                      _16295 };
    assign _16297 = _16296 < _15774;
    assign _16298 = ~ _16297;
    assign _16286 = _15771[6:6];
    assign _16283 = _16278 - _15774;
    assign _16284 = _16280 ? _16283 : _16278;
    assign _16285 = _16284[62:0];
    assign _16287 = { _16285,
                      _16286 };
    assign _16288 = _16287 < _15774;
    assign _16289 = ~ _16288;
    assign _16277 = _15771[7:7];
    assign _16274 = _16269 - _15774;
    assign _16275 = _16271 ? _16274 : _16269;
    assign _16276 = _16275[62:0];
    assign _16278 = { _16276,
                      _16277 };
    assign _16279 = _16278 < _15774;
    assign _16280 = ~ _16279;
    assign _16268 = _15771[8:8];
    assign _16265 = _16260 - _15774;
    assign _16266 = _16262 ? _16265 : _16260;
    assign _16267 = _16266[62:0];
    assign _16269 = { _16267,
                      _16268 };
    assign _16270 = _16269 < _15774;
    assign _16271 = ~ _16270;
    assign _16259 = _15771[9:9];
    assign _16256 = _16251 - _15774;
    assign _16257 = _16253 ? _16256 : _16251;
    assign _16258 = _16257[62:0];
    assign _16260 = { _16258,
                      _16259 };
    assign _16261 = _16260 < _15774;
    assign _16262 = ~ _16261;
    assign _16250 = _15771[10:10];
    assign _16247 = _16242 - _15774;
    assign _16248 = _16244 ? _16247 : _16242;
    assign _16249 = _16248[62:0];
    assign _16251 = { _16249,
                      _16250 };
    assign _16252 = _16251 < _15774;
    assign _16253 = ~ _16252;
    assign _16241 = _15771[11:11];
    assign _16238 = _16233 - _15774;
    assign _16239 = _16235 ? _16238 : _16233;
    assign _16240 = _16239[62:0];
    assign _16242 = { _16240,
                      _16241 };
    assign _16243 = _16242 < _15774;
    assign _16244 = ~ _16243;
    assign _16232 = _15771[12:12];
    assign _16229 = _16224 - _15774;
    assign _16230 = _16226 ? _16229 : _16224;
    assign _16231 = _16230[62:0];
    assign _16233 = { _16231,
                      _16232 };
    assign _16234 = _16233 < _15774;
    assign _16235 = ~ _16234;
    assign _16223 = _15771[13:13];
    assign _16220 = _16215 - _15774;
    assign _16221 = _16217 ? _16220 : _16215;
    assign _16222 = _16221[62:0];
    assign _16224 = { _16222,
                      _16223 };
    assign _16225 = _16224 < _15774;
    assign _16226 = ~ _16225;
    assign _16214 = _15771[14:14];
    assign _16211 = _16206 - _15774;
    assign _16212 = _16208 ? _16211 : _16206;
    assign _16213 = _16212[62:0];
    assign _16215 = { _16213,
                      _16214 };
    assign _16216 = _16215 < _15774;
    assign _16217 = ~ _16216;
    assign _16205 = _15771[15:15];
    assign _16202 = _16197 - _15774;
    assign _16203 = _16199 ? _16202 : _16197;
    assign _16204 = _16203[62:0];
    assign _16206 = { _16204,
                      _16205 };
    assign _16207 = _16206 < _15774;
    assign _16208 = ~ _16207;
    assign _16196 = _15771[16:16];
    assign _16193 = _16188 - _15774;
    assign _16194 = _16190 ? _16193 : _16188;
    assign _16195 = _16194[62:0];
    assign _16197 = { _16195,
                      _16196 };
    assign _16198 = _16197 < _15774;
    assign _16199 = ~ _16198;
    assign _16187 = _15771[17:17];
    assign _16184 = _16179 - _15774;
    assign _16185 = _16181 ? _16184 : _16179;
    assign _16186 = _16185[62:0];
    assign _16188 = { _16186,
                      _16187 };
    assign _16189 = _16188 < _15774;
    assign _16190 = ~ _16189;
    assign _16178 = _15771[18:18];
    assign _16175 = _16170 - _15774;
    assign _16176 = _16172 ? _16175 : _16170;
    assign _16177 = _16176[62:0];
    assign _16179 = { _16177,
                      _16178 };
    assign _16180 = _16179 < _15774;
    assign _16181 = ~ _16180;
    assign _16169 = _15771[19:19];
    assign _16166 = _16161 - _15774;
    assign _16167 = _16163 ? _16166 : _16161;
    assign _16168 = _16167[62:0];
    assign _16170 = { _16168,
                      _16169 };
    assign _16171 = _16170 < _15774;
    assign _16172 = ~ _16171;
    assign _16160 = _15771[20:20];
    assign _16157 = _16152 - _15774;
    assign _16158 = _16154 ? _16157 : _16152;
    assign _16159 = _16158[62:0];
    assign _16161 = { _16159,
                      _16160 };
    assign _16162 = _16161 < _15774;
    assign _16163 = ~ _16162;
    assign _16151 = _15771[21:21];
    assign _16148 = _16143 - _15774;
    assign _16149 = _16145 ? _16148 : _16143;
    assign _16150 = _16149[62:0];
    assign _16152 = { _16150,
                      _16151 };
    assign _16153 = _16152 < _15774;
    assign _16154 = ~ _16153;
    assign _16142 = _15771[22:22];
    assign _16139 = _16134 - _15774;
    assign _16140 = _16136 ? _16139 : _16134;
    assign _16141 = _16140[62:0];
    assign _16143 = { _16141,
                      _16142 };
    assign _16144 = _16143 < _15774;
    assign _16145 = ~ _16144;
    assign _16133 = _15771[23:23];
    assign _16130 = _16125 - _15774;
    assign _16131 = _16127 ? _16130 : _16125;
    assign _16132 = _16131[62:0];
    assign _16134 = { _16132,
                      _16133 };
    assign _16135 = _16134 < _15774;
    assign _16136 = ~ _16135;
    assign _16124 = _15771[24:24];
    assign _16121 = _16116 - _15774;
    assign _16122 = _16118 ? _16121 : _16116;
    assign _16123 = _16122[62:0];
    assign _16125 = { _16123,
                      _16124 };
    assign _16126 = _16125 < _15774;
    assign _16127 = ~ _16126;
    assign _16115 = _15771[25:25];
    assign _16112 = _16107 - _15774;
    assign _16113 = _16109 ? _16112 : _16107;
    assign _16114 = _16113[62:0];
    assign _16116 = { _16114,
                      _16115 };
    assign _16117 = _16116 < _15774;
    assign _16118 = ~ _16117;
    assign _16106 = _15771[26:26];
    assign _16103 = _16098 - _15774;
    assign _16104 = _16100 ? _16103 : _16098;
    assign _16105 = _16104[62:0];
    assign _16107 = { _16105,
                      _16106 };
    assign _16108 = _16107 < _15774;
    assign _16109 = ~ _16108;
    assign _16097 = _15771[27:27];
    assign _16094 = _16089 - _15774;
    assign _16095 = _16091 ? _16094 : _16089;
    assign _16096 = _16095[62:0];
    assign _16098 = { _16096,
                      _16097 };
    assign _16099 = _16098 < _15774;
    assign _16100 = ~ _16099;
    assign _16088 = _15771[28:28];
    assign _16085 = _16080 - _15774;
    assign _16086 = _16082 ? _16085 : _16080;
    assign _16087 = _16086[62:0];
    assign _16089 = { _16087,
                      _16088 };
    assign _16090 = _16089 < _15774;
    assign _16091 = ~ _16090;
    assign _16079 = _15771[29:29];
    assign _16076 = _16071 - _15774;
    assign _16077 = _16073 ? _16076 : _16071;
    assign _16078 = _16077[62:0];
    assign _16080 = { _16078,
                      _16079 };
    assign _16081 = _16080 < _15774;
    assign _16082 = ~ _16081;
    assign _16070 = _15771[30:30];
    assign _16067 = _16062 - _15774;
    assign _16068 = _16064 ? _16067 : _16062;
    assign _16069 = _16068[62:0];
    assign _16071 = { _16069,
                      _16070 };
    assign _16072 = _16071 < _15774;
    assign _16073 = ~ _16072;
    assign _16061 = _15771[31:31];
    assign _16058 = _16053 - _15774;
    assign _16059 = _16055 ? _16058 : _16053;
    assign _16060 = _16059[62:0];
    assign _16062 = { _16060,
                      _16061 };
    assign _16063 = _16062 < _15774;
    assign _16064 = ~ _16063;
    assign _16052 = _15771[32:32];
    assign _16049 = _16044 - _15774;
    assign _16050 = _16046 ? _16049 : _16044;
    assign _16051 = _16050[62:0];
    assign _16053 = { _16051,
                      _16052 };
    assign _16054 = _16053 < _15774;
    assign _16055 = ~ _16054;
    assign _16043 = _15771[33:33];
    assign _16040 = _16035 - _15774;
    assign _16041 = _16037 ? _16040 : _16035;
    assign _16042 = _16041[62:0];
    assign _16044 = { _16042,
                      _16043 };
    assign _16045 = _16044 < _15774;
    assign _16046 = ~ _16045;
    assign _16034 = _15771[34:34];
    assign _16031 = _16026 - _15774;
    assign _16032 = _16028 ? _16031 : _16026;
    assign _16033 = _16032[62:0];
    assign _16035 = { _16033,
                      _16034 };
    assign _16036 = _16035 < _15774;
    assign _16037 = ~ _16036;
    assign _16025 = _15771[35:35];
    assign _16022 = _16017 - _15774;
    assign _16023 = _16019 ? _16022 : _16017;
    assign _16024 = _16023[62:0];
    assign _16026 = { _16024,
                      _16025 };
    assign _16027 = _16026 < _15774;
    assign _16028 = ~ _16027;
    assign _16016 = _15771[36:36];
    assign _16013 = _16008 - _15774;
    assign _16014 = _16010 ? _16013 : _16008;
    assign _16015 = _16014[62:0];
    assign _16017 = { _16015,
                      _16016 };
    assign _16018 = _16017 < _15774;
    assign _16019 = ~ _16018;
    assign _16007 = _15771[37:37];
    assign _16004 = _15999 - _15774;
    assign _16005 = _16001 ? _16004 : _15999;
    assign _16006 = _16005[62:0];
    assign _16008 = { _16006,
                      _16007 };
    assign _16009 = _16008 < _15774;
    assign _16010 = ~ _16009;
    assign _15998 = _15771[38:38];
    assign _15995 = _15990 - _15774;
    assign _15996 = _15992 ? _15995 : _15990;
    assign _15997 = _15996[62:0];
    assign _15999 = { _15997,
                      _15998 };
    assign _16000 = _15999 < _15774;
    assign _16001 = ~ _16000;
    assign _15989 = _15771[39:39];
    assign _15986 = _15981 - _15774;
    assign _15987 = _15983 ? _15986 : _15981;
    assign _15988 = _15987[62:0];
    assign _15990 = { _15988,
                      _15989 };
    assign _15991 = _15990 < _15774;
    assign _15992 = ~ _15991;
    assign _15980 = _15771[40:40];
    assign _15977 = _15972 - _15774;
    assign _15978 = _15974 ? _15977 : _15972;
    assign _15979 = _15978[62:0];
    assign _15981 = { _15979,
                      _15980 };
    assign _15982 = _15981 < _15774;
    assign _15983 = ~ _15982;
    assign _15971 = _15771[41:41];
    assign _15968 = _15963 - _15774;
    assign _15969 = _15965 ? _15968 : _15963;
    assign _15970 = _15969[62:0];
    assign _15972 = { _15970,
                      _15971 };
    assign _15973 = _15972 < _15774;
    assign _15974 = ~ _15973;
    assign _15962 = _15771[42:42];
    assign _15959 = _15954 - _15774;
    assign _15960 = _15956 ? _15959 : _15954;
    assign _15961 = _15960[62:0];
    assign _15963 = { _15961,
                      _15962 };
    assign _15964 = _15963 < _15774;
    assign _15965 = ~ _15964;
    assign _15953 = _15771[43:43];
    assign _15950 = _15945 - _15774;
    assign _15951 = _15947 ? _15950 : _15945;
    assign _15952 = _15951[62:0];
    assign _15954 = { _15952,
                      _15953 };
    assign _15955 = _15954 < _15774;
    assign _15956 = ~ _15955;
    assign _15944 = _15771[44:44];
    assign _15941 = _15936 - _15774;
    assign _15942 = _15938 ? _15941 : _15936;
    assign _15943 = _15942[62:0];
    assign _15945 = { _15943,
                      _15944 };
    assign _15946 = _15945 < _15774;
    assign _15947 = ~ _15946;
    assign _15935 = _15771[45:45];
    assign _15932 = _15927 - _15774;
    assign _15933 = _15929 ? _15932 : _15927;
    assign _15934 = _15933[62:0];
    assign _15936 = { _15934,
                      _15935 };
    assign _15937 = _15936 < _15774;
    assign _15938 = ~ _15937;
    assign _15926 = _15771[46:46];
    assign _15923 = _15918 - _15774;
    assign _15924 = _15920 ? _15923 : _15918;
    assign _15925 = _15924[62:0];
    assign _15927 = { _15925,
                      _15926 };
    assign _15928 = _15927 < _15774;
    assign _15929 = ~ _15928;
    assign _15917 = _15771[47:47];
    assign _15914 = _15909 - _15774;
    assign _15915 = _15911 ? _15914 : _15909;
    assign _15916 = _15915[62:0];
    assign _15918 = { _15916,
                      _15917 };
    assign _15919 = _15918 < _15774;
    assign _15920 = ~ _15919;
    assign _15908 = _15771[48:48];
    assign _15905 = _15900 - _15774;
    assign _15906 = _15902 ? _15905 : _15900;
    assign _15907 = _15906[62:0];
    assign _15909 = { _15907,
                      _15908 };
    assign _15910 = _15909 < _15774;
    assign _15911 = ~ _15910;
    assign _15899 = _15771[49:49];
    assign _15896 = _15891 - _15774;
    assign _15897 = _15893 ? _15896 : _15891;
    assign _15898 = _15897[62:0];
    assign _15900 = { _15898,
                      _15899 };
    assign _15901 = _15900 < _15774;
    assign _15902 = ~ _15901;
    assign _15890 = _15771[50:50];
    assign _15887 = _15882 - _15774;
    assign _15888 = _15884 ? _15887 : _15882;
    assign _15889 = _15888[62:0];
    assign _15891 = { _15889,
                      _15890 };
    assign _15892 = _15891 < _15774;
    assign _15893 = ~ _15892;
    assign _15881 = _15771[51:51];
    assign _15878 = _15873 - _15774;
    assign _15879 = _15875 ? _15878 : _15873;
    assign _15880 = _15879[62:0];
    assign _15882 = { _15880,
                      _15881 };
    assign _15883 = _15882 < _15774;
    assign _15884 = ~ _15883;
    assign _15872 = _15771[52:52];
    assign _15869 = _15864 - _15774;
    assign _15870 = _15866 ? _15869 : _15864;
    assign _15871 = _15870[62:0];
    assign _15873 = { _15871,
                      _15872 };
    assign _15874 = _15873 < _15774;
    assign _15875 = ~ _15874;
    assign _15863 = _15771[53:53];
    assign _15860 = _15855 - _15774;
    assign _15861 = _15857 ? _15860 : _15855;
    assign _15862 = _15861[62:0];
    assign _15864 = { _15862,
                      _15863 };
    assign _15865 = _15864 < _15774;
    assign _15866 = ~ _15865;
    assign _15854 = _15771[54:54];
    assign _15851 = _15846 - _15774;
    assign _15852 = _15848 ? _15851 : _15846;
    assign _15853 = _15852[62:0];
    assign _15855 = { _15853,
                      _15854 };
    assign _15856 = _15855 < _15774;
    assign _15857 = ~ _15856;
    assign _15845 = _15771[55:55];
    assign _15842 = _15837 - _15774;
    assign _15843 = _15839 ? _15842 : _15837;
    assign _15844 = _15843[62:0];
    assign _15846 = { _15844,
                      _15845 };
    assign _15847 = _15846 < _15774;
    assign _15848 = ~ _15847;
    assign _15836 = _15771[56:56];
    assign _15833 = _15828 - _15774;
    assign _15834 = _15830 ? _15833 : _15828;
    assign _15835 = _15834[62:0];
    assign _15837 = { _15835,
                      _15836 };
    assign _15838 = _15837 < _15774;
    assign _15839 = ~ _15838;
    assign _15827 = _15771[57:57];
    assign _15824 = _15819 - _15774;
    assign _15825 = _15821 ? _15824 : _15819;
    assign _15826 = _15825[62:0];
    assign _15828 = { _15826,
                      _15827 };
    assign _15829 = _15828 < _15774;
    assign _15830 = ~ _15829;
    assign _15818 = _15771[58:58];
    assign _15815 = _15810 - _15774;
    assign _15816 = _15812 ? _15815 : _15810;
    assign _15817 = _15816[62:0];
    assign _15819 = { _15817,
                      _15818 };
    assign _15820 = _15819 < _15774;
    assign _15821 = ~ _15820;
    assign _15809 = _15771[59:59];
    assign _15806 = _15801 - _15774;
    assign _15807 = _15803 ? _15806 : _15801;
    assign _15808 = _15807[62:0];
    assign _15810 = { _15808,
                      _15809 };
    assign _15811 = _15810 < _15774;
    assign _15812 = ~ _15811;
    assign _15800 = _15771[60:60];
    assign _15797 = _15792 - _15774;
    assign _15798 = _15794 ? _15797 : _15792;
    assign _15799 = _15798[62:0];
    assign _15801 = { _15799,
                      _15800 };
    assign _15802 = _15801 < _15774;
    assign _15803 = ~ _15802;
    assign _15791 = _15771[61:61];
    assign _15788 = _15783 - _15774;
    assign _15789 = _15785 ? _15788 : _15783;
    assign _15790 = _15789[62:0];
    assign _15792 = { _15790,
                      _15791 };
    assign _15793 = _15792 < _15774;
    assign _15794 = ~ _15793;
    assign _15782 = _15771[62:62];
    assign _15779 = _15773 - _15774;
    assign _15780 = _15776 ? _15779 : _15773;
    assign _15781 = _15780[62:0];
    assign _15783 = { _15781,
                      _15782 };
    assign _15784 = _15783 < _15774;
    assign _15785 = ~ _15784;
    assign _15774 = 64'b0000000000000000000000000000000000000000000011110100011000101001;
    assign _15770 = 64'b0000000000000000000000000000000000000000000011110100011000101000;
    assign _15771 = _3 + _15770;
    assign _15772 = _15771[63:63];
    assign _15773 = { _22185,
                      _15772 };
    assign _15775 = _15773 < _15774;
    assign _15776 = ~ _15775;
    assign _15777 = { _22185,
                      _15776 };
    assign _15778 = _15777[62:0];
    assign _15786 = { _15778,
                      _15785 };
    assign _15787 = _15786[62:0];
    assign _15795 = { _15787,
                      _15794 };
    assign _15796 = _15795[62:0];
    assign _15804 = { _15796,
                      _15803 };
    assign _15805 = _15804[62:0];
    assign _15813 = { _15805,
                      _15812 };
    assign _15814 = _15813[62:0];
    assign _15822 = { _15814,
                      _15821 };
    assign _15823 = _15822[62:0];
    assign _15831 = { _15823,
                      _15830 };
    assign _15832 = _15831[62:0];
    assign _15840 = { _15832,
                      _15839 };
    assign _15841 = _15840[62:0];
    assign _15849 = { _15841,
                      _15848 };
    assign _15850 = _15849[62:0];
    assign _15858 = { _15850,
                      _15857 };
    assign _15859 = _15858[62:0];
    assign _15867 = { _15859,
                      _15866 };
    assign _15868 = _15867[62:0];
    assign _15876 = { _15868,
                      _15875 };
    assign _15877 = _15876[62:0];
    assign _15885 = { _15877,
                      _15884 };
    assign _15886 = _15885[62:0];
    assign _15894 = { _15886,
                      _15893 };
    assign _15895 = _15894[62:0];
    assign _15903 = { _15895,
                      _15902 };
    assign _15904 = _15903[62:0];
    assign _15912 = { _15904,
                      _15911 };
    assign _15913 = _15912[62:0];
    assign _15921 = { _15913,
                      _15920 };
    assign _15922 = _15921[62:0];
    assign _15930 = { _15922,
                      _15929 };
    assign _15931 = _15930[62:0];
    assign _15939 = { _15931,
                      _15938 };
    assign _15940 = _15939[62:0];
    assign _15948 = { _15940,
                      _15947 };
    assign _15949 = _15948[62:0];
    assign _15957 = { _15949,
                      _15956 };
    assign _15958 = _15957[62:0];
    assign _15966 = { _15958,
                      _15965 };
    assign _15967 = _15966[62:0];
    assign _15975 = { _15967,
                      _15974 };
    assign _15976 = _15975[62:0];
    assign _15984 = { _15976,
                      _15983 };
    assign _15985 = _15984[62:0];
    assign _15993 = { _15985,
                      _15992 };
    assign _15994 = _15993[62:0];
    assign _16002 = { _15994,
                      _16001 };
    assign _16003 = _16002[62:0];
    assign _16011 = { _16003,
                      _16010 };
    assign _16012 = _16011[62:0];
    assign _16020 = { _16012,
                      _16019 };
    assign _16021 = _16020[62:0];
    assign _16029 = { _16021,
                      _16028 };
    assign _16030 = _16029[62:0];
    assign _16038 = { _16030,
                      _16037 };
    assign _16039 = _16038[62:0];
    assign _16047 = { _16039,
                      _16046 };
    assign _16048 = _16047[62:0];
    assign _16056 = { _16048,
                      _16055 };
    assign _16057 = _16056[62:0];
    assign _16065 = { _16057,
                      _16064 };
    assign _16066 = _16065[62:0];
    assign _16074 = { _16066,
                      _16073 };
    assign _16075 = _16074[62:0];
    assign _16083 = { _16075,
                      _16082 };
    assign _16084 = _16083[62:0];
    assign _16092 = { _16084,
                      _16091 };
    assign _16093 = _16092[62:0];
    assign _16101 = { _16093,
                      _16100 };
    assign _16102 = _16101[62:0];
    assign _16110 = { _16102,
                      _16109 };
    assign _16111 = _16110[62:0];
    assign _16119 = { _16111,
                      _16118 };
    assign _16120 = _16119[62:0];
    assign _16128 = { _16120,
                      _16127 };
    assign _16129 = _16128[62:0];
    assign _16137 = { _16129,
                      _16136 };
    assign _16138 = _16137[62:0];
    assign _16146 = { _16138,
                      _16145 };
    assign _16147 = _16146[62:0];
    assign _16155 = { _16147,
                      _16154 };
    assign _16156 = _16155[62:0];
    assign _16164 = { _16156,
                      _16163 };
    assign _16165 = _16164[62:0];
    assign _16173 = { _16165,
                      _16172 };
    assign _16174 = _16173[62:0];
    assign _16182 = { _16174,
                      _16181 };
    assign _16183 = _16182[62:0];
    assign _16191 = { _16183,
                      _16190 };
    assign _16192 = _16191[62:0];
    assign _16200 = { _16192,
                      _16199 };
    assign _16201 = _16200[62:0];
    assign _16209 = { _16201,
                      _16208 };
    assign _16210 = _16209[62:0];
    assign _16218 = { _16210,
                      _16217 };
    assign _16219 = _16218[62:0];
    assign _16227 = { _16219,
                      _16226 };
    assign _16228 = _16227[62:0];
    assign _16236 = { _16228,
                      _16235 };
    assign _16237 = _16236[62:0];
    assign _16245 = { _16237,
                      _16244 };
    assign _16246 = _16245[62:0];
    assign _16254 = { _16246,
                      _16253 };
    assign _16255 = _16254[62:0];
    assign _16263 = { _16255,
                      _16262 };
    assign _16264 = _16263[62:0];
    assign _16272 = { _16264,
                      _16271 };
    assign _16273 = _16272[62:0];
    assign _16281 = { _16273,
                      _16280 };
    assign _16282 = _16281[62:0];
    assign _16290 = { _16282,
                      _16289 };
    assign _16291 = _16290[62:0];
    assign _16299 = { _16291,
                      _16298 };
    assign _16300 = _16299[62:0];
    assign _16308 = { _16300,
                      _16307 };
    assign _16309 = _16308[62:0];
    assign _16317 = { _16309,
                      _16316 };
    assign _16318 = _16317[62:0];
    assign _16326 = { _16318,
                      _16325 };
    assign _16327 = _16326[62:0];
    assign _16335 = { _16327,
                      _16334 };
    assign _16336 = _16335[62:0];
    assign _16344 = { _16336,
                      _16343 };
    assign _16345 = _16344 * _15774;
    assign _16346 = _16345[63:0];
    assign _15767 = 64'b0000000000000000000000000000000000000101111101110110100000000100;
    assign _16347 = _15767 < _16346;
    assign _16348 = _16347 ? _16346 : _15767;
    assign _15764 = 64'b0000000000000000000000000000000000111011100110101100100111111111;
    assign _15765 = _5 < _15764;
    assign _15766 = _15765 ? _5 : _15764;
    assign _16349 = _15766 < _16348;
    assign _16350 = ~ _16349;
    assign _17513 = _16350 ? _17512 : _21604;
    assign _15754 = _15185[0:0];
    assign _15751 = _15746 - _22192;
    assign _15752 = _15748 ? _15751 : _15746;
    assign _15753 = _15752[62:0];
    assign _15755 = { _15753,
                      _15754 };
    assign _15756 = _15755 < _22192;
    assign _15757 = ~ _15756;
    assign _15745 = _15185[1:1];
    assign _15742 = _15737 - _22192;
    assign _15743 = _15739 ? _15742 : _15737;
    assign _15744 = _15743[62:0];
    assign _15746 = { _15744,
                      _15745 };
    assign _15747 = _15746 < _22192;
    assign _15748 = ~ _15747;
    assign _15736 = _15185[2:2];
    assign _15733 = _15728 - _22192;
    assign _15734 = _15730 ? _15733 : _15728;
    assign _15735 = _15734[62:0];
    assign _15737 = { _15735,
                      _15736 };
    assign _15738 = _15737 < _22192;
    assign _15739 = ~ _15738;
    assign _15727 = _15185[3:3];
    assign _15724 = _15719 - _22192;
    assign _15725 = _15721 ? _15724 : _15719;
    assign _15726 = _15725[62:0];
    assign _15728 = { _15726,
                      _15727 };
    assign _15729 = _15728 < _22192;
    assign _15730 = ~ _15729;
    assign _15718 = _15185[4:4];
    assign _15715 = _15710 - _22192;
    assign _15716 = _15712 ? _15715 : _15710;
    assign _15717 = _15716[62:0];
    assign _15719 = { _15717,
                      _15718 };
    assign _15720 = _15719 < _22192;
    assign _15721 = ~ _15720;
    assign _15709 = _15185[5:5];
    assign _15706 = _15701 - _22192;
    assign _15707 = _15703 ? _15706 : _15701;
    assign _15708 = _15707[62:0];
    assign _15710 = { _15708,
                      _15709 };
    assign _15711 = _15710 < _22192;
    assign _15712 = ~ _15711;
    assign _15700 = _15185[6:6];
    assign _15697 = _15692 - _22192;
    assign _15698 = _15694 ? _15697 : _15692;
    assign _15699 = _15698[62:0];
    assign _15701 = { _15699,
                      _15700 };
    assign _15702 = _15701 < _22192;
    assign _15703 = ~ _15702;
    assign _15691 = _15185[7:7];
    assign _15688 = _15683 - _22192;
    assign _15689 = _15685 ? _15688 : _15683;
    assign _15690 = _15689[62:0];
    assign _15692 = { _15690,
                      _15691 };
    assign _15693 = _15692 < _22192;
    assign _15694 = ~ _15693;
    assign _15682 = _15185[8:8];
    assign _15679 = _15674 - _22192;
    assign _15680 = _15676 ? _15679 : _15674;
    assign _15681 = _15680[62:0];
    assign _15683 = { _15681,
                      _15682 };
    assign _15684 = _15683 < _22192;
    assign _15685 = ~ _15684;
    assign _15673 = _15185[9:9];
    assign _15670 = _15665 - _22192;
    assign _15671 = _15667 ? _15670 : _15665;
    assign _15672 = _15671[62:0];
    assign _15674 = { _15672,
                      _15673 };
    assign _15675 = _15674 < _22192;
    assign _15676 = ~ _15675;
    assign _15664 = _15185[10:10];
    assign _15661 = _15656 - _22192;
    assign _15662 = _15658 ? _15661 : _15656;
    assign _15663 = _15662[62:0];
    assign _15665 = { _15663,
                      _15664 };
    assign _15666 = _15665 < _22192;
    assign _15667 = ~ _15666;
    assign _15655 = _15185[11:11];
    assign _15652 = _15647 - _22192;
    assign _15653 = _15649 ? _15652 : _15647;
    assign _15654 = _15653[62:0];
    assign _15656 = { _15654,
                      _15655 };
    assign _15657 = _15656 < _22192;
    assign _15658 = ~ _15657;
    assign _15646 = _15185[12:12];
    assign _15643 = _15638 - _22192;
    assign _15644 = _15640 ? _15643 : _15638;
    assign _15645 = _15644[62:0];
    assign _15647 = { _15645,
                      _15646 };
    assign _15648 = _15647 < _22192;
    assign _15649 = ~ _15648;
    assign _15637 = _15185[13:13];
    assign _15634 = _15629 - _22192;
    assign _15635 = _15631 ? _15634 : _15629;
    assign _15636 = _15635[62:0];
    assign _15638 = { _15636,
                      _15637 };
    assign _15639 = _15638 < _22192;
    assign _15640 = ~ _15639;
    assign _15628 = _15185[14:14];
    assign _15625 = _15620 - _22192;
    assign _15626 = _15622 ? _15625 : _15620;
    assign _15627 = _15626[62:0];
    assign _15629 = { _15627,
                      _15628 };
    assign _15630 = _15629 < _22192;
    assign _15631 = ~ _15630;
    assign _15619 = _15185[15:15];
    assign _15616 = _15611 - _22192;
    assign _15617 = _15613 ? _15616 : _15611;
    assign _15618 = _15617[62:0];
    assign _15620 = { _15618,
                      _15619 };
    assign _15621 = _15620 < _22192;
    assign _15622 = ~ _15621;
    assign _15610 = _15185[16:16];
    assign _15607 = _15602 - _22192;
    assign _15608 = _15604 ? _15607 : _15602;
    assign _15609 = _15608[62:0];
    assign _15611 = { _15609,
                      _15610 };
    assign _15612 = _15611 < _22192;
    assign _15613 = ~ _15612;
    assign _15601 = _15185[17:17];
    assign _15598 = _15593 - _22192;
    assign _15599 = _15595 ? _15598 : _15593;
    assign _15600 = _15599[62:0];
    assign _15602 = { _15600,
                      _15601 };
    assign _15603 = _15602 < _22192;
    assign _15604 = ~ _15603;
    assign _15592 = _15185[18:18];
    assign _15589 = _15584 - _22192;
    assign _15590 = _15586 ? _15589 : _15584;
    assign _15591 = _15590[62:0];
    assign _15593 = { _15591,
                      _15592 };
    assign _15594 = _15593 < _22192;
    assign _15595 = ~ _15594;
    assign _15583 = _15185[19:19];
    assign _15580 = _15575 - _22192;
    assign _15581 = _15577 ? _15580 : _15575;
    assign _15582 = _15581[62:0];
    assign _15584 = { _15582,
                      _15583 };
    assign _15585 = _15584 < _22192;
    assign _15586 = ~ _15585;
    assign _15574 = _15185[20:20];
    assign _15571 = _15566 - _22192;
    assign _15572 = _15568 ? _15571 : _15566;
    assign _15573 = _15572[62:0];
    assign _15575 = { _15573,
                      _15574 };
    assign _15576 = _15575 < _22192;
    assign _15577 = ~ _15576;
    assign _15565 = _15185[21:21];
    assign _15562 = _15557 - _22192;
    assign _15563 = _15559 ? _15562 : _15557;
    assign _15564 = _15563[62:0];
    assign _15566 = { _15564,
                      _15565 };
    assign _15567 = _15566 < _22192;
    assign _15568 = ~ _15567;
    assign _15556 = _15185[22:22];
    assign _15553 = _15548 - _22192;
    assign _15554 = _15550 ? _15553 : _15548;
    assign _15555 = _15554[62:0];
    assign _15557 = { _15555,
                      _15556 };
    assign _15558 = _15557 < _22192;
    assign _15559 = ~ _15558;
    assign _15547 = _15185[23:23];
    assign _15544 = _15539 - _22192;
    assign _15545 = _15541 ? _15544 : _15539;
    assign _15546 = _15545[62:0];
    assign _15548 = { _15546,
                      _15547 };
    assign _15549 = _15548 < _22192;
    assign _15550 = ~ _15549;
    assign _15538 = _15185[24:24];
    assign _15535 = _15530 - _22192;
    assign _15536 = _15532 ? _15535 : _15530;
    assign _15537 = _15536[62:0];
    assign _15539 = { _15537,
                      _15538 };
    assign _15540 = _15539 < _22192;
    assign _15541 = ~ _15540;
    assign _15529 = _15185[25:25];
    assign _15526 = _15521 - _22192;
    assign _15527 = _15523 ? _15526 : _15521;
    assign _15528 = _15527[62:0];
    assign _15530 = { _15528,
                      _15529 };
    assign _15531 = _15530 < _22192;
    assign _15532 = ~ _15531;
    assign _15520 = _15185[26:26];
    assign _15517 = _15512 - _22192;
    assign _15518 = _15514 ? _15517 : _15512;
    assign _15519 = _15518[62:0];
    assign _15521 = { _15519,
                      _15520 };
    assign _15522 = _15521 < _22192;
    assign _15523 = ~ _15522;
    assign _15511 = _15185[27:27];
    assign _15508 = _15503 - _22192;
    assign _15509 = _15505 ? _15508 : _15503;
    assign _15510 = _15509[62:0];
    assign _15512 = { _15510,
                      _15511 };
    assign _15513 = _15512 < _22192;
    assign _15514 = ~ _15513;
    assign _15502 = _15185[28:28];
    assign _15499 = _15494 - _22192;
    assign _15500 = _15496 ? _15499 : _15494;
    assign _15501 = _15500[62:0];
    assign _15503 = { _15501,
                      _15502 };
    assign _15504 = _15503 < _22192;
    assign _15505 = ~ _15504;
    assign _15493 = _15185[29:29];
    assign _15490 = _15485 - _22192;
    assign _15491 = _15487 ? _15490 : _15485;
    assign _15492 = _15491[62:0];
    assign _15494 = { _15492,
                      _15493 };
    assign _15495 = _15494 < _22192;
    assign _15496 = ~ _15495;
    assign _15484 = _15185[30:30];
    assign _15481 = _15476 - _22192;
    assign _15482 = _15478 ? _15481 : _15476;
    assign _15483 = _15482[62:0];
    assign _15485 = { _15483,
                      _15484 };
    assign _15486 = _15485 < _22192;
    assign _15487 = ~ _15486;
    assign _15475 = _15185[31:31];
    assign _15472 = _15467 - _22192;
    assign _15473 = _15469 ? _15472 : _15467;
    assign _15474 = _15473[62:0];
    assign _15476 = { _15474,
                      _15475 };
    assign _15477 = _15476 < _22192;
    assign _15478 = ~ _15477;
    assign _15466 = _15185[32:32];
    assign _15463 = _15458 - _22192;
    assign _15464 = _15460 ? _15463 : _15458;
    assign _15465 = _15464[62:0];
    assign _15467 = { _15465,
                      _15466 };
    assign _15468 = _15467 < _22192;
    assign _15469 = ~ _15468;
    assign _15457 = _15185[33:33];
    assign _15454 = _15449 - _22192;
    assign _15455 = _15451 ? _15454 : _15449;
    assign _15456 = _15455[62:0];
    assign _15458 = { _15456,
                      _15457 };
    assign _15459 = _15458 < _22192;
    assign _15460 = ~ _15459;
    assign _15448 = _15185[34:34];
    assign _15445 = _15440 - _22192;
    assign _15446 = _15442 ? _15445 : _15440;
    assign _15447 = _15446[62:0];
    assign _15449 = { _15447,
                      _15448 };
    assign _15450 = _15449 < _22192;
    assign _15451 = ~ _15450;
    assign _15439 = _15185[35:35];
    assign _15436 = _15431 - _22192;
    assign _15437 = _15433 ? _15436 : _15431;
    assign _15438 = _15437[62:0];
    assign _15440 = { _15438,
                      _15439 };
    assign _15441 = _15440 < _22192;
    assign _15442 = ~ _15441;
    assign _15430 = _15185[36:36];
    assign _15427 = _15422 - _22192;
    assign _15428 = _15424 ? _15427 : _15422;
    assign _15429 = _15428[62:0];
    assign _15431 = { _15429,
                      _15430 };
    assign _15432 = _15431 < _22192;
    assign _15433 = ~ _15432;
    assign _15421 = _15185[37:37];
    assign _15418 = _15413 - _22192;
    assign _15419 = _15415 ? _15418 : _15413;
    assign _15420 = _15419[62:0];
    assign _15422 = { _15420,
                      _15421 };
    assign _15423 = _15422 < _22192;
    assign _15424 = ~ _15423;
    assign _15412 = _15185[38:38];
    assign _15409 = _15404 - _22192;
    assign _15410 = _15406 ? _15409 : _15404;
    assign _15411 = _15410[62:0];
    assign _15413 = { _15411,
                      _15412 };
    assign _15414 = _15413 < _22192;
    assign _15415 = ~ _15414;
    assign _15403 = _15185[39:39];
    assign _15400 = _15395 - _22192;
    assign _15401 = _15397 ? _15400 : _15395;
    assign _15402 = _15401[62:0];
    assign _15404 = { _15402,
                      _15403 };
    assign _15405 = _15404 < _22192;
    assign _15406 = ~ _15405;
    assign _15394 = _15185[40:40];
    assign _15391 = _15386 - _22192;
    assign _15392 = _15388 ? _15391 : _15386;
    assign _15393 = _15392[62:0];
    assign _15395 = { _15393,
                      _15394 };
    assign _15396 = _15395 < _22192;
    assign _15397 = ~ _15396;
    assign _15385 = _15185[41:41];
    assign _15382 = _15377 - _22192;
    assign _15383 = _15379 ? _15382 : _15377;
    assign _15384 = _15383[62:0];
    assign _15386 = { _15384,
                      _15385 };
    assign _15387 = _15386 < _22192;
    assign _15388 = ~ _15387;
    assign _15376 = _15185[42:42];
    assign _15373 = _15368 - _22192;
    assign _15374 = _15370 ? _15373 : _15368;
    assign _15375 = _15374[62:0];
    assign _15377 = { _15375,
                      _15376 };
    assign _15378 = _15377 < _22192;
    assign _15379 = ~ _15378;
    assign _15367 = _15185[43:43];
    assign _15364 = _15359 - _22192;
    assign _15365 = _15361 ? _15364 : _15359;
    assign _15366 = _15365[62:0];
    assign _15368 = { _15366,
                      _15367 };
    assign _15369 = _15368 < _22192;
    assign _15370 = ~ _15369;
    assign _15358 = _15185[44:44];
    assign _15355 = _15350 - _22192;
    assign _15356 = _15352 ? _15355 : _15350;
    assign _15357 = _15356[62:0];
    assign _15359 = { _15357,
                      _15358 };
    assign _15360 = _15359 < _22192;
    assign _15361 = ~ _15360;
    assign _15349 = _15185[45:45];
    assign _15346 = _15341 - _22192;
    assign _15347 = _15343 ? _15346 : _15341;
    assign _15348 = _15347[62:0];
    assign _15350 = { _15348,
                      _15349 };
    assign _15351 = _15350 < _22192;
    assign _15352 = ~ _15351;
    assign _15340 = _15185[46:46];
    assign _15337 = _15332 - _22192;
    assign _15338 = _15334 ? _15337 : _15332;
    assign _15339 = _15338[62:0];
    assign _15341 = { _15339,
                      _15340 };
    assign _15342 = _15341 < _22192;
    assign _15343 = ~ _15342;
    assign _15331 = _15185[47:47];
    assign _15328 = _15323 - _22192;
    assign _15329 = _15325 ? _15328 : _15323;
    assign _15330 = _15329[62:0];
    assign _15332 = { _15330,
                      _15331 };
    assign _15333 = _15332 < _22192;
    assign _15334 = ~ _15333;
    assign _15322 = _15185[48:48];
    assign _15319 = _15314 - _22192;
    assign _15320 = _15316 ? _15319 : _15314;
    assign _15321 = _15320[62:0];
    assign _15323 = { _15321,
                      _15322 };
    assign _15324 = _15323 < _22192;
    assign _15325 = ~ _15324;
    assign _15313 = _15185[49:49];
    assign _15310 = _15305 - _22192;
    assign _15311 = _15307 ? _15310 : _15305;
    assign _15312 = _15311[62:0];
    assign _15314 = { _15312,
                      _15313 };
    assign _15315 = _15314 < _22192;
    assign _15316 = ~ _15315;
    assign _15304 = _15185[50:50];
    assign _15301 = _15296 - _22192;
    assign _15302 = _15298 ? _15301 : _15296;
    assign _15303 = _15302[62:0];
    assign _15305 = { _15303,
                      _15304 };
    assign _15306 = _15305 < _22192;
    assign _15307 = ~ _15306;
    assign _15295 = _15185[51:51];
    assign _15292 = _15287 - _22192;
    assign _15293 = _15289 ? _15292 : _15287;
    assign _15294 = _15293[62:0];
    assign _15296 = { _15294,
                      _15295 };
    assign _15297 = _15296 < _22192;
    assign _15298 = ~ _15297;
    assign _15286 = _15185[52:52];
    assign _15283 = _15278 - _22192;
    assign _15284 = _15280 ? _15283 : _15278;
    assign _15285 = _15284[62:0];
    assign _15287 = { _15285,
                      _15286 };
    assign _15288 = _15287 < _22192;
    assign _15289 = ~ _15288;
    assign _15277 = _15185[53:53];
    assign _15274 = _15269 - _22192;
    assign _15275 = _15271 ? _15274 : _15269;
    assign _15276 = _15275[62:0];
    assign _15278 = { _15276,
                      _15277 };
    assign _15279 = _15278 < _22192;
    assign _15280 = ~ _15279;
    assign _15268 = _15185[54:54];
    assign _15265 = _15260 - _22192;
    assign _15266 = _15262 ? _15265 : _15260;
    assign _15267 = _15266[62:0];
    assign _15269 = { _15267,
                      _15268 };
    assign _15270 = _15269 < _22192;
    assign _15271 = ~ _15270;
    assign _15259 = _15185[55:55];
    assign _15256 = _15251 - _22192;
    assign _15257 = _15253 ? _15256 : _15251;
    assign _15258 = _15257[62:0];
    assign _15260 = { _15258,
                      _15259 };
    assign _15261 = _15260 < _22192;
    assign _15262 = ~ _15261;
    assign _15250 = _15185[56:56];
    assign _15247 = _15242 - _22192;
    assign _15248 = _15244 ? _15247 : _15242;
    assign _15249 = _15248[62:0];
    assign _15251 = { _15249,
                      _15250 };
    assign _15252 = _15251 < _22192;
    assign _15253 = ~ _15252;
    assign _15241 = _15185[57:57];
    assign _15238 = _15233 - _22192;
    assign _15239 = _15235 ? _15238 : _15233;
    assign _15240 = _15239[62:0];
    assign _15242 = { _15240,
                      _15241 };
    assign _15243 = _15242 < _22192;
    assign _15244 = ~ _15243;
    assign _15232 = _15185[58:58];
    assign _15229 = _15224 - _22192;
    assign _15230 = _15226 ? _15229 : _15224;
    assign _15231 = _15230[62:0];
    assign _15233 = { _15231,
                      _15232 };
    assign _15234 = _15233 < _22192;
    assign _15235 = ~ _15234;
    assign _15223 = _15185[59:59];
    assign _15220 = _15215 - _22192;
    assign _15221 = _15217 ? _15220 : _15215;
    assign _15222 = _15221[62:0];
    assign _15224 = { _15222,
                      _15223 };
    assign _15225 = _15224 < _22192;
    assign _15226 = ~ _15225;
    assign _15214 = _15185[60:60];
    assign _15211 = _15206 - _22192;
    assign _15212 = _15208 ? _15211 : _15206;
    assign _15213 = _15212[62:0];
    assign _15215 = { _15213,
                      _15214 };
    assign _15216 = _15215 < _22192;
    assign _15217 = ~ _15216;
    assign _15205 = _15185[61:61];
    assign _15202 = _15197 - _22192;
    assign _15203 = _15199 ? _15202 : _15197;
    assign _15204 = _15203[62:0];
    assign _15206 = { _15204,
                      _15205 };
    assign _15207 = _15206 < _22192;
    assign _15208 = ~ _15207;
    assign _15196 = _15185[62:62];
    assign _15193 = _15187 - _22192;
    assign _15194 = _15190 ? _15193 : _15187;
    assign _15195 = _15194[62:0];
    assign _15197 = { _15195,
                      _15196 };
    assign _15198 = _15197 < _22192;
    assign _15199 = ~ _15198;
    assign _15183 = _15175 + _22186;
    assign _15184 = _15175 * _15183;
    assign _15185 = _15184[63:0];
    assign _15186 = _15185[63:63];
    assign _15187 = { _22185,
                      _15186 };
    assign _15189 = _15187 < _22192;
    assign _15190 = ~ _15189;
    assign _15191 = { _22185,
                      _15190 };
    assign _15192 = _15191[62:0];
    assign _15200 = { _15192,
                      _15199 };
    assign _15201 = _15200[62:0];
    assign _15209 = { _15201,
                      _15208 };
    assign _15210 = _15209[62:0];
    assign _15218 = { _15210,
                      _15217 };
    assign _15219 = _15218[62:0];
    assign _15227 = { _15219,
                      _15226 };
    assign _15228 = _15227[62:0];
    assign _15236 = { _15228,
                      _15235 };
    assign _15237 = _15236[62:0];
    assign _15245 = { _15237,
                      _15244 };
    assign _15246 = _15245[62:0];
    assign _15254 = { _15246,
                      _15253 };
    assign _15255 = _15254[62:0];
    assign _15263 = { _15255,
                      _15262 };
    assign _15264 = _15263[62:0];
    assign _15272 = { _15264,
                      _15271 };
    assign _15273 = _15272[62:0];
    assign _15281 = { _15273,
                      _15280 };
    assign _15282 = _15281[62:0];
    assign _15290 = { _15282,
                      _15289 };
    assign _15291 = _15290[62:0];
    assign _15299 = { _15291,
                      _15298 };
    assign _15300 = _15299[62:0];
    assign _15308 = { _15300,
                      _15307 };
    assign _15309 = _15308[62:0];
    assign _15317 = { _15309,
                      _15316 };
    assign _15318 = _15317[62:0];
    assign _15326 = { _15318,
                      _15325 };
    assign _15327 = _15326[62:0];
    assign _15335 = { _15327,
                      _15334 };
    assign _15336 = _15335[62:0];
    assign _15344 = { _15336,
                      _15343 };
    assign _15345 = _15344[62:0];
    assign _15353 = { _15345,
                      _15352 };
    assign _15354 = _15353[62:0];
    assign _15362 = { _15354,
                      _15361 };
    assign _15363 = _15362[62:0];
    assign _15371 = { _15363,
                      _15370 };
    assign _15372 = _15371[62:0];
    assign _15380 = { _15372,
                      _15379 };
    assign _15381 = _15380[62:0];
    assign _15389 = { _15381,
                      _15388 };
    assign _15390 = _15389[62:0];
    assign _15398 = { _15390,
                      _15397 };
    assign _15399 = _15398[62:0];
    assign _15407 = { _15399,
                      _15406 };
    assign _15408 = _15407[62:0];
    assign _15416 = { _15408,
                      _15415 };
    assign _15417 = _15416[62:0];
    assign _15425 = { _15417,
                      _15424 };
    assign _15426 = _15425[62:0];
    assign _15434 = { _15426,
                      _15433 };
    assign _15435 = _15434[62:0];
    assign _15443 = { _15435,
                      _15442 };
    assign _15444 = _15443[62:0];
    assign _15452 = { _15444,
                      _15451 };
    assign _15453 = _15452[62:0];
    assign _15461 = { _15453,
                      _15460 };
    assign _15462 = _15461[62:0];
    assign _15470 = { _15462,
                      _15469 };
    assign _15471 = _15470[62:0];
    assign _15479 = { _15471,
                      _15478 };
    assign _15480 = _15479[62:0];
    assign _15488 = { _15480,
                      _15487 };
    assign _15489 = _15488[62:0];
    assign _15497 = { _15489,
                      _15496 };
    assign _15498 = _15497[62:0];
    assign _15506 = { _15498,
                      _15505 };
    assign _15507 = _15506[62:0];
    assign _15515 = { _15507,
                      _15514 };
    assign _15516 = _15515[62:0];
    assign _15524 = { _15516,
                      _15523 };
    assign _15525 = _15524[62:0];
    assign _15533 = { _15525,
                      _15532 };
    assign _15534 = _15533[62:0];
    assign _15542 = { _15534,
                      _15541 };
    assign _15543 = _15542[62:0];
    assign _15551 = { _15543,
                      _15550 };
    assign _15552 = _15551[62:0];
    assign _15560 = { _15552,
                      _15559 };
    assign _15561 = _15560[62:0];
    assign _15569 = { _15561,
                      _15568 };
    assign _15570 = _15569[62:0];
    assign _15578 = { _15570,
                      _15577 };
    assign _15579 = _15578[62:0];
    assign _15587 = { _15579,
                      _15586 };
    assign _15588 = _15587[62:0];
    assign _15596 = { _15588,
                      _15595 };
    assign _15597 = _15596[62:0];
    assign _15605 = { _15597,
                      _15604 };
    assign _15606 = _15605[62:0];
    assign _15614 = { _15606,
                      _15613 };
    assign _15615 = _15614[62:0];
    assign _15623 = { _15615,
                      _15622 };
    assign _15624 = _15623[62:0];
    assign _15632 = { _15624,
                      _15631 };
    assign _15633 = _15632[62:0];
    assign _15641 = { _15633,
                      _15640 };
    assign _15642 = _15641[62:0];
    assign _15650 = { _15642,
                      _15649 };
    assign _15651 = _15650[62:0];
    assign _15659 = { _15651,
                      _15658 };
    assign _15660 = _15659[62:0];
    assign _15668 = { _15660,
                      _15667 };
    assign _15669 = _15668[62:0];
    assign _15677 = { _15669,
                      _15676 };
    assign _15678 = _15677[62:0];
    assign _15686 = { _15678,
                      _15685 };
    assign _15687 = _15686[62:0];
    assign _15695 = { _15687,
                      _15694 };
    assign _15696 = _15695[62:0];
    assign _15704 = { _15696,
                      _15703 };
    assign _15705 = _15704[62:0];
    assign _15713 = { _15705,
                      _15712 };
    assign _15714 = _15713[62:0];
    assign _15722 = { _15714,
                      _15721 };
    assign _15723 = _15722[62:0];
    assign _15731 = { _15723,
                      _15730 };
    assign _15732 = _15731[62:0];
    assign _15740 = { _15732,
                      _15739 };
    assign _15741 = _15740[62:0];
    assign _15749 = { _15741,
                      _15748 };
    assign _15750 = _15749[62:0];
    assign _15758 = { _15750,
                      _15757 };
    assign _15759 = _14023 * _15758;
    assign _15760 = _15759[63:0];
    assign _15171 = _14603[0:0];
    assign _15168 = _15163 - _14023;
    assign _15169 = _15165 ? _15168 : _15163;
    assign _15170 = _15169[62:0];
    assign _15172 = { _15170,
                      _15171 };
    assign _15173 = _15172 < _14023;
    assign _15174 = ~ _15173;
    assign _15162 = _14603[1:1];
    assign _15159 = _15154 - _14023;
    assign _15160 = _15156 ? _15159 : _15154;
    assign _15161 = _15160[62:0];
    assign _15163 = { _15161,
                      _15162 };
    assign _15164 = _15163 < _14023;
    assign _15165 = ~ _15164;
    assign _15153 = _14603[2:2];
    assign _15150 = _15145 - _14023;
    assign _15151 = _15147 ? _15150 : _15145;
    assign _15152 = _15151[62:0];
    assign _15154 = { _15152,
                      _15153 };
    assign _15155 = _15154 < _14023;
    assign _15156 = ~ _15155;
    assign _15144 = _14603[3:3];
    assign _15141 = _15136 - _14023;
    assign _15142 = _15138 ? _15141 : _15136;
    assign _15143 = _15142[62:0];
    assign _15145 = { _15143,
                      _15144 };
    assign _15146 = _15145 < _14023;
    assign _15147 = ~ _15146;
    assign _15135 = _14603[4:4];
    assign _15132 = _15127 - _14023;
    assign _15133 = _15129 ? _15132 : _15127;
    assign _15134 = _15133[62:0];
    assign _15136 = { _15134,
                      _15135 };
    assign _15137 = _15136 < _14023;
    assign _15138 = ~ _15137;
    assign _15126 = _14603[5:5];
    assign _15123 = _15118 - _14023;
    assign _15124 = _15120 ? _15123 : _15118;
    assign _15125 = _15124[62:0];
    assign _15127 = { _15125,
                      _15126 };
    assign _15128 = _15127 < _14023;
    assign _15129 = ~ _15128;
    assign _15117 = _14603[6:6];
    assign _15114 = _15109 - _14023;
    assign _15115 = _15111 ? _15114 : _15109;
    assign _15116 = _15115[62:0];
    assign _15118 = { _15116,
                      _15117 };
    assign _15119 = _15118 < _14023;
    assign _15120 = ~ _15119;
    assign _15108 = _14603[7:7];
    assign _15105 = _15100 - _14023;
    assign _15106 = _15102 ? _15105 : _15100;
    assign _15107 = _15106[62:0];
    assign _15109 = { _15107,
                      _15108 };
    assign _15110 = _15109 < _14023;
    assign _15111 = ~ _15110;
    assign _15099 = _14603[8:8];
    assign _15096 = _15091 - _14023;
    assign _15097 = _15093 ? _15096 : _15091;
    assign _15098 = _15097[62:0];
    assign _15100 = { _15098,
                      _15099 };
    assign _15101 = _15100 < _14023;
    assign _15102 = ~ _15101;
    assign _15090 = _14603[9:9];
    assign _15087 = _15082 - _14023;
    assign _15088 = _15084 ? _15087 : _15082;
    assign _15089 = _15088[62:0];
    assign _15091 = { _15089,
                      _15090 };
    assign _15092 = _15091 < _14023;
    assign _15093 = ~ _15092;
    assign _15081 = _14603[10:10];
    assign _15078 = _15073 - _14023;
    assign _15079 = _15075 ? _15078 : _15073;
    assign _15080 = _15079[62:0];
    assign _15082 = { _15080,
                      _15081 };
    assign _15083 = _15082 < _14023;
    assign _15084 = ~ _15083;
    assign _15072 = _14603[11:11];
    assign _15069 = _15064 - _14023;
    assign _15070 = _15066 ? _15069 : _15064;
    assign _15071 = _15070[62:0];
    assign _15073 = { _15071,
                      _15072 };
    assign _15074 = _15073 < _14023;
    assign _15075 = ~ _15074;
    assign _15063 = _14603[12:12];
    assign _15060 = _15055 - _14023;
    assign _15061 = _15057 ? _15060 : _15055;
    assign _15062 = _15061[62:0];
    assign _15064 = { _15062,
                      _15063 };
    assign _15065 = _15064 < _14023;
    assign _15066 = ~ _15065;
    assign _15054 = _14603[13:13];
    assign _15051 = _15046 - _14023;
    assign _15052 = _15048 ? _15051 : _15046;
    assign _15053 = _15052[62:0];
    assign _15055 = { _15053,
                      _15054 };
    assign _15056 = _15055 < _14023;
    assign _15057 = ~ _15056;
    assign _15045 = _14603[14:14];
    assign _15042 = _15037 - _14023;
    assign _15043 = _15039 ? _15042 : _15037;
    assign _15044 = _15043[62:0];
    assign _15046 = { _15044,
                      _15045 };
    assign _15047 = _15046 < _14023;
    assign _15048 = ~ _15047;
    assign _15036 = _14603[15:15];
    assign _15033 = _15028 - _14023;
    assign _15034 = _15030 ? _15033 : _15028;
    assign _15035 = _15034[62:0];
    assign _15037 = { _15035,
                      _15036 };
    assign _15038 = _15037 < _14023;
    assign _15039 = ~ _15038;
    assign _15027 = _14603[16:16];
    assign _15024 = _15019 - _14023;
    assign _15025 = _15021 ? _15024 : _15019;
    assign _15026 = _15025[62:0];
    assign _15028 = { _15026,
                      _15027 };
    assign _15029 = _15028 < _14023;
    assign _15030 = ~ _15029;
    assign _15018 = _14603[17:17];
    assign _15015 = _15010 - _14023;
    assign _15016 = _15012 ? _15015 : _15010;
    assign _15017 = _15016[62:0];
    assign _15019 = { _15017,
                      _15018 };
    assign _15020 = _15019 < _14023;
    assign _15021 = ~ _15020;
    assign _15009 = _14603[18:18];
    assign _15006 = _15001 - _14023;
    assign _15007 = _15003 ? _15006 : _15001;
    assign _15008 = _15007[62:0];
    assign _15010 = { _15008,
                      _15009 };
    assign _15011 = _15010 < _14023;
    assign _15012 = ~ _15011;
    assign _15000 = _14603[19:19];
    assign _14997 = _14992 - _14023;
    assign _14998 = _14994 ? _14997 : _14992;
    assign _14999 = _14998[62:0];
    assign _15001 = { _14999,
                      _15000 };
    assign _15002 = _15001 < _14023;
    assign _15003 = ~ _15002;
    assign _14991 = _14603[20:20];
    assign _14988 = _14983 - _14023;
    assign _14989 = _14985 ? _14988 : _14983;
    assign _14990 = _14989[62:0];
    assign _14992 = { _14990,
                      _14991 };
    assign _14993 = _14992 < _14023;
    assign _14994 = ~ _14993;
    assign _14982 = _14603[21:21];
    assign _14979 = _14974 - _14023;
    assign _14980 = _14976 ? _14979 : _14974;
    assign _14981 = _14980[62:0];
    assign _14983 = { _14981,
                      _14982 };
    assign _14984 = _14983 < _14023;
    assign _14985 = ~ _14984;
    assign _14973 = _14603[22:22];
    assign _14970 = _14965 - _14023;
    assign _14971 = _14967 ? _14970 : _14965;
    assign _14972 = _14971[62:0];
    assign _14974 = { _14972,
                      _14973 };
    assign _14975 = _14974 < _14023;
    assign _14976 = ~ _14975;
    assign _14964 = _14603[23:23];
    assign _14961 = _14956 - _14023;
    assign _14962 = _14958 ? _14961 : _14956;
    assign _14963 = _14962[62:0];
    assign _14965 = { _14963,
                      _14964 };
    assign _14966 = _14965 < _14023;
    assign _14967 = ~ _14966;
    assign _14955 = _14603[24:24];
    assign _14952 = _14947 - _14023;
    assign _14953 = _14949 ? _14952 : _14947;
    assign _14954 = _14953[62:0];
    assign _14956 = { _14954,
                      _14955 };
    assign _14957 = _14956 < _14023;
    assign _14958 = ~ _14957;
    assign _14946 = _14603[25:25];
    assign _14943 = _14938 - _14023;
    assign _14944 = _14940 ? _14943 : _14938;
    assign _14945 = _14944[62:0];
    assign _14947 = { _14945,
                      _14946 };
    assign _14948 = _14947 < _14023;
    assign _14949 = ~ _14948;
    assign _14937 = _14603[26:26];
    assign _14934 = _14929 - _14023;
    assign _14935 = _14931 ? _14934 : _14929;
    assign _14936 = _14935[62:0];
    assign _14938 = { _14936,
                      _14937 };
    assign _14939 = _14938 < _14023;
    assign _14940 = ~ _14939;
    assign _14928 = _14603[27:27];
    assign _14925 = _14920 - _14023;
    assign _14926 = _14922 ? _14925 : _14920;
    assign _14927 = _14926[62:0];
    assign _14929 = { _14927,
                      _14928 };
    assign _14930 = _14929 < _14023;
    assign _14931 = ~ _14930;
    assign _14919 = _14603[28:28];
    assign _14916 = _14911 - _14023;
    assign _14917 = _14913 ? _14916 : _14911;
    assign _14918 = _14917[62:0];
    assign _14920 = { _14918,
                      _14919 };
    assign _14921 = _14920 < _14023;
    assign _14922 = ~ _14921;
    assign _14910 = _14603[29:29];
    assign _14907 = _14902 - _14023;
    assign _14908 = _14904 ? _14907 : _14902;
    assign _14909 = _14908[62:0];
    assign _14911 = { _14909,
                      _14910 };
    assign _14912 = _14911 < _14023;
    assign _14913 = ~ _14912;
    assign _14901 = _14603[30:30];
    assign _14898 = _14893 - _14023;
    assign _14899 = _14895 ? _14898 : _14893;
    assign _14900 = _14899[62:0];
    assign _14902 = { _14900,
                      _14901 };
    assign _14903 = _14902 < _14023;
    assign _14904 = ~ _14903;
    assign _14892 = _14603[31:31];
    assign _14889 = _14884 - _14023;
    assign _14890 = _14886 ? _14889 : _14884;
    assign _14891 = _14890[62:0];
    assign _14893 = { _14891,
                      _14892 };
    assign _14894 = _14893 < _14023;
    assign _14895 = ~ _14894;
    assign _14883 = _14603[32:32];
    assign _14880 = _14875 - _14023;
    assign _14881 = _14877 ? _14880 : _14875;
    assign _14882 = _14881[62:0];
    assign _14884 = { _14882,
                      _14883 };
    assign _14885 = _14884 < _14023;
    assign _14886 = ~ _14885;
    assign _14874 = _14603[33:33];
    assign _14871 = _14866 - _14023;
    assign _14872 = _14868 ? _14871 : _14866;
    assign _14873 = _14872[62:0];
    assign _14875 = { _14873,
                      _14874 };
    assign _14876 = _14875 < _14023;
    assign _14877 = ~ _14876;
    assign _14865 = _14603[34:34];
    assign _14862 = _14857 - _14023;
    assign _14863 = _14859 ? _14862 : _14857;
    assign _14864 = _14863[62:0];
    assign _14866 = { _14864,
                      _14865 };
    assign _14867 = _14866 < _14023;
    assign _14868 = ~ _14867;
    assign _14856 = _14603[35:35];
    assign _14853 = _14848 - _14023;
    assign _14854 = _14850 ? _14853 : _14848;
    assign _14855 = _14854[62:0];
    assign _14857 = { _14855,
                      _14856 };
    assign _14858 = _14857 < _14023;
    assign _14859 = ~ _14858;
    assign _14847 = _14603[36:36];
    assign _14844 = _14839 - _14023;
    assign _14845 = _14841 ? _14844 : _14839;
    assign _14846 = _14845[62:0];
    assign _14848 = { _14846,
                      _14847 };
    assign _14849 = _14848 < _14023;
    assign _14850 = ~ _14849;
    assign _14838 = _14603[37:37];
    assign _14835 = _14830 - _14023;
    assign _14836 = _14832 ? _14835 : _14830;
    assign _14837 = _14836[62:0];
    assign _14839 = { _14837,
                      _14838 };
    assign _14840 = _14839 < _14023;
    assign _14841 = ~ _14840;
    assign _14829 = _14603[38:38];
    assign _14826 = _14821 - _14023;
    assign _14827 = _14823 ? _14826 : _14821;
    assign _14828 = _14827[62:0];
    assign _14830 = { _14828,
                      _14829 };
    assign _14831 = _14830 < _14023;
    assign _14832 = ~ _14831;
    assign _14820 = _14603[39:39];
    assign _14817 = _14812 - _14023;
    assign _14818 = _14814 ? _14817 : _14812;
    assign _14819 = _14818[62:0];
    assign _14821 = { _14819,
                      _14820 };
    assign _14822 = _14821 < _14023;
    assign _14823 = ~ _14822;
    assign _14811 = _14603[40:40];
    assign _14808 = _14803 - _14023;
    assign _14809 = _14805 ? _14808 : _14803;
    assign _14810 = _14809[62:0];
    assign _14812 = { _14810,
                      _14811 };
    assign _14813 = _14812 < _14023;
    assign _14814 = ~ _14813;
    assign _14802 = _14603[41:41];
    assign _14799 = _14794 - _14023;
    assign _14800 = _14796 ? _14799 : _14794;
    assign _14801 = _14800[62:0];
    assign _14803 = { _14801,
                      _14802 };
    assign _14804 = _14803 < _14023;
    assign _14805 = ~ _14804;
    assign _14793 = _14603[42:42];
    assign _14790 = _14785 - _14023;
    assign _14791 = _14787 ? _14790 : _14785;
    assign _14792 = _14791[62:0];
    assign _14794 = { _14792,
                      _14793 };
    assign _14795 = _14794 < _14023;
    assign _14796 = ~ _14795;
    assign _14784 = _14603[43:43];
    assign _14781 = _14776 - _14023;
    assign _14782 = _14778 ? _14781 : _14776;
    assign _14783 = _14782[62:0];
    assign _14785 = { _14783,
                      _14784 };
    assign _14786 = _14785 < _14023;
    assign _14787 = ~ _14786;
    assign _14775 = _14603[44:44];
    assign _14772 = _14767 - _14023;
    assign _14773 = _14769 ? _14772 : _14767;
    assign _14774 = _14773[62:0];
    assign _14776 = { _14774,
                      _14775 };
    assign _14777 = _14776 < _14023;
    assign _14778 = ~ _14777;
    assign _14766 = _14603[45:45];
    assign _14763 = _14758 - _14023;
    assign _14764 = _14760 ? _14763 : _14758;
    assign _14765 = _14764[62:0];
    assign _14767 = { _14765,
                      _14766 };
    assign _14768 = _14767 < _14023;
    assign _14769 = ~ _14768;
    assign _14757 = _14603[46:46];
    assign _14754 = _14749 - _14023;
    assign _14755 = _14751 ? _14754 : _14749;
    assign _14756 = _14755[62:0];
    assign _14758 = { _14756,
                      _14757 };
    assign _14759 = _14758 < _14023;
    assign _14760 = ~ _14759;
    assign _14748 = _14603[47:47];
    assign _14745 = _14740 - _14023;
    assign _14746 = _14742 ? _14745 : _14740;
    assign _14747 = _14746[62:0];
    assign _14749 = { _14747,
                      _14748 };
    assign _14750 = _14749 < _14023;
    assign _14751 = ~ _14750;
    assign _14739 = _14603[48:48];
    assign _14736 = _14731 - _14023;
    assign _14737 = _14733 ? _14736 : _14731;
    assign _14738 = _14737[62:0];
    assign _14740 = { _14738,
                      _14739 };
    assign _14741 = _14740 < _14023;
    assign _14742 = ~ _14741;
    assign _14730 = _14603[49:49];
    assign _14727 = _14722 - _14023;
    assign _14728 = _14724 ? _14727 : _14722;
    assign _14729 = _14728[62:0];
    assign _14731 = { _14729,
                      _14730 };
    assign _14732 = _14731 < _14023;
    assign _14733 = ~ _14732;
    assign _14721 = _14603[50:50];
    assign _14718 = _14713 - _14023;
    assign _14719 = _14715 ? _14718 : _14713;
    assign _14720 = _14719[62:0];
    assign _14722 = { _14720,
                      _14721 };
    assign _14723 = _14722 < _14023;
    assign _14724 = ~ _14723;
    assign _14712 = _14603[51:51];
    assign _14709 = _14704 - _14023;
    assign _14710 = _14706 ? _14709 : _14704;
    assign _14711 = _14710[62:0];
    assign _14713 = { _14711,
                      _14712 };
    assign _14714 = _14713 < _14023;
    assign _14715 = ~ _14714;
    assign _14703 = _14603[52:52];
    assign _14700 = _14695 - _14023;
    assign _14701 = _14697 ? _14700 : _14695;
    assign _14702 = _14701[62:0];
    assign _14704 = { _14702,
                      _14703 };
    assign _14705 = _14704 < _14023;
    assign _14706 = ~ _14705;
    assign _14694 = _14603[53:53];
    assign _14691 = _14686 - _14023;
    assign _14692 = _14688 ? _14691 : _14686;
    assign _14693 = _14692[62:0];
    assign _14695 = { _14693,
                      _14694 };
    assign _14696 = _14695 < _14023;
    assign _14697 = ~ _14696;
    assign _14685 = _14603[54:54];
    assign _14682 = _14677 - _14023;
    assign _14683 = _14679 ? _14682 : _14677;
    assign _14684 = _14683[62:0];
    assign _14686 = { _14684,
                      _14685 };
    assign _14687 = _14686 < _14023;
    assign _14688 = ~ _14687;
    assign _14676 = _14603[55:55];
    assign _14673 = _14668 - _14023;
    assign _14674 = _14670 ? _14673 : _14668;
    assign _14675 = _14674[62:0];
    assign _14677 = { _14675,
                      _14676 };
    assign _14678 = _14677 < _14023;
    assign _14679 = ~ _14678;
    assign _14667 = _14603[56:56];
    assign _14664 = _14659 - _14023;
    assign _14665 = _14661 ? _14664 : _14659;
    assign _14666 = _14665[62:0];
    assign _14668 = { _14666,
                      _14667 };
    assign _14669 = _14668 < _14023;
    assign _14670 = ~ _14669;
    assign _14658 = _14603[57:57];
    assign _14655 = _14650 - _14023;
    assign _14656 = _14652 ? _14655 : _14650;
    assign _14657 = _14656[62:0];
    assign _14659 = { _14657,
                      _14658 };
    assign _14660 = _14659 < _14023;
    assign _14661 = ~ _14660;
    assign _14649 = _14603[58:58];
    assign _14646 = _14641 - _14023;
    assign _14647 = _14643 ? _14646 : _14641;
    assign _14648 = _14647[62:0];
    assign _14650 = { _14648,
                      _14649 };
    assign _14651 = _14650 < _14023;
    assign _14652 = ~ _14651;
    assign _14640 = _14603[59:59];
    assign _14637 = _14632 - _14023;
    assign _14638 = _14634 ? _14637 : _14632;
    assign _14639 = _14638[62:0];
    assign _14641 = { _14639,
                      _14640 };
    assign _14642 = _14641 < _14023;
    assign _14643 = ~ _14642;
    assign _14631 = _14603[60:60];
    assign _14628 = _14623 - _14023;
    assign _14629 = _14625 ? _14628 : _14623;
    assign _14630 = _14629[62:0];
    assign _14632 = { _14630,
                      _14631 };
    assign _14633 = _14632 < _14023;
    assign _14634 = ~ _14633;
    assign _14622 = _14603[61:61];
    assign _14619 = _14614 - _14023;
    assign _14620 = _14616 ? _14619 : _14614;
    assign _14621 = _14620[62:0];
    assign _14623 = { _14621,
                      _14622 };
    assign _14624 = _14623 < _14023;
    assign _14625 = ~ _14624;
    assign _14613 = _14603[62:62];
    assign _14610 = _14605 - _14023;
    assign _14611 = _14607 ? _14610 : _14605;
    assign _14612 = _14611[62:0];
    assign _14614 = { _14612,
                      _14613 };
    assign _14615 = _14614 < _14023;
    assign _14616 = ~ _14615;
    assign _14603 = _14015 - _14597;
    assign _14604 = _14603[63:63];
    assign _14605 = { _22185,
                      _14604 };
    assign _14606 = _14605 < _14023;
    assign _14607 = ~ _14606;
    assign _14608 = { _22185,
                      _14607 };
    assign _14609 = _14608[62:0];
    assign _14617 = { _14609,
                      _14616 };
    assign _14618 = _14617[62:0];
    assign _14626 = { _14618,
                      _14625 };
    assign _14627 = _14626[62:0];
    assign _14635 = { _14627,
                      _14634 };
    assign _14636 = _14635[62:0];
    assign _14644 = { _14636,
                      _14643 };
    assign _14645 = _14644[62:0];
    assign _14653 = { _14645,
                      _14652 };
    assign _14654 = _14653[62:0];
    assign _14662 = { _14654,
                      _14661 };
    assign _14663 = _14662[62:0];
    assign _14671 = { _14663,
                      _14670 };
    assign _14672 = _14671[62:0];
    assign _14680 = { _14672,
                      _14679 };
    assign _14681 = _14680[62:0];
    assign _14689 = { _14681,
                      _14688 };
    assign _14690 = _14689[62:0];
    assign _14698 = { _14690,
                      _14697 };
    assign _14699 = _14698[62:0];
    assign _14707 = { _14699,
                      _14706 };
    assign _14708 = _14707[62:0];
    assign _14716 = { _14708,
                      _14715 };
    assign _14717 = _14716[62:0];
    assign _14725 = { _14717,
                      _14724 };
    assign _14726 = _14725[62:0];
    assign _14734 = { _14726,
                      _14733 };
    assign _14735 = _14734[62:0];
    assign _14743 = { _14735,
                      _14742 };
    assign _14744 = _14743[62:0];
    assign _14752 = { _14744,
                      _14751 };
    assign _14753 = _14752[62:0];
    assign _14761 = { _14753,
                      _14760 };
    assign _14762 = _14761[62:0];
    assign _14770 = { _14762,
                      _14769 };
    assign _14771 = _14770[62:0];
    assign _14779 = { _14771,
                      _14778 };
    assign _14780 = _14779[62:0];
    assign _14788 = { _14780,
                      _14787 };
    assign _14789 = _14788[62:0];
    assign _14797 = { _14789,
                      _14796 };
    assign _14798 = _14797[62:0];
    assign _14806 = { _14798,
                      _14805 };
    assign _14807 = _14806[62:0];
    assign _14815 = { _14807,
                      _14814 };
    assign _14816 = _14815[62:0];
    assign _14824 = { _14816,
                      _14823 };
    assign _14825 = _14824[62:0];
    assign _14833 = { _14825,
                      _14832 };
    assign _14834 = _14833[62:0];
    assign _14842 = { _14834,
                      _14841 };
    assign _14843 = _14842[62:0];
    assign _14851 = { _14843,
                      _14850 };
    assign _14852 = _14851[62:0];
    assign _14860 = { _14852,
                      _14859 };
    assign _14861 = _14860[62:0];
    assign _14869 = { _14861,
                      _14868 };
    assign _14870 = _14869[62:0];
    assign _14878 = { _14870,
                      _14877 };
    assign _14879 = _14878[62:0];
    assign _14887 = { _14879,
                      _14886 };
    assign _14888 = _14887[62:0];
    assign _14896 = { _14888,
                      _14895 };
    assign _14897 = _14896[62:0];
    assign _14905 = { _14897,
                      _14904 };
    assign _14906 = _14905[62:0];
    assign _14914 = { _14906,
                      _14913 };
    assign _14915 = _14914[62:0];
    assign _14923 = { _14915,
                      _14922 };
    assign _14924 = _14923[62:0];
    assign _14932 = { _14924,
                      _14931 };
    assign _14933 = _14932[62:0];
    assign _14941 = { _14933,
                      _14940 };
    assign _14942 = _14941[62:0];
    assign _14950 = { _14942,
                      _14949 };
    assign _14951 = _14950[62:0];
    assign _14959 = { _14951,
                      _14958 };
    assign _14960 = _14959[62:0];
    assign _14968 = { _14960,
                      _14967 };
    assign _14969 = _14968[62:0];
    assign _14977 = { _14969,
                      _14976 };
    assign _14978 = _14977[62:0];
    assign _14986 = { _14978,
                      _14985 };
    assign _14987 = _14986[62:0];
    assign _14995 = { _14987,
                      _14994 };
    assign _14996 = _14995[62:0];
    assign _15004 = { _14996,
                      _15003 };
    assign _15005 = _15004[62:0];
    assign _15013 = { _15005,
                      _15012 };
    assign _15014 = _15013[62:0];
    assign _15022 = { _15014,
                      _15021 };
    assign _15023 = _15022[62:0];
    assign _15031 = { _15023,
                      _15030 };
    assign _15032 = _15031[62:0];
    assign _15040 = { _15032,
                      _15039 };
    assign _15041 = _15040[62:0];
    assign _15049 = { _15041,
                      _15048 };
    assign _15050 = _15049[62:0];
    assign _15058 = { _15050,
                      _15057 };
    assign _15059 = _15058[62:0];
    assign _15067 = { _15059,
                      _15066 };
    assign _15068 = _15067[62:0];
    assign _15076 = { _15068,
                      _15075 };
    assign _15077 = _15076[62:0];
    assign _15085 = { _15077,
                      _15084 };
    assign _15086 = _15085[62:0];
    assign _15094 = { _15086,
                      _15093 };
    assign _15095 = _15094[62:0];
    assign _15103 = { _15095,
                      _15102 };
    assign _15104 = _15103[62:0];
    assign _15112 = { _15104,
                      _15111 };
    assign _15113 = _15112[62:0];
    assign _15121 = { _15113,
                      _15120 };
    assign _15122 = _15121[62:0];
    assign _15130 = { _15122,
                      _15129 };
    assign _15131 = _15130[62:0];
    assign _15139 = { _15131,
                      _15138 };
    assign _15140 = _15139[62:0];
    assign _15148 = { _15140,
                      _15147 };
    assign _15149 = _15148[62:0];
    assign _15157 = { _15149,
                      _15156 };
    assign _15158 = _15157[62:0];
    assign _15166 = { _15158,
                      _15165 };
    assign _15167 = _15166[62:0];
    assign _15175 = { _15167,
                      _15174 };
    assign _15177 = _15175 + _22186;
    assign _15178 = _15177 * _14597;
    assign _15179 = _15178[63:0];
    assign _15761 = _15179 + _15760;
    assign _14589 = _14020[0:0];
    assign _14586 = _14581 - _14023;
    assign _14587 = _14583 ? _14586 : _14581;
    assign _14588 = _14587[62:0];
    assign _14590 = { _14588,
                      _14589 };
    assign _14591 = _14590 < _14023;
    assign _14592 = ~ _14591;
    assign _14580 = _14020[1:1];
    assign _14577 = _14572 - _14023;
    assign _14578 = _14574 ? _14577 : _14572;
    assign _14579 = _14578[62:0];
    assign _14581 = { _14579,
                      _14580 };
    assign _14582 = _14581 < _14023;
    assign _14583 = ~ _14582;
    assign _14571 = _14020[2:2];
    assign _14568 = _14563 - _14023;
    assign _14569 = _14565 ? _14568 : _14563;
    assign _14570 = _14569[62:0];
    assign _14572 = { _14570,
                      _14571 };
    assign _14573 = _14572 < _14023;
    assign _14574 = ~ _14573;
    assign _14562 = _14020[3:3];
    assign _14559 = _14554 - _14023;
    assign _14560 = _14556 ? _14559 : _14554;
    assign _14561 = _14560[62:0];
    assign _14563 = { _14561,
                      _14562 };
    assign _14564 = _14563 < _14023;
    assign _14565 = ~ _14564;
    assign _14553 = _14020[4:4];
    assign _14550 = _14545 - _14023;
    assign _14551 = _14547 ? _14550 : _14545;
    assign _14552 = _14551[62:0];
    assign _14554 = { _14552,
                      _14553 };
    assign _14555 = _14554 < _14023;
    assign _14556 = ~ _14555;
    assign _14544 = _14020[5:5];
    assign _14541 = _14536 - _14023;
    assign _14542 = _14538 ? _14541 : _14536;
    assign _14543 = _14542[62:0];
    assign _14545 = { _14543,
                      _14544 };
    assign _14546 = _14545 < _14023;
    assign _14547 = ~ _14546;
    assign _14535 = _14020[6:6];
    assign _14532 = _14527 - _14023;
    assign _14533 = _14529 ? _14532 : _14527;
    assign _14534 = _14533[62:0];
    assign _14536 = { _14534,
                      _14535 };
    assign _14537 = _14536 < _14023;
    assign _14538 = ~ _14537;
    assign _14526 = _14020[7:7];
    assign _14523 = _14518 - _14023;
    assign _14524 = _14520 ? _14523 : _14518;
    assign _14525 = _14524[62:0];
    assign _14527 = { _14525,
                      _14526 };
    assign _14528 = _14527 < _14023;
    assign _14529 = ~ _14528;
    assign _14517 = _14020[8:8];
    assign _14514 = _14509 - _14023;
    assign _14515 = _14511 ? _14514 : _14509;
    assign _14516 = _14515[62:0];
    assign _14518 = { _14516,
                      _14517 };
    assign _14519 = _14518 < _14023;
    assign _14520 = ~ _14519;
    assign _14508 = _14020[9:9];
    assign _14505 = _14500 - _14023;
    assign _14506 = _14502 ? _14505 : _14500;
    assign _14507 = _14506[62:0];
    assign _14509 = { _14507,
                      _14508 };
    assign _14510 = _14509 < _14023;
    assign _14511 = ~ _14510;
    assign _14499 = _14020[10:10];
    assign _14496 = _14491 - _14023;
    assign _14497 = _14493 ? _14496 : _14491;
    assign _14498 = _14497[62:0];
    assign _14500 = { _14498,
                      _14499 };
    assign _14501 = _14500 < _14023;
    assign _14502 = ~ _14501;
    assign _14490 = _14020[11:11];
    assign _14487 = _14482 - _14023;
    assign _14488 = _14484 ? _14487 : _14482;
    assign _14489 = _14488[62:0];
    assign _14491 = { _14489,
                      _14490 };
    assign _14492 = _14491 < _14023;
    assign _14493 = ~ _14492;
    assign _14481 = _14020[12:12];
    assign _14478 = _14473 - _14023;
    assign _14479 = _14475 ? _14478 : _14473;
    assign _14480 = _14479[62:0];
    assign _14482 = { _14480,
                      _14481 };
    assign _14483 = _14482 < _14023;
    assign _14484 = ~ _14483;
    assign _14472 = _14020[13:13];
    assign _14469 = _14464 - _14023;
    assign _14470 = _14466 ? _14469 : _14464;
    assign _14471 = _14470[62:0];
    assign _14473 = { _14471,
                      _14472 };
    assign _14474 = _14473 < _14023;
    assign _14475 = ~ _14474;
    assign _14463 = _14020[14:14];
    assign _14460 = _14455 - _14023;
    assign _14461 = _14457 ? _14460 : _14455;
    assign _14462 = _14461[62:0];
    assign _14464 = { _14462,
                      _14463 };
    assign _14465 = _14464 < _14023;
    assign _14466 = ~ _14465;
    assign _14454 = _14020[15:15];
    assign _14451 = _14446 - _14023;
    assign _14452 = _14448 ? _14451 : _14446;
    assign _14453 = _14452[62:0];
    assign _14455 = { _14453,
                      _14454 };
    assign _14456 = _14455 < _14023;
    assign _14457 = ~ _14456;
    assign _14445 = _14020[16:16];
    assign _14442 = _14437 - _14023;
    assign _14443 = _14439 ? _14442 : _14437;
    assign _14444 = _14443[62:0];
    assign _14446 = { _14444,
                      _14445 };
    assign _14447 = _14446 < _14023;
    assign _14448 = ~ _14447;
    assign _14436 = _14020[17:17];
    assign _14433 = _14428 - _14023;
    assign _14434 = _14430 ? _14433 : _14428;
    assign _14435 = _14434[62:0];
    assign _14437 = { _14435,
                      _14436 };
    assign _14438 = _14437 < _14023;
    assign _14439 = ~ _14438;
    assign _14427 = _14020[18:18];
    assign _14424 = _14419 - _14023;
    assign _14425 = _14421 ? _14424 : _14419;
    assign _14426 = _14425[62:0];
    assign _14428 = { _14426,
                      _14427 };
    assign _14429 = _14428 < _14023;
    assign _14430 = ~ _14429;
    assign _14418 = _14020[19:19];
    assign _14415 = _14410 - _14023;
    assign _14416 = _14412 ? _14415 : _14410;
    assign _14417 = _14416[62:0];
    assign _14419 = { _14417,
                      _14418 };
    assign _14420 = _14419 < _14023;
    assign _14421 = ~ _14420;
    assign _14409 = _14020[20:20];
    assign _14406 = _14401 - _14023;
    assign _14407 = _14403 ? _14406 : _14401;
    assign _14408 = _14407[62:0];
    assign _14410 = { _14408,
                      _14409 };
    assign _14411 = _14410 < _14023;
    assign _14412 = ~ _14411;
    assign _14400 = _14020[21:21];
    assign _14397 = _14392 - _14023;
    assign _14398 = _14394 ? _14397 : _14392;
    assign _14399 = _14398[62:0];
    assign _14401 = { _14399,
                      _14400 };
    assign _14402 = _14401 < _14023;
    assign _14403 = ~ _14402;
    assign _14391 = _14020[22:22];
    assign _14388 = _14383 - _14023;
    assign _14389 = _14385 ? _14388 : _14383;
    assign _14390 = _14389[62:0];
    assign _14392 = { _14390,
                      _14391 };
    assign _14393 = _14392 < _14023;
    assign _14394 = ~ _14393;
    assign _14382 = _14020[23:23];
    assign _14379 = _14374 - _14023;
    assign _14380 = _14376 ? _14379 : _14374;
    assign _14381 = _14380[62:0];
    assign _14383 = { _14381,
                      _14382 };
    assign _14384 = _14383 < _14023;
    assign _14385 = ~ _14384;
    assign _14373 = _14020[24:24];
    assign _14370 = _14365 - _14023;
    assign _14371 = _14367 ? _14370 : _14365;
    assign _14372 = _14371[62:0];
    assign _14374 = { _14372,
                      _14373 };
    assign _14375 = _14374 < _14023;
    assign _14376 = ~ _14375;
    assign _14364 = _14020[25:25];
    assign _14361 = _14356 - _14023;
    assign _14362 = _14358 ? _14361 : _14356;
    assign _14363 = _14362[62:0];
    assign _14365 = { _14363,
                      _14364 };
    assign _14366 = _14365 < _14023;
    assign _14367 = ~ _14366;
    assign _14355 = _14020[26:26];
    assign _14352 = _14347 - _14023;
    assign _14353 = _14349 ? _14352 : _14347;
    assign _14354 = _14353[62:0];
    assign _14356 = { _14354,
                      _14355 };
    assign _14357 = _14356 < _14023;
    assign _14358 = ~ _14357;
    assign _14346 = _14020[27:27];
    assign _14343 = _14338 - _14023;
    assign _14344 = _14340 ? _14343 : _14338;
    assign _14345 = _14344[62:0];
    assign _14347 = { _14345,
                      _14346 };
    assign _14348 = _14347 < _14023;
    assign _14349 = ~ _14348;
    assign _14337 = _14020[28:28];
    assign _14334 = _14329 - _14023;
    assign _14335 = _14331 ? _14334 : _14329;
    assign _14336 = _14335[62:0];
    assign _14338 = { _14336,
                      _14337 };
    assign _14339 = _14338 < _14023;
    assign _14340 = ~ _14339;
    assign _14328 = _14020[29:29];
    assign _14325 = _14320 - _14023;
    assign _14326 = _14322 ? _14325 : _14320;
    assign _14327 = _14326[62:0];
    assign _14329 = { _14327,
                      _14328 };
    assign _14330 = _14329 < _14023;
    assign _14331 = ~ _14330;
    assign _14319 = _14020[30:30];
    assign _14316 = _14311 - _14023;
    assign _14317 = _14313 ? _14316 : _14311;
    assign _14318 = _14317[62:0];
    assign _14320 = { _14318,
                      _14319 };
    assign _14321 = _14320 < _14023;
    assign _14322 = ~ _14321;
    assign _14310 = _14020[31:31];
    assign _14307 = _14302 - _14023;
    assign _14308 = _14304 ? _14307 : _14302;
    assign _14309 = _14308[62:0];
    assign _14311 = { _14309,
                      _14310 };
    assign _14312 = _14311 < _14023;
    assign _14313 = ~ _14312;
    assign _14301 = _14020[32:32];
    assign _14298 = _14293 - _14023;
    assign _14299 = _14295 ? _14298 : _14293;
    assign _14300 = _14299[62:0];
    assign _14302 = { _14300,
                      _14301 };
    assign _14303 = _14302 < _14023;
    assign _14304 = ~ _14303;
    assign _14292 = _14020[33:33];
    assign _14289 = _14284 - _14023;
    assign _14290 = _14286 ? _14289 : _14284;
    assign _14291 = _14290[62:0];
    assign _14293 = { _14291,
                      _14292 };
    assign _14294 = _14293 < _14023;
    assign _14295 = ~ _14294;
    assign _14283 = _14020[34:34];
    assign _14280 = _14275 - _14023;
    assign _14281 = _14277 ? _14280 : _14275;
    assign _14282 = _14281[62:0];
    assign _14284 = { _14282,
                      _14283 };
    assign _14285 = _14284 < _14023;
    assign _14286 = ~ _14285;
    assign _14274 = _14020[35:35];
    assign _14271 = _14266 - _14023;
    assign _14272 = _14268 ? _14271 : _14266;
    assign _14273 = _14272[62:0];
    assign _14275 = { _14273,
                      _14274 };
    assign _14276 = _14275 < _14023;
    assign _14277 = ~ _14276;
    assign _14265 = _14020[36:36];
    assign _14262 = _14257 - _14023;
    assign _14263 = _14259 ? _14262 : _14257;
    assign _14264 = _14263[62:0];
    assign _14266 = { _14264,
                      _14265 };
    assign _14267 = _14266 < _14023;
    assign _14268 = ~ _14267;
    assign _14256 = _14020[37:37];
    assign _14253 = _14248 - _14023;
    assign _14254 = _14250 ? _14253 : _14248;
    assign _14255 = _14254[62:0];
    assign _14257 = { _14255,
                      _14256 };
    assign _14258 = _14257 < _14023;
    assign _14259 = ~ _14258;
    assign _14247 = _14020[38:38];
    assign _14244 = _14239 - _14023;
    assign _14245 = _14241 ? _14244 : _14239;
    assign _14246 = _14245[62:0];
    assign _14248 = { _14246,
                      _14247 };
    assign _14249 = _14248 < _14023;
    assign _14250 = ~ _14249;
    assign _14238 = _14020[39:39];
    assign _14235 = _14230 - _14023;
    assign _14236 = _14232 ? _14235 : _14230;
    assign _14237 = _14236[62:0];
    assign _14239 = { _14237,
                      _14238 };
    assign _14240 = _14239 < _14023;
    assign _14241 = ~ _14240;
    assign _14229 = _14020[40:40];
    assign _14226 = _14221 - _14023;
    assign _14227 = _14223 ? _14226 : _14221;
    assign _14228 = _14227[62:0];
    assign _14230 = { _14228,
                      _14229 };
    assign _14231 = _14230 < _14023;
    assign _14232 = ~ _14231;
    assign _14220 = _14020[41:41];
    assign _14217 = _14212 - _14023;
    assign _14218 = _14214 ? _14217 : _14212;
    assign _14219 = _14218[62:0];
    assign _14221 = { _14219,
                      _14220 };
    assign _14222 = _14221 < _14023;
    assign _14223 = ~ _14222;
    assign _14211 = _14020[42:42];
    assign _14208 = _14203 - _14023;
    assign _14209 = _14205 ? _14208 : _14203;
    assign _14210 = _14209[62:0];
    assign _14212 = { _14210,
                      _14211 };
    assign _14213 = _14212 < _14023;
    assign _14214 = ~ _14213;
    assign _14202 = _14020[43:43];
    assign _14199 = _14194 - _14023;
    assign _14200 = _14196 ? _14199 : _14194;
    assign _14201 = _14200[62:0];
    assign _14203 = { _14201,
                      _14202 };
    assign _14204 = _14203 < _14023;
    assign _14205 = ~ _14204;
    assign _14193 = _14020[44:44];
    assign _14190 = _14185 - _14023;
    assign _14191 = _14187 ? _14190 : _14185;
    assign _14192 = _14191[62:0];
    assign _14194 = { _14192,
                      _14193 };
    assign _14195 = _14194 < _14023;
    assign _14196 = ~ _14195;
    assign _14184 = _14020[45:45];
    assign _14181 = _14176 - _14023;
    assign _14182 = _14178 ? _14181 : _14176;
    assign _14183 = _14182[62:0];
    assign _14185 = { _14183,
                      _14184 };
    assign _14186 = _14185 < _14023;
    assign _14187 = ~ _14186;
    assign _14175 = _14020[46:46];
    assign _14172 = _14167 - _14023;
    assign _14173 = _14169 ? _14172 : _14167;
    assign _14174 = _14173[62:0];
    assign _14176 = { _14174,
                      _14175 };
    assign _14177 = _14176 < _14023;
    assign _14178 = ~ _14177;
    assign _14166 = _14020[47:47];
    assign _14163 = _14158 - _14023;
    assign _14164 = _14160 ? _14163 : _14158;
    assign _14165 = _14164[62:0];
    assign _14167 = { _14165,
                      _14166 };
    assign _14168 = _14167 < _14023;
    assign _14169 = ~ _14168;
    assign _14157 = _14020[48:48];
    assign _14154 = _14149 - _14023;
    assign _14155 = _14151 ? _14154 : _14149;
    assign _14156 = _14155[62:0];
    assign _14158 = { _14156,
                      _14157 };
    assign _14159 = _14158 < _14023;
    assign _14160 = ~ _14159;
    assign _14148 = _14020[49:49];
    assign _14145 = _14140 - _14023;
    assign _14146 = _14142 ? _14145 : _14140;
    assign _14147 = _14146[62:0];
    assign _14149 = { _14147,
                      _14148 };
    assign _14150 = _14149 < _14023;
    assign _14151 = ~ _14150;
    assign _14139 = _14020[50:50];
    assign _14136 = _14131 - _14023;
    assign _14137 = _14133 ? _14136 : _14131;
    assign _14138 = _14137[62:0];
    assign _14140 = { _14138,
                      _14139 };
    assign _14141 = _14140 < _14023;
    assign _14142 = ~ _14141;
    assign _14130 = _14020[51:51];
    assign _14127 = _14122 - _14023;
    assign _14128 = _14124 ? _14127 : _14122;
    assign _14129 = _14128[62:0];
    assign _14131 = { _14129,
                      _14130 };
    assign _14132 = _14131 < _14023;
    assign _14133 = ~ _14132;
    assign _14121 = _14020[52:52];
    assign _14118 = _14113 - _14023;
    assign _14119 = _14115 ? _14118 : _14113;
    assign _14120 = _14119[62:0];
    assign _14122 = { _14120,
                      _14121 };
    assign _14123 = _14122 < _14023;
    assign _14124 = ~ _14123;
    assign _14112 = _14020[53:53];
    assign _14109 = _14104 - _14023;
    assign _14110 = _14106 ? _14109 : _14104;
    assign _14111 = _14110[62:0];
    assign _14113 = { _14111,
                      _14112 };
    assign _14114 = _14113 < _14023;
    assign _14115 = ~ _14114;
    assign _14103 = _14020[54:54];
    assign _14100 = _14095 - _14023;
    assign _14101 = _14097 ? _14100 : _14095;
    assign _14102 = _14101[62:0];
    assign _14104 = { _14102,
                      _14103 };
    assign _14105 = _14104 < _14023;
    assign _14106 = ~ _14105;
    assign _14094 = _14020[55:55];
    assign _14091 = _14086 - _14023;
    assign _14092 = _14088 ? _14091 : _14086;
    assign _14093 = _14092[62:0];
    assign _14095 = { _14093,
                      _14094 };
    assign _14096 = _14095 < _14023;
    assign _14097 = ~ _14096;
    assign _14085 = _14020[56:56];
    assign _14082 = _14077 - _14023;
    assign _14083 = _14079 ? _14082 : _14077;
    assign _14084 = _14083[62:0];
    assign _14086 = { _14084,
                      _14085 };
    assign _14087 = _14086 < _14023;
    assign _14088 = ~ _14087;
    assign _14076 = _14020[57:57];
    assign _14073 = _14068 - _14023;
    assign _14074 = _14070 ? _14073 : _14068;
    assign _14075 = _14074[62:0];
    assign _14077 = { _14075,
                      _14076 };
    assign _14078 = _14077 < _14023;
    assign _14079 = ~ _14078;
    assign _14067 = _14020[58:58];
    assign _14064 = _14059 - _14023;
    assign _14065 = _14061 ? _14064 : _14059;
    assign _14066 = _14065[62:0];
    assign _14068 = { _14066,
                      _14067 };
    assign _14069 = _14068 < _14023;
    assign _14070 = ~ _14069;
    assign _14058 = _14020[59:59];
    assign _14055 = _14050 - _14023;
    assign _14056 = _14052 ? _14055 : _14050;
    assign _14057 = _14056[62:0];
    assign _14059 = { _14057,
                      _14058 };
    assign _14060 = _14059 < _14023;
    assign _14061 = ~ _14060;
    assign _14049 = _14020[60:60];
    assign _14046 = _14041 - _14023;
    assign _14047 = _14043 ? _14046 : _14041;
    assign _14048 = _14047[62:0];
    assign _14050 = { _14048,
                      _14049 };
    assign _14051 = _14050 < _14023;
    assign _14052 = ~ _14051;
    assign _14040 = _14020[61:61];
    assign _14037 = _14032 - _14023;
    assign _14038 = _14034 ? _14037 : _14032;
    assign _14039 = _14038[62:0];
    assign _14041 = { _14039,
                      _14040 };
    assign _14042 = _14041 < _14023;
    assign _14043 = ~ _14042;
    assign _14031 = _14020[62:62];
    assign _14028 = _14022 - _14023;
    assign _14029 = _14025 ? _14028 : _14022;
    assign _14030 = _14029[62:0];
    assign _14032 = { _14030,
                      _14031 };
    assign _14033 = _14032 < _14023;
    assign _14034 = ~ _14033;
    assign _14023 = 64'b0000000000000000000000000000000000000000000100001111010001000111;
    assign _14019 = 64'b0000000000000000000000000000000000000000000100001111010001000110;
    assign _14020 = _3 + _14019;
    assign _14021 = _14020[63:63];
    assign _14022 = { _22185,
                      _14021 };
    assign _14024 = _14022 < _14023;
    assign _14025 = ~ _14024;
    assign _14026 = { _22185,
                      _14025 };
    assign _14027 = _14026[62:0];
    assign _14035 = { _14027,
                      _14034 };
    assign _14036 = _14035[62:0];
    assign _14044 = { _14036,
                      _14043 };
    assign _14045 = _14044[62:0];
    assign _14053 = { _14045,
                      _14052 };
    assign _14054 = _14053[62:0];
    assign _14062 = { _14054,
                      _14061 };
    assign _14063 = _14062[62:0];
    assign _14071 = { _14063,
                      _14070 };
    assign _14072 = _14071[62:0];
    assign _14080 = { _14072,
                      _14079 };
    assign _14081 = _14080[62:0];
    assign _14089 = { _14081,
                      _14088 };
    assign _14090 = _14089[62:0];
    assign _14098 = { _14090,
                      _14097 };
    assign _14099 = _14098[62:0];
    assign _14107 = { _14099,
                      _14106 };
    assign _14108 = _14107[62:0];
    assign _14116 = { _14108,
                      _14115 };
    assign _14117 = _14116[62:0];
    assign _14125 = { _14117,
                      _14124 };
    assign _14126 = _14125[62:0];
    assign _14134 = { _14126,
                      _14133 };
    assign _14135 = _14134[62:0];
    assign _14143 = { _14135,
                      _14142 };
    assign _14144 = _14143[62:0];
    assign _14152 = { _14144,
                      _14151 };
    assign _14153 = _14152[62:0];
    assign _14161 = { _14153,
                      _14160 };
    assign _14162 = _14161[62:0];
    assign _14170 = { _14162,
                      _14169 };
    assign _14171 = _14170[62:0];
    assign _14179 = { _14171,
                      _14178 };
    assign _14180 = _14179[62:0];
    assign _14188 = { _14180,
                      _14187 };
    assign _14189 = _14188[62:0];
    assign _14197 = { _14189,
                      _14196 };
    assign _14198 = _14197[62:0];
    assign _14206 = { _14198,
                      _14205 };
    assign _14207 = _14206[62:0];
    assign _14215 = { _14207,
                      _14214 };
    assign _14216 = _14215[62:0];
    assign _14224 = { _14216,
                      _14223 };
    assign _14225 = _14224[62:0];
    assign _14233 = { _14225,
                      _14232 };
    assign _14234 = _14233[62:0];
    assign _14242 = { _14234,
                      _14241 };
    assign _14243 = _14242[62:0];
    assign _14251 = { _14243,
                      _14250 };
    assign _14252 = _14251[62:0];
    assign _14260 = { _14252,
                      _14259 };
    assign _14261 = _14260[62:0];
    assign _14269 = { _14261,
                      _14268 };
    assign _14270 = _14269[62:0];
    assign _14278 = { _14270,
                      _14277 };
    assign _14279 = _14278[62:0];
    assign _14287 = { _14279,
                      _14286 };
    assign _14288 = _14287[62:0];
    assign _14296 = { _14288,
                      _14295 };
    assign _14297 = _14296[62:0];
    assign _14305 = { _14297,
                      _14304 };
    assign _14306 = _14305[62:0];
    assign _14314 = { _14306,
                      _14313 };
    assign _14315 = _14314[62:0];
    assign _14323 = { _14315,
                      _14322 };
    assign _14324 = _14323[62:0];
    assign _14332 = { _14324,
                      _14331 };
    assign _14333 = _14332[62:0];
    assign _14341 = { _14333,
                      _14340 };
    assign _14342 = _14341[62:0];
    assign _14350 = { _14342,
                      _14349 };
    assign _14351 = _14350[62:0];
    assign _14359 = { _14351,
                      _14358 };
    assign _14360 = _14359[62:0];
    assign _14368 = { _14360,
                      _14367 };
    assign _14369 = _14368[62:0];
    assign _14377 = { _14369,
                      _14376 };
    assign _14378 = _14377[62:0];
    assign _14386 = { _14378,
                      _14385 };
    assign _14387 = _14386[62:0];
    assign _14395 = { _14387,
                      _14394 };
    assign _14396 = _14395[62:0];
    assign _14404 = { _14396,
                      _14403 };
    assign _14405 = _14404[62:0];
    assign _14413 = { _14405,
                      _14412 };
    assign _14414 = _14413[62:0];
    assign _14422 = { _14414,
                      _14421 };
    assign _14423 = _14422[62:0];
    assign _14431 = { _14423,
                      _14430 };
    assign _14432 = _14431[62:0];
    assign _14440 = { _14432,
                      _14439 };
    assign _14441 = _14440[62:0];
    assign _14449 = { _14441,
                      _14448 };
    assign _14450 = _14449[62:0];
    assign _14458 = { _14450,
                      _14457 };
    assign _14459 = _14458[62:0];
    assign _14467 = { _14459,
                      _14466 };
    assign _14468 = _14467[62:0];
    assign _14476 = { _14468,
                      _14475 };
    assign _14477 = _14476[62:0];
    assign _14485 = { _14477,
                      _14484 };
    assign _14486 = _14485[62:0];
    assign _14494 = { _14486,
                      _14493 };
    assign _14495 = _14494[62:0];
    assign _14503 = { _14495,
                      _14502 };
    assign _14504 = _14503[62:0];
    assign _14512 = { _14504,
                      _14511 };
    assign _14513 = _14512[62:0];
    assign _14521 = { _14513,
                      _14520 };
    assign _14522 = _14521[62:0];
    assign _14530 = { _14522,
                      _14529 };
    assign _14531 = _14530[62:0];
    assign _14539 = { _14531,
                      _14538 };
    assign _14540 = _14539[62:0];
    assign _14548 = { _14540,
                      _14547 };
    assign _14549 = _14548[62:0];
    assign _14557 = { _14549,
                      _14556 };
    assign _14558 = _14557[62:0];
    assign _14566 = { _14558,
                      _14565 };
    assign _14567 = _14566[62:0];
    assign _14575 = { _14567,
                      _14574 };
    assign _14576 = _14575[62:0];
    assign _14584 = { _14576,
                      _14583 };
    assign _14585 = _14584[62:0];
    assign _14593 = { _14585,
                      _14592 };
    assign _14594 = _14593 * _14023;
    assign _14595 = _14594[63:0];
    assign _14596 = _14023 < _14595;
    assign _14597 = _14596 ? _14595 : _14023;
    assign _14013 = 64'b0000000000000000000000000000000000000000100110001001011001111111;
    assign _14014 = _5 < _14013;
    assign _14015 = _14014 ? _5 : _14013;
    assign _14598 = _14015 < _14597;
    assign _14599 = ~ _14598;
    assign _15762 = _14599 ? _15761 : _21604;
    assign _14003 = _13434[0:0];
    assign _14000 = _13995 - _22192;
    assign _14001 = _13997 ? _14000 : _13995;
    assign _14002 = _14001[62:0];
    assign _14004 = { _14002,
                      _14003 };
    assign _14005 = _14004 < _22192;
    assign _14006 = ~ _14005;
    assign _13994 = _13434[1:1];
    assign _13991 = _13986 - _22192;
    assign _13992 = _13988 ? _13991 : _13986;
    assign _13993 = _13992[62:0];
    assign _13995 = { _13993,
                      _13994 };
    assign _13996 = _13995 < _22192;
    assign _13997 = ~ _13996;
    assign _13985 = _13434[2:2];
    assign _13982 = _13977 - _22192;
    assign _13983 = _13979 ? _13982 : _13977;
    assign _13984 = _13983[62:0];
    assign _13986 = { _13984,
                      _13985 };
    assign _13987 = _13986 < _22192;
    assign _13988 = ~ _13987;
    assign _13976 = _13434[3:3];
    assign _13973 = _13968 - _22192;
    assign _13974 = _13970 ? _13973 : _13968;
    assign _13975 = _13974[62:0];
    assign _13977 = { _13975,
                      _13976 };
    assign _13978 = _13977 < _22192;
    assign _13979 = ~ _13978;
    assign _13967 = _13434[4:4];
    assign _13964 = _13959 - _22192;
    assign _13965 = _13961 ? _13964 : _13959;
    assign _13966 = _13965[62:0];
    assign _13968 = { _13966,
                      _13967 };
    assign _13969 = _13968 < _22192;
    assign _13970 = ~ _13969;
    assign _13958 = _13434[5:5];
    assign _13955 = _13950 - _22192;
    assign _13956 = _13952 ? _13955 : _13950;
    assign _13957 = _13956[62:0];
    assign _13959 = { _13957,
                      _13958 };
    assign _13960 = _13959 < _22192;
    assign _13961 = ~ _13960;
    assign _13949 = _13434[6:6];
    assign _13946 = _13941 - _22192;
    assign _13947 = _13943 ? _13946 : _13941;
    assign _13948 = _13947[62:0];
    assign _13950 = { _13948,
                      _13949 };
    assign _13951 = _13950 < _22192;
    assign _13952 = ~ _13951;
    assign _13940 = _13434[7:7];
    assign _13937 = _13932 - _22192;
    assign _13938 = _13934 ? _13937 : _13932;
    assign _13939 = _13938[62:0];
    assign _13941 = { _13939,
                      _13940 };
    assign _13942 = _13941 < _22192;
    assign _13943 = ~ _13942;
    assign _13931 = _13434[8:8];
    assign _13928 = _13923 - _22192;
    assign _13929 = _13925 ? _13928 : _13923;
    assign _13930 = _13929[62:0];
    assign _13932 = { _13930,
                      _13931 };
    assign _13933 = _13932 < _22192;
    assign _13934 = ~ _13933;
    assign _13922 = _13434[9:9];
    assign _13919 = _13914 - _22192;
    assign _13920 = _13916 ? _13919 : _13914;
    assign _13921 = _13920[62:0];
    assign _13923 = { _13921,
                      _13922 };
    assign _13924 = _13923 < _22192;
    assign _13925 = ~ _13924;
    assign _13913 = _13434[10:10];
    assign _13910 = _13905 - _22192;
    assign _13911 = _13907 ? _13910 : _13905;
    assign _13912 = _13911[62:0];
    assign _13914 = { _13912,
                      _13913 };
    assign _13915 = _13914 < _22192;
    assign _13916 = ~ _13915;
    assign _13904 = _13434[11:11];
    assign _13901 = _13896 - _22192;
    assign _13902 = _13898 ? _13901 : _13896;
    assign _13903 = _13902[62:0];
    assign _13905 = { _13903,
                      _13904 };
    assign _13906 = _13905 < _22192;
    assign _13907 = ~ _13906;
    assign _13895 = _13434[12:12];
    assign _13892 = _13887 - _22192;
    assign _13893 = _13889 ? _13892 : _13887;
    assign _13894 = _13893[62:0];
    assign _13896 = { _13894,
                      _13895 };
    assign _13897 = _13896 < _22192;
    assign _13898 = ~ _13897;
    assign _13886 = _13434[13:13];
    assign _13883 = _13878 - _22192;
    assign _13884 = _13880 ? _13883 : _13878;
    assign _13885 = _13884[62:0];
    assign _13887 = { _13885,
                      _13886 };
    assign _13888 = _13887 < _22192;
    assign _13889 = ~ _13888;
    assign _13877 = _13434[14:14];
    assign _13874 = _13869 - _22192;
    assign _13875 = _13871 ? _13874 : _13869;
    assign _13876 = _13875[62:0];
    assign _13878 = { _13876,
                      _13877 };
    assign _13879 = _13878 < _22192;
    assign _13880 = ~ _13879;
    assign _13868 = _13434[15:15];
    assign _13865 = _13860 - _22192;
    assign _13866 = _13862 ? _13865 : _13860;
    assign _13867 = _13866[62:0];
    assign _13869 = { _13867,
                      _13868 };
    assign _13870 = _13869 < _22192;
    assign _13871 = ~ _13870;
    assign _13859 = _13434[16:16];
    assign _13856 = _13851 - _22192;
    assign _13857 = _13853 ? _13856 : _13851;
    assign _13858 = _13857[62:0];
    assign _13860 = { _13858,
                      _13859 };
    assign _13861 = _13860 < _22192;
    assign _13862 = ~ _13861;
    assign _13850 = _13434[17:17];
    assign _13847 = _13842 - _22192;
    assign _13848 = _13844 ? _13847 : _13842;
    assign _13849 = _13848[62:0];
    assign _13851 = { _13849,
                      _13850 };
    assign _13852 = _13851 < _22192;
    assign _13853 = ~ _13852;
    assign _13841 = _13434[18:18];
    assign _13838 = _13833 - _22192;
    assign _13839 = _13835 ? _13838 : _13833;
    assign _13840 = _13839[62:0];
    assign _13842 = { _13840,
                      _13841 };
    assign _13843 = _13842 < _22192;
    assign _13844 = ~ _13843;
    assign _13832 = _13434[19:19];
    assign _13829 = _13824 - _22192;
    assign _13830 = _13826 ? _13829 : _13824;
    assign _13831 = _13830[62:0];
    assign _13833 = { _13831,
                      _13832 };
    assign _13834 = _13833 < _22192;
    assign _13835 = ~ _13834;
    assign _13823 = _13434[20:20];
    assign _13820 = _13815 - _22192;
    assign _13821 = _13817 ? _13820 : _13815;
    assign _13822 = _13821[62:0];
    assign _13824 = { _13822,
                      _13823 };
    assign _13825 = _13824 < _22192;
    assign _13826 = ~ _13825;
    assign _13814 = _13434[21:21];
    assign _13811 = _13806 - _22192;
    assign _13812 = _13808 ? _13811 : _13806;
    assign _13813 = _13812[62:0];
    assign _13815 = { _13813,
                      _13814 };
    assign _13816 = _13815 < _22192;
    assign _13817 = ~ _13816;
    assign _13805 = _13434[22:22];
    assign _13802 = _13797 - _22192;
    assign _13803 = _13799 ? _13802 : _13797;
    assign _13804 = _13803[62:0];
    assign _13806 = { _13804,
                      _13805 };
    assign _13807 = _13806 < _22192;
    assign _13808 = ~ _13807;
    assign _13796 = _13434[23:23];
    assign _13793 = _13788 - _22192;
    assign _13794 = _13790 ? _13793 : _13788;
    assign _13795 = _13794[62:0];
    assign _13797 = { _13795,
                      _13796 };
    assign _13798 = _13797 < _22192;
    assign _13799 = ~ _13798;
    assign _13787 = _13434[24:24];
    assign _13784 = _13779 - _22192;
    assign _13785 = _13781 ? _13784 : _13779;
    assign _13786 = _13785[62:0];
    assign _13788 = { _13786,
                      _13787 };
    assign _13789 = _13788 < _22192;
    assign _13790 = ~ _13789;
    assign _13778 = _13434[25:25];
    assign _13775 = _13770 - _22192;
    assign _13776 = _13772 ? _13775 : _13770;
    assign _13777 = _13776[62:0];
    assign _13779 = { _13777,
                      _13778 };
    assign _13780 = _13779 < _22192;
    assign _13781 = ~ _13780;
    assign _13769 = _13434[26:26];
    assign _13766 = _13761 - _22192;
    assign _13767 = _13763 ? _13766 : _13761;
    assign _13768 = _13767[62:0];
    assign _13770 = { _13768,
                      _13769 };
    assign _13771 = _13770 < _22192;
    assign _13772 = ~ _13771;
    assign _13760 = _13434[27:27];
    assign _13757 = _13752 - _22192;
    assign _13758 = _13754 ? _13757 : _13752;
    assign _13759 = _13758[62:0];
    assign _13761 = { _13759,
                      _13760 };
    assign _13762 = _13761 < _22192;
    assign _13763 = ~ _13762;
    assign _13751 = _13434[28:28];
    assign _13748 = _13743 - _22192;
    assign _13749 = _13745 ? _13748 : _13743;
    assign _13750 = _13749[62:0];
    assign _13752 = { _13750,
                      _13751 };
    assign _13753 = _13752 < _22192;
    assign _13754 = ~ _13753;
    assign _13742 = _13434[29:29];
    assign _13739 = _13734 - _22192;
    assign _13740 = _13736 ? _13739 : _13734;
    assign _13741 = _13740[62:0];
    assign _13743 = { _13741,
                      _13742 };
    assign _13744 = _13743 < _22192;
    assign _13745 = ~ _13744;
    assign _13733 = _13434[30:30];
    assign _13730 = _13725 - _22192;
    assign _13731 = _13727 ? _13730 : _13725;
    assign _13732 = _13731[62:0];
    assign _13734 = { _13732,
                      _13733 };
    assign _13735 = _13734 < _22192;
    assign _13736 = ~ _13735;
    assign _13724 = _13434[31:31];
    assign _13721 = _13716 - _22192;
    assign _13722 = _13718 ? _13721 : _13716;
    assign _13723 = _13722[62:0];
    assign _13725 = { _13723,
                      _13724 };
    assign _13726 = _13725 < _22192;
    assign _13727 = ~ _13726;
    assign _13715 = _13434[32:32];
    assign _13712 = _13707 - _22192;
    assign _13713 = _13709 ? _13712 : _13707;
    assign _13714 = _13713[62:0];
    assign _13716 = { _13714,
                      _13715 };
    assign _13717 = _13716 < _22192;
    assign _13718 = ~ _13717;
    assign _13706 = _13434[33:33];
    assign _13703 = _13698 - _22192;
    assign _13704 = _13700 ? _13703 : _13698;
    assign _13705 = _13704[62:0];
    assign _13707 = { _13705,
                      _13706 };
    assign _13708 = _13707 < _22192;
    assign _13709 = ~ _13708;
    assign _13697 = _13434[34:34];
    assign _13694 = _13689 - _22192;
    assign _13695 = _13691 ? _13694 : _13689;
    assign _13696 = _13695[62:0];
    assign _13698 = { _13696,
                      _13697 };
    assign _13699 = _13698 < _22192;
    assign _13700 = ~ _13699;
    assign _13688 = _13434[35:35];
    assign _13685 = _13680 - _22192;
    assign _13686 = _13682 ? _13685 : _13680;
    assign _13687 = _13686[62:0];
    assign _13689 = { _13687,
                      _13688 };
    assign _13690 = _13689 < _22192;
    assign _13691 = ~ _13690;
    assign _13679 = _13434[36:36];
    assign _13676 = _13671 - _22192;
    assign _13677 = _13673 ? _13676 : _13671;
    assign _13678 = _13677[62:0];
    assign _13680 = { _13678,
                      _13679 };
    assign _13681 = _13680 < _22192;
    assign _13682 = ~ _13681;
    assign _13670 = _13434[37:37];
    assign _13667 = _13662 - _22192;
    assign _13668 = _13664 ? _13667 : _13662;
    assign _13669 = _13668[62:0];
    assign _13671 = { _13669,
                      _13670 };
    assign _13672 = _13671 < _22192;
    assign _13673 = ~ _13672;
    assign _13661 = _13434[38:38];
    assign _13658 = _13653 - _22192;
    assign _13659 = _13655 ? _13658 : _13653;
    assign _13660 = _13659[62:0];
    assign _13662 = { _13660,
                      _13661 };
    assign _13663 = _13662 < _22192;
    assign _13664 = ~ _13663;
    assign _13652 = _13434[39:39];
    assign _13649 = _13644 - _22192;
    assign _13650 = _13646 ? _13649 : _13644;
    assign _13651 = _13650[62:0];
    assign _13653 = { _13651,
                      _13652 };
    assign _13654 = _13653 < _22192;
    assign _13655 = ~ _13654;
    assign _13643 = _13434[40:40];
    assign _13640 = _13635 - _22192;
    assign _13641 = _13637 ? _13640 : _13635;
    assign _13642 = _13641[62:0];
    assign _13644 = { _13642,
                      _13643 };
    assign _13645 = _13644 < _22192;
    assign _13646 = ~ _13645;
    assign _13634 = _13434[41:41];
    assign _13631 = _13626 - _22192;
    assign _13632 = _13628 ? _13631 : _13626;
    assign _13633 = _13632[62:0];
    assign _13635 = { _13633,
                      _13634 };
    assign _13636 = _13635 < _22192;
    assign _13637 = ~ _13636;
    assign _13625 = _13434[42:42];
    assign _13622 = _13617 - _22192;
    assign _13623 = _13619 ? _13622 : _13617;
    assign _13624 = _13623[62:0];
    assign _13626 = { _13624,
                      _13625 };
    assign _13627 = _13626 < _22192;
    assign _13628 = ~ _13627;
    assign _13616 = _13434[43:43];
    assign _13613 = _13608 - _22192;
    assign _13614 = _13610 ? _13613 : _13608;
    assign _13615 = _13614[62:0];
    assign _13617 = { _13615,
                      _13616 };
    assign _13618 = _13617 < _22192;
    assign _13619 = ~ _13618;
    assign _13607 = _13434[44:44];
    assign _13604 = _13599 - _22192;
    assign _13605 = _13601 ? _13604 : _13599;
    assign _13606 = _13605[62:0];
    assign _13608 = { _13606,
                      _13607 };
    assign _13609 = _13608 < _22192;
    assign _13610 = ~ _13609;
    assign _13598 = _13434[45:45];
    assign _13595 = _13590 - _22192;
    assign _13596 = _13592 ? _13595 : _13590;
    assign _13597 = _13596[62:0];
    assign _13599 = { _13597,
                      _13598 };
    assign _13600 = _13599 < _22192;
    assign _13601 = ~ _13600;
    assign _13589 = _13434[46:46];
    assign _13586 = _13581 - _22192;
    assign _13587 = _13583 ? _13586 : _13581;
    assign _13588 = _13587[62:0];
    assign _13590 = { _13588,
                      _13589 };
    assign _13591 = _13590 < _22192;
    assign _13592 = ~ _13591;
    assign _13580 = _13434[47:47];
    assign _13577 = _13572 - _22192;
    assign _13578 = _13574 ? _13577 : _13572;
    assign _13579 = _13578[62:0];
    assign _13581 = { _13579,
                      _13580 };
    assign _13582 = _13581 < _22192;
    assign _13583 = ~ _13582;
    assign _13571 = _13434[48:48];
    assign _13568 = _13563 - _22192;
    assign _13569 = _13565 ? _13568 : _13563;
    assign _13570 = _13569[62:0];
    assign _13572 = { _13570,
                      _13571 };
    assign _13573 = _13572 < _22192;
    assign _13574 = ~ _13573;
    assign _13562 = _13434[49:49];
    assign _13559 = _13554 - _22192;
    assign _13560 = _13556 ? _13559 : _13554;
    assign _13561 = _13560[62:0];
    assign _13563 = { _13561,
                      _13562 };
    assign _13564 = _13563 < _22192;
    assign _13565 = ~ _13564;
    assign _13553 = _13434[50:50];
    assign _13550 = _13545 - _22192;
    assign _13551 = _13547 ? _13550 : _13545;
    assign _13552 = _13551[62:0];
    assign _13554 = { _13552,
                      _13553 };
    assign _13555 = _13554 < _22192;
    assign _13556 = ~ _13555;
    assign _13544 = _13434[51:51];
    assign _13541 = _13536 - _22192;
    assign _13542 = _13538 ? _13541 : _13536;
    assign _13543 = _13542[62:0];
    assign _13545 = { _13543,
                      _13544 };
    assign _13546 = _13545 < _22192;
    assign _13547 = ~ _13546;
    assign _13535 = _13434[52:52];
    assign _13532 = _13527 - _22192;
    assign _13533 = _13529 ? _13532 : _13527;
    assign _13534 = _13533[62:0];
    assign _13536 = { _13534,
                      _13535 };
    assign _13537 = _13536 < _22192;
    assign _13538 = ~ _13537;
    assign _13526 = _13434[53:53];
    assign _13523 = _13518 - _22192;
    assign _13524 = _13520 ? _13523 : _13518;
    assign _13525 = _13524[62:0];
    assign _13527 = { _13525,
                      _13526 };
    assign _13528 = _13527 < _22192;
    assign _13529 = ~ _13528;
    assign _13517 = _13434[54:54];
    assign _13514 = _13509 - _22192;
    assign _13515 = _13511 ? _13514 : _13509;
    assign _13516 = _13515[62:0];
    assign _13518 = { _13516,
                      _13517 };
    assign _13519 = _13518 < _22192;
    assign _13520 = ~ _13519;
    assign _13508 = _13434[55:55];
    assign _13505 = _13500 - _22192;
    assign _13506 = _13502 ? _13505 : _13500;
    assign _13507 = _13506[62:0];
    assign _13509 = { _13507,
                      _13508 };
    assign _13510 = _13509 < _22192;
    assign _13511 = ~ _13510;
    assign _13499 = _13434[56:56];
    assign _13496 = _13491 - _22192;
    assign _13497 = _13493 ? _13496 : _13491;
    assign _13498 = _13497[62:0];
    assign _13500 = { _13498,
                      _13499 };
    assign _13501 = _13500 < _22192;
    assign _13502 = ~ _13501;
    assign _13490 = _13434[57:57];
    assign _13487 = _13482 - _22192;
    assign _13488 = _13484 ? _13487 : _13482;
    assign _13489 = _13488[62:0];
    assign _13491 = { _13489,
                      _13490 };
    assign _13492 = _13491 < _22192;
    assign _13493 = ~ _13492;
    assign _13481 = _13434[58:58];
    assign _13478 = _13473 - _22192;
    assign _13479 = _13475 ? _13478 : _13473;
    assign _13480 = _13479[62:0];
    assign _13482 = { _13480,
                      _13481 };
    assign _13483 = _13482 < _22192;
    assign _13484 = ~ _13483;
    assign _13472 = _13434[59:59];
    assign _13469 = _13464 - _22192;
    assign _13470 = _13466 ? _13469 : _13464;
    assign _13471 = _13470[62:0];
    assign _13473 = { _13471,
                      _13472 };
    assign _13474 = _13473 < _22192;
    assign _13475 = ~ _13474;
    assign _13463 = _13434[60:60];
    assign _13460 = _13455 - _22192;
    assign _13461 = _13457 ? _13460 : _13455;
    assign _13462 = _13461[62:0];
    assign _13464 = { _13462,
                      _13463 };
    assign _13465 = _13464 < _22192;
    assign _13466 = ~ _13465;
    assign _13454 = _13434[61:61];
    assign _13451 = _13446 - _22192;
    assign _13452 = _13448 ? _13451 : _13446;
    assign _13453 = _13452[62:0];
    assign _13455 = { _13453,
                      _13454 };
    assign _13456 = _13455 < _22192;
    assign _13457 = ~ _13456;
    assign _13445 = _13434[62:62];
    assign _13442 = _13436 - _22192;
    assign _13443 = _13439 ? _13442 : _13436;
    assign _13444 = _13443[62:0];
    assign _13446 = { _13444,
                      _13445 };
    assign _13447 = _13446 < _22192;
    assign _13448 = ~ _13447;
    assign _13432 = _13424 + _22186;
    assign _13433 = _13424 * _13432;
    assign _13434 = _13433[63:0];
    assign _13435 = _13434[63:63];
    assign _13436 = { _22185,
                      _13435 };
    assign _13438 = _13436 < _22192;
    assign _13439 = ~ _13438;
    assign _13440 = { _22185,
                      _13439 };
    assign _13441 = _13440[62:0];
    assign _13449 = { _13441,
                      _13448 };
    assign _13450 = _13449[62:0];
    assign _13458 = { _13450,
                      _13457 };
    assign _13459 = _13458[62:0];
    assign _13467 = { _13459,
                      _13466 };
    assign _13468 = _13467[62:0];
    assign _13476 = { _13468,
                      _13475 };
    assign _13477 = _13476[62:0];
    assign _13485 = { _13477,
                      _13484 };
    assign _13486 = _13485[62:0];
    assign _13494 = { _13486,
                      _13493 };
    assign _13495 = _13494[62:0];
    assign _13503 = { _13495,
                      _13502 };
    assign _13504 = _13503[62:0];
    assign _13512 = { _13504,
                      _13511 };
    assign _13513 = _13512[62:0];
    assign _13521 = { _13513,
                      _13520 };
    assign _13522 = _13521[62:0];
    assign _13530 = { _13522,
                      _13529 };
    assign _13531 = _13530[62:0];
    assign _13539 = { _13531,
                      _13538 };
    assign _13540 = _13539[62:0];
    assign _13548 = { _13540,
                      _13547 };
    assign _13549 = _13548[62:0];
    assign _13557 = { _13549,
                      _13556 };
    assign _13558 = _13557[62:0];
    assign _13566 = { _13558,
                      _13565 };
    assign _13567 = _13566[62:0];
    assign _13575 = { _13567,
                      _13574 };
    assign _13576 = _13575[62:0];
    assign _13584 = { _13576,
                      _13583 };
    assign _13585 = _13584[62:0];
    assign _13593 = { _13585,
                      _13592 };
    assign _13594 = _13593[62:0];
    assign _13602 = { _13594,
                      _13601 };
    assign _13603 = _13602[62:0];
    assign _13611 = { _13603,
                      _13610 };
    assign _13612 = _13611[62:0];
    assign _13620 = { _13612,
                      _13619 };
    assign _13621 = _13620[62:0];
    assign _13629 = { _13621,
                      _13628 };
    assign _13630 = _13629[62:0];
    assign _13638 = { _13630,
                      _13637 };
    assign _13639 = _13638[62:0];
    assign _13647 = { _13639,
                      _13646 };
    assign _13648 = _13647[62:0];
    assign _13656 = { _13648,
                      _13655 };
    assign _13657 = _13656[62:0];
    assign _13665 = { _13657,
                      _13664 };
    assign _13666 = _13665[62:0];
    assign _13674 = { _13666,
                      _13673 };
    assign _13675 = _13674[62:0];
    assign _13683 = { _13675,
                      _13682 };
    assign _13684 = _13683[62:0];
    assign _13692 = { _13684,
                      _13691 };
    assign _13693 = _13692[62:0];
    assign _13701 = { _13693,
                      _13700 };
    assign _13702 = _13701[62:0];
    assign _13710 = { _13702,
                      _13709 };
    assign _13711 = _13710[62:0];
    assign _13719 = { _13711,
                      _13718 };
    assign _13720 = _13719[62:0];
    assign _13728 = { _13720,
                      _13727 };
    assign _13729 = _13728[62:0];
    assign _13737 = { _13729,
                      _13736 };
    assign _13738 = _13737[62:0];
    assign _13746 = { _13738,
                      _13745 };
    assign _13747 = _13746[62:0];
    assign _13755 = { _13747,
                      _13754 };
    assign _13756 = _13755[62:0];
    assign _13764 = { _13756,
                      _13763 };
    assign _13765 = _13764[62:0];
    assign _13773 = { _13765,
                      _13772 };
    assign _13774 = _13773[62:0];
    assign _13782 = { _13774,
                      _13781 };
    assign _13783 = _13782[62:0];
    assign _13791 = { _13783,
                      _13790 };
    assign _13792 = _13791[62:0];
    assign _13800 = { _13792,
                      _13799 };
    assign _13801 = _13800[62:0];
    assign _13809 = { _13801,
                      _13808 };
    assign _13810 = _13809[62:0];
    assign _13818 = { _13810,
                      _13817 };
    assign _13819 = _13818[62:0];
    assign _13827 = { _13819,
                      _13826 };
    assign _13828 = _13827[62:0];
    assign _13836 = { _13828,
                      _13835 };
    assign _13837 = _13836[62:0];
    assign _13845 = { _13837,
                      _13844 };
    assign _13846 = _13845[62:0];
    assign _13854 = { _13846,
                      _13853 };
    assign _13855 = _13854[62:0];
    assign _13863 = { _13855,
                      _13862 };
    assign _13864 = _13863[62:0];
    assign _13872 = { _13864,
                      _13871 };
    assign _13873 = _13872[62:0];
    assign _13881 = { _13873,
                      _13880 };
    assign _13882 = _13881[62:0];
    assign _13890 = { _13882,
                      _13889 };
    assign _13891 = _13890[62:0];
    assign _13899 = { _13891,
                      _13898 };
    assign _13900 = _13899[62:0];
    assign _13908 = { _13900,
                      _13907 };
    assign _13909 = _13908[62:0];
    assign _13917 = { _13909,
                      _13916 };
    assign _13918 = _13917[62:0];
    assign _13926 = { _13918,
                      _13925 };
    assign _13927 = _13926[62:0];
    assign _13935 = { _13927,
                      _13934 };
    assign _13936 = _13935[62:0];
    assign _13944 = { _13936,
                      _13943 };
    assign _13945 = _13944[62:0];
    assign _13953 = { _13945,
                      _13952 };
    assign _13954 = _13953[62:0];
    assign _13962 = { _13954,
                      _13961 };
    assign _13963 = _13962[62:0];
    assign _13971 = { _13963,
                      _13970 };
    assign _13972 = _13971[62:0];
    assign _13980 = { _13972,
                      _13979 };
    assign _13981 = _13980[62:0];
    assign _13989 = { _13981,
                      _13988 };
    assign _13990 = _13989[62:0];
    assign _13998 = { _13990,
                      _13997 };
    assign _13999 = _13998[62:0];
    assign _14007 = { _13999,
                      _14006 };
    assign _14008 = _12272 * _14007;
    assign _14009 = _14008[63:0];
    assign _13420 = _12852[0:0];
    assign _13417 = _13412 - _12272;
    assign _13418 = _13414 ? _13417 : _13412;
    assign _13419 = _13418[62:0];
    assign _13421 = { _13419,
                      _13420 };
    assign _13422 = _13421 < _12272;
    assign _13423 = ~ _13422;
    assign _13411 = _12852[1:1];
    assign _13408 = _13403 - _12272;
    assign _13409 = _13405 ? _13408 : _13403;
    assign _13410 = _13409[62:0];
    assign _13412 = { _13410,
                      _13411 };
    assign _13413 = _13412 < _12272;
    assign _13414 = ~ _13413;
    assign _13402 = _12852[2:2];
    assign _13399 = _13394 - _12272;
    assign _13400 = _13396 ? _13399 : _13394;
    assign _13401 = _13400[62:0];
    assign _13403 = { _13401,
                      _13402 };
    assign _13404 = _13403 < _12272;
    assign _13405 = ~ _13404;
    assign _13393 = _12852[3:3];
    assign _13390 = _13385 - _12272;
    assign _13391 = _13387 ? _13390 : _13385;
    assign _13392 = _13391[62:0];
    assign _13394 = { _13392,
                      _13393 };
    assign _13395 = _13394 < _12272;
    assign _13396 = ~ _13395;
    assign _13384 = _12852[4:4];
    assign _13381 = _13376 - _12272;
    assign _13382 = _13378 ? _13381 : _13376;
    assign _13383 = _13382[62:0];
    assign _13385 = { _13383,
                      _13384 };
    assign _13386 = _13385 < _12272;
    assign _13387 = ~ _13386;
    assign _13375 = _12852[5:5];
    assign _13372 = _13367 - _12272;
    assign _13373 = _13369 ? _13372 : _13367;
    assign _13374 = _13373[62:0];
    assign _13376 = { _13374,
                      _13375 };
    assign _13377 = _13376 < _12272;
    assign _13378 = ~ _13377;
    assign _13366 = _12852[6:6];
    assign _13363 = _13358 - _12272;
    assign _13364 = _13360 ? _13363 : _13358;
    assign _13365 = _13364[62:0];
    assign _13367 = { _13365,
                      _13366 };
    assign _13368 = _13367 < _12272;
    assign _13369 = ~ _13368;
    assign _13357 = _12852[7:7];
    assign _13354 = _13349 - _12272;
    assign _13355 = _13351 ? _13354 : _13349;
    assign _13356 = _13355[62:0];
    assign _13358 = { _13356,
                      _13357 };
    assign _13359 = _13358 < _12272;
    assign _13360 = ~ _13359;
    assign _13348 = _12852[8:8];
    assign _13345 = _13340 - _12272;
    assign _13346 = _13342 ? _13345 : _13340;
    assign _13347 = _13346[62:0];
    assign _13349 = { _13347,
                      _13348 };
    assign _13350 = _13349 < _12272;
    assign _13351 = ~ _13350;
    assign _13339 = _12852[9:9];
    assign _13336 = _13331 - _12272;
    assign _13337 = _13333 ? _13336 : _13331;
    assign _13338 = _13337[62:0];
    assign _13340 = { _13338,
                      _13339 };
    assign _13341 = _13340 < _12272;
    assign _13342 = ~ _13341;
    assign _13330 = _12852[10:10];
    assign _13327 = _13322 - _12272;
    assign _13328 = _13324 ? _13327 : _13322;
    assign _13329 = _13328[62:0];
    assign _13331 = { _13329,
                      _13330 };
    assign _13332 = _13331 < _12272;
    assign _13333 = ~ _13332;
    assign _13321 = _12852[11:11];
    assign _13318 = _13313 - _12272;
    assign _13319 = _13315 ? _13318 : _13313;
    assign _13320 = _13319[62:0];
    assign _13322 = { _13320,
                      _13321 };
    assign _13323 = _13322 < _12272;
    assign _13324 = ~ _13323;
    assign _13312 = _12852[12:12];
    assign _13309 = _13304 - _12272;
    assign _13310 = _13306 ? _13309 : _13304;
    assign _13311 = _13310[62:0];
    assign _13313 = { _13311,
                      _13312 };
    assign _13314 = _13313 < _12272;
    assign _13315 = ~ _13314;
    assign _13303 = _12852[13:13];
    assign _13300 = _13295 - _12272;
    assign _13301 = _13297 ? _13300 : _13295;
    assign _13302 = _13301[62:0];
    assign _13304 = { _13302,
                      _13303 };
    assign _13305 = _13304 < _12272;
    assign _13306 = ~ _13305;
    assign _13294 = _12852[14:14];
    assign _13291 = _13286 - _12272;
    assign _13292 = _13288 ? _13291 : _13286;
    assign _13293 = _13292[62:0];
    assign _13295 = { _13293,
                      _13294 };
    assign _13296 = _13295 < _12272;
    assign _13297 = ~ _13296;
    assign _13285 = _12852[15:15];
    assign _13282 = _13277 - _12272;
    assign _13283 = _13279 ? _13282 : _13277;
    assign _13284 = _13283[62:0];
    assign _13286 = { _13284,
                      _13285 };
    assign _13287 = _13286 < _12272;
    assign _13288 = ~ _13287;
    assign _13276 = _12852[16:16];
    assign _13273 = _13268 - _12272;
    assign _13274 = _13270 ? _13273 : _13268;
    assign _13275 = _13274[62:0];
    assign _13277 = { _13275,
                      _13276 };
    assign _13278 = _13277 < _12272;
    assign _13279 = ~ _13278;
    assign _13267 = _12852[17:17];
    assign _13264 = _13259 - _12272;
    assign _13265 = _13261 ? _13264 : _13259;
    assign _13266 = _13265[62:0];
    assign _13268 = { _13266,
                      _13267 };
    assign _13269 = _13268 < _12272;
    assign _13270 = ~ _13269;
    assign _13258 = _12852[18:18];
    assign _13255 = _13250 - _12272;
    assign _13256 = _13252 ? _13255 : _13250;
    assign _13257 = _13256[62:0];
    assign _13259 = { _13257,
                      _13258 };
    assign _13260 = _13259 < _12272;
    assign _13261 = ~ _13260;
    assign _13249 = _12852[19:19];
    assign _13246 = _13241 - _12272;
    assign _13247 = _13243 ? _13246 : _13241;
    assign _13248 = _13247[62:0];
    assign _13250 = { _13248,
                      _13249 };
    assign _13251 = _13250 < _12272;
    assign _13252 = ~ _13251;
    assign _13240 = _12852[20:20];
    assign _13237 = _13232 - _12272;
    assign _13238 = _13234 ? _13237 : _13232;
    assign _13239 = _13238[62:0];
    assign _13241 = { _13239,
                      _13240 };
    assign _13242 = _13241 < _12272;
    assign _13243 = ~ _13242;
    assign _13231 = _12852[21:21];
    assign _13228 = _13223 - _12272;
    assign _13229 = _13225 ? _13228 : _13223;
    assign _13230 = _13229[62:0];
    assign _13232 = { _13230,
                      _13231 };
    assign _13233 = _13232 < _12272;
    assign _13234 = ~ _13233;
    assign _13222 = _12852[22:22];
    assign _13219 = _13214 - _12272;
    assign _13220 = _13216 ? _13219 : _13214;
    assign _13221 = _13220[62:0];
    assign _13223 = { _13221,
                      _13222 };
    assign _13224 = _13223 < _12272;
    assign _13225 = ~ _13224;
    assign _13213 = _12852[23:23];
    assign _13210 = _13205 - _12272;
    assign _13211 = _13207 ? _13210 : _13205;
    assign _13212 = _13211[62:0];
    assign _13214 = { _13212,
                      _13213 };
    assign _13215 = _13214 < _12272;
    assign _13216 = ~ _13215;
    assign _13204 = _12852[24:24];
    assign _13201 = _13196 - _12272;
    assign _13202 = _13198 ? _13201 : _13196;
    assign _13203 = _13202[62:0];
    assign _13205 = { _13203,
                      _13204 };
    assign _13206 = _13205 < _12272;
    assign _13207 = ~ _13206;
    assign _13195 = _12852[25:25];
    assign _13192 = _13187 - _12272;
    assign _13193 = _13189 ? _13192 : _13187;
    assign _13194 = _13193[62:0];
    assign _13196 = { _13194,
                      _13195 };
    assign _13197 = _13196 < _12272;
    assign _13198 = ~ _13197;
    assign _13186 = _12852[26:26];
    assign _13183 = _13178 - _12272;
    assign _13184 = _13180 ? _13183 : _13178;
    assign _13185 = _13184[62:0];
    assign _13187 = { _13185,
                      _13186 };
    assign _13188 = _13187 < _12272;
    assign _13189 = ~ _13188;
    assign _13177 = _12852[27:27];
    assign _13174 = _13169 - _12272;
    assign _13175 = _13171 ? _13174 : _13169;
    assign _13176 = _13175[62:0];
    assign _13178 = { _13176,
                      _13177 };
    assign _13179 = _13178 < _12272;
    assign _13180 = ~ _13179;
    assign _13168 = _12852[28:28];
    assign _13165 = _13160 - _12272;
    assign _13166 = _13162 ? _13165 : _13160;
    assign _13167 = _13166[62:0];
    assign _13169 = { _13167,
                      _13168 };
    assign _13170 = _13169 < _12272;
    assign _13171 = ~ _13170;
    assign _13159 = _12852[29:29];
    assign _13156 = _13151 - _12272;
    assign _13157 = _13153 ? _13156 : _13151;
    assign _13158 = _13157[62:0];
    assign _13160 = { _13158,
                      _13159 };
    assign _13161 = _13160 < _12272;
    assign _13162 = ~ _13161;
    assign _13150 = _12852[30:30];
    assign _13147 = _13142 - _12272;
    assign _13148 = _13144 ? _13147 : _13142;
    assign _13149 = _13148[62:0];
    assign _13151 = { _13149,
                      _13150 };
    assign _13152 = _13151 < _12272;
    assign _13153 = ~ _13152;
    assign _13141 = _12852[31:31];
    assign _13138 = _13133 - _12272;
    assign _13139 = _13135 ? _13138 : _13133;
    assign _13140 = _13139[62:0];
    assign _13142 = { _13140,
                      _13141 };
    assign _13143 = _13142 < _12272;
    assign _13144 = ~ _13143;
    assign _13132 = _12852[32:32];
    assign _13129 = _13124 - _12272;
    assign _13130 = _13126 ? _13129 : _13124;
    assign _13131 = _13130[62:0];
    assign _13133 = { _13131,
                      _13132 };
    assign _13134 = _13133 < _12272;
    assign _13135 = ~ _13134;
    assign _13123 = _12852[33:33];
    assign _13120 = _13115 - _12272;
    assign _13121 = _13117 ? _13120 : _13115;
    assign _13122 = _13121[62:0];
    assign _13124 = { _13122,
                      _13123 };
    assign _13125 = _13124 < _12272;
    assign _13126 = ~ _13125;
    assign _13114 = _12852[34:34];
    assign _13111 = _13106 - _12272;
    assign _13112 = _13108 ? _13111 : _13106;
    assign _13113 = _13112[62:0];
    assign _13115 = { _13113,
                      _13114 };
    assign _13116 = _13115 < _12272;
    assign _13117 = ~ _13116;
    assign _13105 = _12852[35:35];
    assign _13102 = _13097 - _12272;
    assign _13103 = _13099 ? _13102 : _13097;
    assign _13104 = _13103[62:0];
    assign _13106 = { _13104,
                      _13105 };
    assign _13107 = _13106 < _12272;
    assign _13108 = ~ _13107;
    assign _13096 = _12852[36:36];
    assign _13093 = _13088 - _12272;
    assign _13094 = _13090 ? _13093 : _13088;
    assign _13095 = _13094[62:0];
    assign _13097 = { _13095,
                      _13096 };
    assign _13098 = _13097 < _12272;
    assign _13099 = ~ _13098;
    assign _13087 = _12852[37:37];
    assign _13084 = _13079 - _12272;
    assign _13085 = _13081 ? _13084 : _13079;
    assign _13086 = _13085[62:0];
    assign _13088 = { _13086,
                      _13087 };
    assign _13089 = _13088 < _12272;
    assign _13090 = ~ _13089;
    assign _13078 = _12852[38:38];
    assign _13075 = _13070 - _12272;
    assign _13076 = _13072 ? _13075 : _13070;
    assign _13077 = _13076[62:0];
    assign _13079 = { _13077,
                      _13078 };
    assign _13080 = _13079 < _12272;
    assign _13081 = ~ _13080;
    assign _13069 = _12852[39:39];
    assign _13066 = _13061 - _12272;
    assign _13067 = _13063 ? _13066 : _13061;
    assign _13068 = _13067[62:0];
    assign _13070 = { _13068,
                      _13069 };
    assign _13071 = _13070 < _12272;
    assign _13072 = ~ _13071;
    assign _13060 = _12852[40:40];
    assign _13057 = _13052 - _12272;
    assign _13058 = _13054 ? _13057 : _13052;
    assign _13059 = _13058[62:0];
    assign _13061 = { _13059,
                      _13060 };
    assign _13062 = _13061 < _12272;
    assign _13063 = ~ _13062;
    assign _13051 = _12852[41:41];
    assign _13048 = _13043 - _12272;
    assign _13049 = _13045 ? _13048 : _13043;
    assign _13050 = _13049[62:0];
    assign _13052 = { _13050,
                      _13051 };
    assign _13053 = _13052 < _12272;
    assign _13054 = ~ _13053;
    assign _13042 = _12852[42:42];
    assign _13039 = _13034 - _12272;
    assign _13040 = _13036 ? _13039 : _13034;
    assign _13041 = _13040[62:0];
    assign _13043 = { _13041,
                      _13042 };
    assign _13044 = _13043 < _12272;
    assign _13045 = ~ _13044;
    assign _13033 = _12852[43:43];
    assign _13030 = _13025 - _12272;
    assign _13031 = _13027 ? _13030 : _13025;
    assign _13032 = _13031[62:0];
    assign _13034 = { _13032,
                      _13033 };
    assign _13035 = _13034 < _12272;
    assign _13036 = ~ _13035;
    assign _13024 = _12852[44:44];
    assign _13021 = _13016 - _12272;
    assign _13022 = _13018 ? _13021 : _13016;
    assign _13023 = _13022[62:0];
    assign _13025 = { _13023,
                      _13024 };
    assign _13026 = _13025 < _12272;
    assign _13027 = ~ _13026;
    assign _13015 = _12852[45:45];
    assign _13012 = _13007 - _12272;
    assign _13013 = _13009 ? _13012 : _13007;
    assign _13014 = _13013[62:0];
    assign _13016 = { _13014,
                      _13015 };
    assign _13017 = _13016 < _12272;
    assign _13018 = ~ _13017;
    assign _13006 = _12852[46:46];
    assign _13003 = _12998 - _12272;
    assign _13004 = _13000 ? _13003 : _12998;
    assign _13005 = _13004[62:0];
    assign _13007 = { _13005,
                      _13006 };
    assign _13008 = _13007 < _12272;
    assign _13009 = ~ _13008;
    assign _12997 = _12852[47:47];
    assign _12994 = _12989 - _12272;
    assign _12995 = _12991 ? _12994 : _12989;
    assign _12996 = _12995[62:0];
    assign _12998 = { _12996,
                      _12997 };
    assign _12999 = _12998 < _12272;
    assign _13000 = ~ _12999;
    assign _12988 = _12852[48:48];
    assign _12985 = _12980 - _12272;
    assign _12986 = _12982 ? _12985 : _12980;
    assign _12987 = _12986[62:0];
    assign _12989 = { _12987,
                      _12988 };
    assign _12990 = _12989 < _12272;
    assign _12991 = ~ _12990;
    assign _12979 = _12852[49:49];
    assign _12976 = _12971 - _12272;
    assign _12977 = _12973 ? _12976 : _12971;
    assign _12978 = _12977[62:0];
    assign _12980 = { _12978,
                      _12979 };
    assign _12981 = _12980 < _12272;
    assign _12982 = ~ _12981;
    assign _12970 = _12852[50:50];
    assign _12967 = _12962 - _12272;
    assign _12968 = _12964 ? _12967 : _12962;
    assign _12969 = _12968[62:0];
    assign _12971 = { _12969,
                      _12970 };
    assign _12972 = _12971 < _12272;
    assign _12973 = ~ _12972;
    assign _12961 = _12852[51:51];
    assign _12958 = _12953 - _12272;
    assign _12959 = _12955 ? _12958 : _12953;
    assign _12960 = _12959[62:0];
    assign _12962 = { _12960,
                      _12961 };
    assign _12963 = _12962 < _12272;
    assign _12964 = ~ _12963;
    assign _12952 = _12852[52:52];
    assign _12949 = _12944 - _12272;
    assign _12950 = _12946 ? _12949 : _12944;
    assign _12951 = _12950[62:0];
    assign _12953 = { _12951,
                      _12952 };
    assign _12954 = _12953 < _12272;
    assign _12955 = ~ _12954;
    assign _12943 = _12852[53:53];
    assign _12940 = _12935 - _12272;
    assign _12941 = _12937 ? _12940 : _12935;
    assign _12942 = _12941[62:0];
    assign _12944 = { _12942,
                      _12943 };
    assign _12945 = _12944 < _12272;
    assign _12946 = ~ _12945;
    assign _12934 = _12852[54:54];
    assign _12931 = _12926 - _12272;
    assign _12932 = _12928 ? _12931 : _12926;
    assign _12933 = _12932[62:0];
    assign _12935 = { _12933,
                      _12934 };
    assign _12936 = _12935 < _12272;
    assign _12937 = ~ _12936;
    assign _12925 = _12852[55:55];
    assign _12922 = _12917 - _12272;
    assign _12923 = _12919 ? _12922 : _12917;
    assign _12924 = _12923[62:0];
    assign _12926 = { _12924,
                      _12925 };
    assign _12927 = _12926 < _12272;
    assign _12928 = ~ _12927;
    assign _12916 = _12852[56:56];
    assign _12913 = _12908 - _12272;
    assign _12914 = _12910 ? _12913 : _12908;
    assign _12915 = _12914[62:0];
    assign _12917 = { _12915,
                      _12916 };
    assign _12918 = _12917 < _12272;
    assign _12919 = ~ _12918;
    assign _12907 = _12852[57:57];
    assign _12904 = _12899 - _12272;
    assign _12905 = _12901 ? _12904 : _12899;
    assign _12906 = _12905[62:0];
    assign _12908 = { _12906,
                      _12907 };
    assign _12909 = _12908 < _12272;
    assign _12910 = ~ _12909;
    assign _12898 = _12852[58:58];
    assign _12895 = _12890 - _12272;
    assign _12896 = _12892 ? _12895 : _12890;
    assign _12897 = _12896[62:0];
    assign _12899 = { _12897,
                      _12898 };
    assign _12900 = _12899 < _12272;
    assign _12901 = ~ _12900;
    assign _12889 = _12852[59:59];
    assign _12886 = _12881 - _12272;
    assign _12887 = _12883 ? _12886 : _12881;
    assign _12888 = _12887[62:0];
    assign _12890 = { _12888,
                      _12889 };
    assign _12891 = _12890 < _12272;
    assign _12892 = ~ _12891;
    assign _12880 = _12852[60:60];
    assign _12877 = _12872 - _12272;
    assign _12878 = _12874 ? _12877 : _12872;
    assign _12879 = _12878[62:0];
    assign _12881 = { _12879,
                      _12880 };
    assign _12882 = _12881 < _12272;
    assign _12883 = ~ _12882;
    assign _12871 = _12852[61:61];
    assign _12868 = _12863 - _12272;
    assign _12869 = _12865 ? _12868 : _12863;
    assign _12870 = _12869[62:0];
    assign _12872 = { _12870,
                      _12871 };
    assign _12873 = _12872 < _12272;
    assign _12874 = ~ _12873;
    assign _12862 = _12852[62:62];
    assign _12859 = _12854 - _12272;
    assign _12860 = _12856 ? _12859 : _12854;
    assign _12861 = _12860[62:0];
    assign _12863 = { _12861,
                      _12862 };
    assign _12864 = _12863 < _12272;
    assign _12865 = ~ _12864;
    assign _12852 = _12264 - _12846;
    assign _12853 = _12852[63:63];
    assign _12854 = { _22185,
                      _12853 };
    assign _12855 = _12854 < _12272;
    assign _12856 = ~ _12855;
    assign _12857 = { _22185,
                      _12856 };
    assign _12858 = _12857[62:0];
    assign _12866 = { _12858,
                      _12865 };
    assign _12867 = _12866[62:0];
    assign _12875 = { _12867,
                      _12874 };
    assign _12876 = _12875[62:0];
    assign _12884 = { _12876,
                      _12883 };
    assign _12885 = _12884[62:0];
    assign _12893 = { _12885,
                      _12892 };
    assign _12894 = _12893[62:0];
    assign _12902 = { _12894,
                      _12901 };
    assign _12903 = _12902[62:0];
    assign _12911 = { _12903,
                      _12910 };
    assign _12912 = _12911[62:0];
    assign _12920 = { _12912,
                      _12919 };
    assign _12921 = _12920[62:0];
    assign _12929 = { _12921,
                      _12928 };
    assign _12930 = _12929[62:0];
    assign _12938 = { _12930,
                      _12937 };
    assign _12939 = _12938[62:0];
    assign _12947 = { _12939,
                      _12946 };
    assign _12948 = _12947[62:0];
    assign _12956 = { _12948,
                      _12955 };
    assign _12957 = _12956[62:0];
    assign _12965 = { _12957,
                      _12964 };
    assign _12966 = _12965[62:0];
    assign _12974 = { _12966,
                      _12973 };
    assign _12975 = _12974[62:0];
    assign _12983 = { _12975,
                      _12982 };
    assign _12984 = _12983[62:0];
    assign _12992 = { _12984,
                      _12991 };
    assign _12993 = _12992[62:0];
    assign _13001 = { _12993,
                      _13000 };
    assign _13002 = _13001[62:0];
    assign _13010 = { _13002,
                      _13009 };
    assign _13011 = _13010[62:0];
    assign _13019 = { _13011,
                      _13018 };
    assign _13020 = _13019[62:0];
    assign _13028 = { _13020,
                      _13027 };
    assign _13029 = _13028[62:0];
    assign _13037 = { _13029,
                      _13036 };
    assign _13038 = _13037[62:0];
    assign _13046 = { _13038,
                      _13045 };
    assign _13047 = _13046[62:0];
    assign _13055 = { _13047,
                      _13054 };
    assign _13056 = _13055[62:0];
    assign _13064 = { _13056,
                      _13063 };
    assign _13065 = _13064[62:0];
    assign _13073 = { _13065,
                      _13072 };
    assign _13074 = _13073[62:0];
    assign _13082 = { _13074,
                      _13081 };
    assign _13083 = _13082[62:0];
    assign _13091 = { _13083,
                      _13090 };
    assign _13092 = _13091[62:0];
    assign _13100 = { _13092,
                      _13099 };
    assign _13101 = _13100[62:0];
    assign _13109 = { _13101,
                      _13108 };
    assign _13110 = _13109[62:0];
    assign _13118 = { _13110,
                      _13117 };
    assign _13119 = _13118[62:0];
    assign _13127 = { _13119,
                      _13126 };
    assign _13128 = _13127[62:0];
    assign _13136 = { _13128,
                      _13135 };
    assign _13137 = _13136[62:0];
    assign _13145 = { _13137,
                      _13144 };
    assign _13146 = _13145[62:0];
    assign _13154 = { _13146,
                      _13153 };
    assign _13155 = _13154[62:0];
    assign _13163 = { _13155,
                      _13162 };
    assign _13164 = _13163[62:0];
    assign _13172 = { _13164,
                      _13171 };
    assign _13173 = _13172[62:0];
    assign _13181 = { _13173,
                      _13180 };
    assign _13182 = _13181[62:0];
    assign _13190 = { _13182,
                      _13189 };
    assign _13191 = _13190[62:0];
    assign _13199 = { _13191,
                      _13198 };
    assign _13200 = _13199[62:0];
    assign _13208 = { _13200,
                      _13207 };
    assign _13209 = _13208[62:0];
    assign _13217 = { _13209,
                      _13216 };
    assign _13218 = _13217[62:0];
    assign _13226 = { _13218,
                      _13225 };
    assign _13227 = _13226[62:0];
    assign _13235 = { _13227,
                      _13234 };
    assign _13236 = _13235[62:0];
    assign _13244 = { _13236,
                      _13243 };
    assign _13245 = _13244[62:0];
    assign _13253 = { _13245,
                      _13252 };
    assign _13254 = _13253[62:0];
    assign _13262 = { _13254,
                      _13261 };
    assign _13263 = _13262[62:0];
    assign _13271 = { _13263,
                      _13270 };
    assign _13272 = _13271[62:0];
    assign _13280 = { _13272,
                      _13279 };
    assign _13281 = _13280[62:0];
    assign _13289 = { _13281,
                      _13288 };
    assign _13290 = _13289[62:0];
    assign _13298 = { _13290,
                      _13297 };
    assign _13299 = _13298[62:0];
    assign _13307 = { _13299,
                      _13306 };
    assign _13308 = _13307[62:0];
    assign _13316 = { _13308,
                      _13315 };
    assign _13317 = _13316[62:0];
    assign _13325 = { _13317,
                      _13324 };
    assign _13326 = _13325[62:0];
    assign _13334 = { _13326,
                      _13333 };
    assign _13335 = _13334[62:0];
    assign _13343 = { _13335,
                      _13342 };
    assign _13344 = _13343[62:0];
    assign _13352 = { _13344,
                      _13351 };
    assign _13353 = _13352[62:0];
    assign _13361 = { _13353,
                      _13360 };
    assign _13362 = _13361[62:0];
    assign _13370 = { _13362,
                      _13369 };
    assign _13371 = _13370[62:0];
    assign _13379 = { _13371,
                      _13378 };
    assign _13380 = _13379[62:0];
    assign _13388 = { _13380,
                      _13387 };
    assign _13389 = _13388[62:0];
    assign _13397 = { _13389,
                      _13396 };
    assign _13398 = _13397[62:0];
    assign _13406 = { _13398,
                      _13405 };
    assign _13407 = _13406[62:0];
    assign _13415 = { _13407,
                      _13414 };
    assign _13416 = _13415[62:0];
    assign _13424 = { _13416,
                      _13423 };
    assign _13426 = _13424 + _22186;
    assign _13427 = _13426 * _12846;
    assign _13428 = _13427[63:0];
    assign _14010 = _13428 + _14009;
    assign _12838 = _12269[0:0];
    assign _12835 = _12830 - _12272;
    assign _12836 = _12832 ? _12835 : _12830;
    assign _12837 = _12836[62:0];
    assign _12839 = { _12837,
                      _12838 };
    assign _12840 = _12839 < _12272;
    assign _12841 = ~ _12840;
    assign _12829 = _12269[1:1];
    assign _12826 = _12821 - _12272;
    assign _12827 = _12823 ? _12826 : _12821;
    assign _12828 = _12827[62:0];
    assign _12830 = { _12828,
                      _12829 };
    assign _12831 = _12830 < _12272;
    assign _12832 = ~ _12831;
    assign _12820 = _12269[2:2];
    assign _12817 = _12812 - _12272;
    assign _12818 = _12814 ? _12817 : _12812;
    assign _12819 = _12818[62:0];
    assign _12821 = { _12819,
                      _12820 };
    assign _12822 = _12821 < _12272;
    assign _12823 = ~ _12822;
    assign _12811 = _12269[3:3];
    assign _12808 = _12803 - _12272;
    assign _12809 = _12805 ? _12808 : _12803;
    assign _12810 = _12809[62:0];
    assign _12812 = { _12810,
                      _12811 };
    assign _12813 = _12812 < _12272;
    assign _12814 = ~ _12813;
    assign _12802 = _12269[4:4];
    assign _12799 = _12794 - _12272;
    assign _12800 = _12796 ? _12799 : _12794;
    assign _12801 = _12800[62:0];
    assign _12803 = { _12801,
                      _12802 };
    assign _12804 = _12803 < _12272;
    assign _12805 = ~ _12804;
    assign _12793 = _12269[5:5];
    assign _12790 = _12785 - _12272;
    assign _12791 = _12787 ? _12790 : _12785;
    assign _12792 = _12791[62:0];
    assign _12794 = { _12792,
                      _12793 };
    assign _12795 = _12794 < _12272;
    assign _12796 = ~ _12795;
    assign _12784 = _12269[6:6];
    assign _12781 = _12776 - _12272;
    assign _12782 = _12778 ? _12781 : _12776;
    assign _12783 = _12782[62:0];
    assign _12785 = { _12783,
                      _12784 };
    assign _12786 = _12785 < _12272;
    assign _12787 = ~ _12786;
    assign _12775 = _12269[7:7];
    assign _12772 = _12767 - _12272;
    assign _12773 = _12769 ? _12772 : _12767;
    assign _12774 = _12773[62:0];
    assign _12776 = { _12774,
                      _12775 };
    assign _12777 = _12776 < _12272;
    assign _12778 = ~ _12777;
    assign _12766 = _12269[8:8];
    assign _12763 = _12758 - _12272;
    assign _12764 = _12760 ? _12763 : _12758;
    assign _12765 = _12764[62:0];
    assign _12767 = { _12765,
                      _12766 };
    assign _12768 = _12767 < _12272;
    assign _12769 = ~ _12768;
    assign _12757 = _12269[9:9];
    assign _12754 = _12749 - _12272;
    assign _12755 = _12751 ? _12754 : _12749;
    assign _12756 = _12755[62:0];
    assign _12758 = { _12756,
                      _12757 };
    assign _12759 = _12758 < _12272;
    assign _12760 = ~ _12759;
    assign _12748 = _12269[10:10];
    assign _12745 = _12740 - _12272;
    assign _12746 = _12742 ? _12745 : _12740;
    assign _12747 = _12746[62:0];
    assign _12749 = { _12747,
                      _12748 };
    assign _12750 = _12749 < _12272;
    assign _12751 = ~ _12750;
    assign _12739 = _12269[11:11];
    assign _12736 = _12731 - _12272;
    assign _12737 = _12733 ? _12736 : _12731;
    assign _12738 = _12737[62:0];
    assign _12740 = { _12738,
                      _12739 };
    assign _12741 = _12740 < _12272;
    assign _12742 = ~ _12741;
    assign _12730 = _12269[12:12];
    assign _12727 = _12722 - _12272;
    assign _12728 = _12724 ? _12727 : _12722;
    assign _12729 = _12728[62:0];
    assign _12731 = { _12729,
                      _12730 };
    assign _12732 = _12731 < _12272;
    assign _12733 = ~ _12732;
    assign _12721 = _12269[13:13];
    assign _12718 = _12713 - _12272;
    assign _12719 = _12715 ? _12718 : _12713;
    assign _12720 = _12719[62:0];
    assign _12722 = { _12720,
                      _12721 };
    assign _12723 = _12722 < _12272;
    assign _12724 = ~ _12723;
    assign _12712 = _12269[14:14];
    assign _12709 = _12704 - _12272;
    assign _12710 = _12706 ? _12709 : _12704;
    assign _12711 = _12710[62:0];
    assign _12713 = { _12711,
                      _12712 };
    assign _12714 = _12713 < _12272;
    assign _12715 = ~ _12714;
    assign _12703 = _12269[15:15];
    assign _12700 = _12695 - _12272;
    assign _12701 = _12697 ? _12700 : _12695;
    assign _12702 = _12701[62:0];
    assign _12704 = { _12702,
                      _12703 };
    assign _12705 = _12704 < _12272;
    assign _12706 = ~ _12705;
    assign _12694 = _12269[16:16];
    assign _12691 = _12686 - _12272;
    assign _12692 = _12688 ? _12691 : _12686;
    assign _12693 = _12692[62:0];
    assign _12695 = { _12693,
                      _12694 };
    assign _12696 = _12695 < _12272;
    assign _12697 = ~ _12696;
    assign _12685 = _12269[17:17];
    assign _12682 = _12677 - _12272;
    assign _12683 = _12679 ? _12682 : _12677;
    assign _12684 = _12683[62:0];
    assign _12686 = { _12684,
                      _12685 };
    assign _12687 = _12686 < _12272;
    assign _12688 = ~ _12687;
    assign _12676 = _12269[18:18];
    assign _12673 = _12668 - _12272;
    assign _12674 = _12670 ? _12673 : _12668;
    assign _12675 = _12674[62:0];
    assign _12677 = { _12675,
                      _12676 };
    assign _12678 = _12677 < _12272;
    assign _12679 = ~ _12678;
    assign _12667 = _12269[19:19];
    assign _12664 = _12659 - _12272;
    assign _12665 = _12661 ? _12664 : _12659;
    assign _12666 = _12665[62:0];
    assign _12668 = { _12666,
                      _12667 };
    assign _12669 = _12668 < _12272;
    assign _12670 = ~ _12669;
    assign _12658 = _12269[20:20];
    assign _12655 = _12650 - _12272;
    assign _12656 = _12652 ? _12655 : _12650;
    assign _12657 = _12656[62:0];
    assign _12659 = { _12657,
                      _12658 };
    assign _12660 = _12659 < _12272;
    assign _12661 = ~ _12660;
    assign _12649 = _12269[21:21];
    assign _12646 = _12641 - _12272;
    assign _12647 = _12643 ? _12646 : _12641;
    assign _12648 = _12647[62:0];
    assign _12650 = { _12648,
                      _12649 };
    assign _12651 = _12650 < _12272;
    assign _12652 = ~ _12651;
    assign _12640 = _12269[22:22];
    assign _12637 = _12632 - _12272;
    assign _12638 = _12634 ? _12637 : _12632;
    assign _12639 = _12638[62:0];
    assign _12641 = { _12639,
                      _12640 };
    assign _12642 = _12641 < _12272;
    assign _12643 = ~ _12642;
    assign _12631 = _12269[23:23];
    assign _12628 = _12623 - _12272;
    assign _12629 = _12625 ? _12628 : _12623;
    assign _12630 = _12629[62:0];
    assign _12632 = { _12630,
                      _12631 };
    assign _12633 = _12632 < _12272;
    assign _12634 = ~ _12633;
    assign _12622 = _12269[24:24];
    assign _12619 = _12614 - _12272;
    assign _12620 = _12616 ? _12619 : _12614;
    assign _12621 = _12620[62:0];
    assign _12623 = { _12621,
                      _12622 };
    assign _12624 = _12623 < _12272;
    assign _12625 = ~ _12624;
    assign _12613 = _12269[25:25];
    assign _12610 = _12605 - _12272;
    assign _12611 = _12607 ? _12610 : _12605;
    assign _12612 = _12611[62:0];
    assign _12614 = { _12612,
                      _12613 };
    assign _12615 = _12614 < _12272;
    assign _12616 = ~ _12615;
    assign _12604 = _12269[26:26];
    assign _12601 = _12596 - _12272;
    assign _12602 = _12598 ? _12601 : _12596;
    assign _12603 = _12602[62:0];
    assign _12605 = { _12603,
                      _12604 };
    assign _12606 = _12605 < _12272;
    assign _12607 = ~ _12606;
    assign _12595 = _12269[27:27];
    assign _12592 = _12587 - _12272;
    assign _12593 = _12589 ? _12592 : _12587;
    assign _12594 = _12593[62:0];
    assign _12596 = { _12594,
                      _12595 };
    assign _12597 = _12596 < _12272;
    assign _12598 = ~ _12597;
    assign _12586 = _12269[28:28];
    assign _12583 = _12578 - _12272;
    assign _12584 = _12580 ? _12583 : _12578;
    assign _12585 = _12584[62:0];
    assign _12587 = { _12585,
                      _12586 };
    assign _12588 = _12587 < _12272;
    assign _12589 = ~ _12588;
    assign _12577 = _12269[29:29];
    assign _12574 = _12569 - _12272;
    assign _12575 = _12571 ? _12574 : _12569;
    assign _12576 = _12575[62:0];
    assign _12578 = { _12576,
                      _12577 };
    assign _12579 = _12578 < _12272;
    assign _12580 = ~ _12579;
    assign _12568 = _12269[30:30];
    assign _12565 = _12560 - _12272;
    assign _12566 = _12562 ? _12565 : _12560;
    assign _12567 = _12566[62:0];
    assign _12569 = { _12567,
                      _12568 };
    assign _12570 = _12569 < _12272;
    assign _12571 = ~ _12570;
    assign _12559 = _12269[31:31];
    assign _12556 = _12551 - _12272;
    assign _12557 = _12553 ? _12556 : _12551;
    assign _12558 = _12557[62:0];
    assign _12560 = { _12558,
                      _12559 };
    assign _12561 = _12560 < _12272;
    assign _12562 = ~ _12561;
    assign _12550 = _12269[32:32];
    assign _12547 = _12542 - _12272;
    assign _12548 = _12544 ? _12547 : _12542;
    assign _12549 = _12548[62:0];
    assign _12551 = { _12549,
                      _12550 };
    assign _12552 = _12551 < _12272;
    assign _12553 = ~ _12552;
    assign _12541 = _12269[33:33];
    assign _12538 = _12533 - _12272;
    assign _12539 = _12535 ? _12538 : _12533;
    assign _12540 = _12539[62:0];
    assign _12542 = { _12540,
                      _12541 };
    assign _12543 = _12542 < _12272;
    assign _12544 = ~ _12543;
    assign _12532 = _12269[34:34];
    assign _12529 = _12524 - _12272;
    assign _12530 = _12526 ? _12529 : _12524;
    assign _12531 = _12530[62:0];
    assign _12533 = { _12531,
                      _12532 };
    assign _12534 = _12533 < _12272;
    assign _12535 = ~ _12534;
    assign _12523 = _12269[35:35];
    assign _12520 = _12515 - _12272;
    assign _12521 = _12517 ? _12520 : _12515;
    assign _12522 = _12521[62:0];
    assign _12524 = { _12522,
                      _12523 };
    assign _12525 = _12524 < _12272;
    assign _12526 = ~ _12525;
    assign _12514 = _12269[36:36];
    assign _12511 = _12506 - _12272;
    assign _12512 = _12508 ? _12511 : _12506;
    assign _12513 = _12512[62:0];
    assign _12515 = { _12513,
                      _12514 };
    assign _12516 = _12515 < _12272;
    assign _12517 = ~ _12516;
    assign _12505 = _12269[37:37];
    assign _12502 = _12497 - _12272;
    assign _12503 = _12499 ? _12502 : _12497;
    assign _12504 = _12503[62:0];
    assign _12506 = { _12504,
                      _12505 };
    assign _12507 = _12506 < _12272;
    assign _12508 = ~ _12507;
    assign _12496 = _12269[38:38];
    assign _12493 = _12488 - _12272;
    assign _12494 = _12490 ? _12493 : _12488;
    assign _12495 = _12494[62:0];
    assign _12497 = { _12495,
                      _12496 };
    assign _12498 = _12497 < _12272;
    assign _12499 = ~ _12498;
    assign _12487 = _12269[39:39];
    assign _12484 = _12479 - _12272;
    assign _12485 = _12481 ? _12484 : _12479;
    assign _12486 = _12485[62:0];
    assign _12488 = { _12486,
                      _12487 };
    assign _12489 = _12488 < _12272;
    assign _12490 = ~ _12489;
    assign _12478 = _12269[40:40];
    assign _12475 = _12470 - _12272;
    assign _12476 = _12472 ? _12475 : _12470;
    assign _12477 = _12476[62:0];
    assign _12479 = { _12477,
                      _12478 };
    assign _12480 = _12479 < _12272;
    assign _12481 = ~ _12480;
    assign _12469 = _12269[41:41];
    assign _12466 = _12461 - _12272;
    assign _12467 = _12463 ? _12466 : _12461;
    assign _12468 = _12467[62:0];
    assign _12470 = { _12468,
                      _12469 };
    assign _12471 = _12470 < _12272;
    assign _12472 = ~ _12471;
    assign _12460 = _12269[42:42];
    assign _12457 = _12452 - _12272;
    assign _12458 = _12454 ? _12457 : _12452;
    assign _12459 = _12458[62:0];
    assign _12461 = { _12459,
                      _12460 };
    assign _12462 = _12461 < _12272;
    assign _12463 = ~ _12462;
    assign _12451 = _12269[43:43];
    assign _12448 = _12443 - _12272;
    assign _12449 = _12445 ? _12448 : _12443;
    assign _12450 = _12449[62:0];
    assign _12452 = { _12450,
                      _12451 };
    assign _12453 = _12452 < _12272;
    assign _12454 = ~ _12453;
    assign _12442 = _12269[44:44];
    assign _12439 = _12434 - _12272;
    assign _12440 = _12436 ? _12439 : _12434;
    assign _12441 = _12440[62:0];
    assign _12443 = { _12441,
                      _12442 };
    assign _12444 = _12443 < _12272;
    assign _12445 = ~ _12444;
    assign _12433 = _12269[45:45];
    assign _12430 = _12425 - _12272;
    assign _12431 = _12427 ? _12430 : _12425;
    assign _12432 = _12431[62:0];
    assign _12434 = { _12432,
                      _12433 };
    assign _12435 = _12434 < _12272;
    assign _12436 = ~ _12435;
    assign _12424 = _12269[46:46];
    assign _12421 = _12416 - _12272;
    assign _12422 = _12418 ? _12421 : _12416;
    assign _12423 = _12422[62:0];
    assign _12425 = { _12423,
                      _12424 };
    assign _12426 = _12425 < _12272;
    assign _12427 = ~ _12426;
    assign _12415 = _12269[47:47];
    assign _12412 = _12407 - _12272;
    assign _12413 = _12409 ? _12412 : _12407;
    assign _12414 = _12413[62:0];
    assign _12416 = { _12414,
                      _12415 };
    assign _12417 = _12416 < _12272;
    assign _12418 = ~ _12417;
    assign _12406 = _12269[48:48];
    assign _12403 = _12398 - _12272;
    assign _12404 = _12400 ? _12403 : _12398;
    assign _12405 = _12404[62:0];
    assign _12407 = { _12405,
                      _12406 };
    assign _12408 = _12407 < _12272;
    assign _12409 = ~ _12408;
    assign _12397 = _12269[49:49];
    assign _12394 = _12389 - _12272;
    assign _12395 = _12391 ? _12394 : _12389;
    assign _12396 = _12395[62:0];
    assign _12398 = { _12396,
                      _12397 };
    assign _12399 = _12398 < _12272;
    assign _12400 = ~ _12399;
    assign _12388 = _12269[50:50];
    assign _12385 = _12380 - _12272;
    assign _12386 = _12382 ? _12385 : _12380;
    assign _12387 = _12386[62:0];
    assign _12389 = { _12387,
                      _12388 };
    assign _12390 = _12389 < _12272;
    assign _12391 = ~ _12390;
    assign _12379 = _12269[51:51];
    assign _12376 = _12371 - _12272;
    assign _12377 = _12373 ? _12376 : _12371;
    assign _12378 = _12377[62:0];
    assign _12380 = { _12378,
                      _12379 };
    assign _12381 = _12380 < _12272;
    assign _12382 = ~ _12381;
    assign _12370 = _12269[52:52];
    assign _12367 = _12362 - _12272;
    assign _12368 = _12364 ? _12367 : _12362;
    assign _12369 = _12368[62:0];
    assign _12371 = { _12369,
                      _12370 };
    assign _12372 = _12371 < _12272;
    assign _12373 = ~ _12372;
    assign _12361 = _12269[53:53];
    assign _12358 = _12353 - _12272;
    assign _12359 = _12355 ? _12358 : _12353;
    assign _12360 = _12359[62:0];
    assign _12362 = { _12360,
                      _12361 };
    assign _12363 = _12362 < _12272;
    assign _12364 = ~ _12363;
    assign _12352 = _12269[54:54];
    assign _12349 = _12344 - _12272;
    assign _12350 = _12346 ? _12349 : _12344;
    assign _12351 = _12350[62:0];
    assign _12353 = { _12351,
                      _12352 };
    assign _12354 = _12353 < _12272;
    assign _12355 = ~ _12354;
    assign _12343 = _12269[55:55];
    assign _12340 = _12335 - _12272;
    assign _12341 = _12337 ? _12340 : _12335;
    assign _12342 = _12341[62:0];
    assign _12344 = { _12342,
                      _12343 };
    assign _12345 = _12344 < _12272;
    assign _12346 = ~ _12345;
    assign _12334 = _12269[56:56];
    assign _12331 = _12326 - _12272;
    assign _12332 = _12328 ? _12331 : _12326;
    assign _12333 = _12332[62:0];
    assign _12335 = { _12333,
                      _12334 };
    assign _12336 = _12335 < _12272;
    assign _12337 = ~ _12336;
    assign _12325 = _12269[57:57];
    assign _12322 = _12317 - _12272;
    assign _12323 = _12319 ? _12322 : _12317;
    assign _12324 = _12323[62:0];
    assign _12326 = { _12324,
                      _12325 };
    assign _12327 = _12326 < _12272;
    assign _12328 = ~ _12327;
    assign _12316 = _12269[58:58];
    assign _12313 = _12308 - _12272;
    assign _12314 = _12310 ? _12313 : _12308;
    assign _12315 = _12314[62:0];
    assign _12317 = { _12315,
                      _12316 };
    assign _12318 = _12317 < _12272;
    assign _12319 = ~ _12318;
    assign _12307 = _12269[59:59];
    assign _12304 = _12299 - _12272;
    assign _12305 = _12301 ? _12304 : _12299;
    assign _12306 = _12305[62:0];
    assign _12308 = { _12306,
                      _12307 };
    assign _12309 = _12308 < _12272;
    assign _12310 = ~ _12309;
    assign _12298 = _12269[60:60];
    assign _12295 = _12290 - _12272;
    assign _12296 = _12292 ? _12295 : _12290;
    assign _12297 = _12296[62:0];
    assign _12299 = { _12297,
                      _12298 };
    assign _12300 = _12299 < _12272;
    assign _12301 = ~ _12300;
    assign _12289 = _12269[61:61];
    assign _12286 = _12281 - _12272;
    assign _12287 = _12283 ? _12286 : _12281;
    assign _12288 = _12287[62:0];
    assign _12290 = { _12288,
                      _12289 };
    assign _12291 = _12290 < _12272;
    assign _12292 = ~ _12291;
    assign _12280 = _12269[62:62];
    assign _12277 = _12271 - _12272;
    assign _12278 = _12274 ? _12277 : _12271;
    assign _12279 = _12278[62:0];
    assign _12281 = { _12279,
                      _12280 };
    assign _12282 = _12281 < _12272;
    assign _12283 = ~ _12282;
    assign _12272 = 64'b0000000000000000000000000000000000000000000000000010011101110101;
    assign _12268 = 64'b0000000000000000000000000000000000000000000000000010011101110100;
    assign _12269 = _3 + _12268;
    assign _12270 = _12269[63:63];
    assign _12271 = { _22185,
                      _12270 };
    assign _12273 = _12271 < _12272;
    assign _12274 = ~ _12273;
    assign _12275 = { _22185,
                      _12274 };
    assign _12276 = _12275[62:0];
    assign _12284 = { _12276,
                      _12283 };
    assign _12285 = _12284[62:0];
    assign _12293 = { _12285,
                      _12292 };
    assign _12294 = _12293[62:0];
    assign _12302 = { _12294,
                      _12301 };
    assign _12303 = _12302[62:0];
    assign _12311 = { _12303,
                      _12310 };
    assign _12312 = _12311[62:0];
    assign _12320 = { _12312,
                      _12319 };
    assign _12321 = _12320[62:0];
    assign _12329 = { _12321,
                      _12328 };
    assign _12330 = _12329[62:0];
    assign _12338 = { _12330,
                      _12337 };
    assign _12339 = _12338[62:0];
    assign _12347 = { _12339,
                      _12346 };
    assign _12348 = _12347[62:0];
    assign _12356 = { _12348,
                      _12355 };
    assign _12357 = _12356[62:0];
    assign _12365 = { _12357,
                      _12364 };
    assign _12366 = _12365[62:0];
    assign _12374 = { _12366,
                      _12373 };
    assign _12375 = _12374[62:0];
    assign _12383 = { _12375,
                      _12382 };
    assign _12384 = _12383[62:0];
    assign _12392 = { _12384,
                      _12391 };
    assign _12393 = _12392[62:0];
    assign _12401 = { _12393,
                      _12400 };
    assign _12402 = _12401[62:0];
    assign _12410 = { _12402,
                      _12409 };
    assign _12411 = _12410[62:0];
    assign _12419 = { _12411,
                      _12418 };
    assign _12420 = _12419[62:0];
    assign _12428 = { _12420,
                      _12427 };
    assign _12429 = _12428[62:0];
    assign _12437 = { _12429,
                      _12436 };
    assign _12438 = _12437[62:0];
    assign _12446 = { _12438,
                      _12445 };
    assign _12447 = _12446[62:0];
    assign _12455 = { _12447,
                      _12454 };
    assign _12456 = _12455[62:0];
    assign _12464 = { _12456,
                      _12463 };
    assign _12465 = _12464[62:0];
    assign _12473 = { _12465,
                      _12472 };
    assign _12474 = _12473[62:0];
    assign _12482 = { _12474,
                      _12481 };
    assign _12483 = _12482[62:0];
    assign _12491 = { _12483,
                      _12490 };
    assign _12492 = _12491[62:0];
    assign _12500 = { _12492,
                      _12499 };
    assign _12501 = _12500[62:0];
    assign _12509 = { _12501,
                      _12508 };
    assign _12510 = _12509[62:0];
    assign _12518 = { _12510,
                      _12517 };
    assign _12519 = _12518[62:0];
    assign _12527 = { _12519,
                      _12526 };
    assign _12528 = _12527[62:0];
    assign _12536 = { _12528,
                      _12535 };
    assign _12537 = _12536[62:0];
    assign _12545 = { _12537,
                      _12544 };
    assign _12546 = _12545[62:0];
    assign _12554 = { _12546,
                      _12553 };
    assign _12555 = _12554[62:0];
    assign _12563 = { _12555,
                      _12562 };
    assign _12564 = _12563[62:0];
    assign _12572 = { _12564,
                      _12571 };
    assign _12573 = _12572[62:0];
    assign _12581 = { _12573,
                      _12580 };
    assign _12582 = _12581[62:0];
    assign _12590 = { _12582,
                      _12589 };
    assign _12591 = _12590[62:0];
    assign _12599 = { _12591,
                      _12598 };
    assign _12600 = _12599[62:0];
    assign _12608 = { _12600,
                      _12607 };
    assign _12609 = _12608[62:0];
    assign _12617 = { _12609,
                      _12616 };
    assign _12618 = _12617[62:0];
    assign _12626 = { _12618,
                      _12625 };
    assign _12627 = _12626[62:0];
    assign _12635 = { _12627,
                      _12634 };
    assign _12636 = _12635[62:0];
    assign _12644 = { _12636,
                      _12643 };
    assign _12645 = _12644[62:0];
    assign _12653 = { _12645,
                      _12652 };
    assign _12654 = _12653[62:0];
    assign _12662 = { _12654,
                      _12661 };
    assign _12663 = _12662[62:0];
    assign _12671 = { _12663,
                      _12670 };
    assign _12672 = _12671[62:0];
    assign _12680 = { _12672,
                      _12679 };
    assign _12681 = _12680[62:0];
    assign _12689 = { _12681,
                      _12688 };
    assign _12690 = _12689[62:0];
    assign _12698 = { _12690,
                      _12697 };
    assign _12699 = _12698[62:0];
    assign _12707 = { _12699,
                      _12706 };
    assign _12708 = _12707[62:0];
    assign _12716 = { _12708,
                      _12715 };
    assign _12717 = _12716[62:0];
    assign _12725 = { _12717,
                      _12724 };
    assign _12726 = _12725[62:0];
    assign _12734 = { _12726,
                      _12733 };
    assign _12735 = _12734[62:0];
    assign _12743 = { _12735,
                      _12742 };
    assign _12744 = _12743[62:0];
    assign _12752 = { _12744,
                      _12751 };
    assign _12753 = _12752[62:0];
    assign _12761 = { _12753,
                      _12760 };
    assign _12762 = _12761[62:0];
    assign _12770 = { _12762,
                      _12769 };
    assign _12771 = _12770[62:0];
    assign _12779 = { _12771,
                      _12778 };
    assign _12780 = _12779[62:0];
    assign _12788 = { _12780,
                      _12787 };
    assign _12789 = _12788[62:0];
    assign _12797 = { _12789,
                      _12796 };
    assign _12798 = _12797[62:0];
    assign _12806 = { _12798,
                      _12805 };
    assign _12807 = _12806[62:0];
    assign _12815 = { _12807,
                      _12814 };
    assign _12816 = _12815[62:0];
    assign _12824 = { _12816,
                      _12823 };
    assign _12825 = _12824[62:0];
    assign _12833 = { _12825,
                      _12832 };
    assign _12834 = _12833[62:0];
    assign _12842 = { _12834,
                      _12841 };
    assign _12843 = _12842 * _12272;
    assign _12844 = _12843[63:0];
    assign _12265 = 64'b0000000000000000000000000000000000000000000000011000101010010010;
    assign _12845 = _12265 < _12844;
    assign _12846 = _12845 ? _12844 : _12265;
    assign _12263 = _5 < _19267;
    assign _12264 = _12263 ? _5 : _19267;
    assign _12847 = _12264 < _12846;
    assign _12848 = ~ _12847;
    assign _14011 = _12848 ? _14010 : _21604;
    assign _12252 = _11683[0:0];
    assign _12249 = _12244 - _22192;
    assign _12250 = _12246 ? _12249 : _12244;
    assign _12251 = _12250[62:0];
    assign _12253 = { _12251,
                      _12252 };
    assign _12254 = _12253 < _22192;
    assign _12255 = ~ _12254;
    assign _12243 = _11683[1:1];
    assign _12240 = _12235 - _22192;
    assign _12241 = _12237 ? _12240 : _12235;
    assign _12242 = _12241[62:0];
    assign _12244 = { _12242,
                      _12243 };
    assign _12245 = _12244 < _22192;
    assign _12246 = ~ _12245;
    assign _12234 = _11683[2:2];
    assign _12231 = _12226 - _22192;
    assign _12232 = _12228 ? _12231 : _12226;
    assign _12233 = _12232[62:0];
    assign _12235 = { _12233,
                      _12234 };
    assign _12236 = _12235 < _22192;
    assign _12237 = ~ _12236;
    assign _12225 = _11683[3:3];
    assign _12222 = _12217 - _22192;
    assign _12223 = _12219 ? _12222 : _12217;
    assign _12224 = _12223[62:0];
    assign _12226 = { _12224,
                      _12225 };
    assign _12227 = _12226 < _22192;
    assign _12228 = ~ _12227;
    assign _12216 = _11683[4:4];
    assign _12213 = _12208 - _22192;
    assign _12214 = _12210 ? _12213 : _12208;
    assign _12215 = _12214[62:0];
    assign _12217 = { _12215,
                      _12216 };
    assign _12218 = _12217 < _22192;
    assign _12219 = ~ _12218;
    assign _12207 = _11683[5:5];
    assign _12204 = _12199 - _22192;
    assign _12205 = _12201 ? _12204 : _12199;
    assign _12206 = _12205[62:0];
    assign _12208 = { _12206,
                      _12207 };
    assign _12209 = _12208 < _22192;
    assign _12210 = ~ _12209;
    assign _12198 = _11683[6:6];
    assign _12195 = _12190 - _22192;
    assign _12196 = _12192 ? _12195 : _12190;
    assign _12197 = _12196[62:0];
    assign _12199 = { _12197,
                      _12198 };
    assign _12200 = _12199 < _22192;
    assign _12201 = ~ _12200;
    assign _12189 = _11683[7:7];
    assign _12186 = _12181 - _22192;
    assign _12187 = _12183 ? _12186 : _12181;
    assign _12188 = _12187[62:0];
    assign _12190 = { _12188,
                      _12189 };
    assign _12191 = _12190 < _22192;
    assign _12192 = ~ _12191;
    assign _12180 = _11683[8:8];
    assign _12177 = _12172 - _22192;
    assign _12178 = _12174 ? _12177 : _12172;
    assign _12179 = _12178[62:0];
    assign _12181 = { _12179,
                      _12180 };
    assign _12182 = _12181 < _22192;
    assign _12183 = ~ _12182;
    assign _12171 = _11683[9:9];
    assign _12168 = _12163 - _22192;
    assign _12169 = _12165 ? _12168 : _12163;
    assign _12170 = _12169[62:0];
    assign _12172 = { _12170,
                      _12171 };
    assign _12173 = _12172 < _22192;
    assign _12174 = ~ _12173;
    assign _12162 = _11683[10:10];
    assign _12159 = _12154 - _22192;
    assign _12160 = _12156 ? _12159 : _12154;
    assign _12161 = _12160[62:0];
    assign _12163 = { _12161,
                      _12162 };
    assign _12164 = _12163 < _22192;
    assign _12165 = ~ _12164;
    assign _12153 = _11683[11:11];
    assign _12150 = _12145 - _22192;
    assign _12151 = _12147 ? _12150 : _12145;
    assign _12152 = _12151[62:0];
    assign _12154 = { _12152,
                      _12153 };
    assign _12155 = _12154 < _22192;
    assign _12156 = ~ _12155;
    assign _12144 = _11683[12:12];
    assign _12141 = _12136 - _22192;
    assign _12142 = _12138 ? _12141 : _12136;
    assign _12143 = _12142[62:0];
    assign _12145 = { _12143,
                      _12144 };
    assign _12146 = _12145 < _22192;
    assign _12147 = ~ _12146;
    assign _12135 = _11683[13:13];
    assign _12132 = _12127 - _22192;
    assign _12133 = _12129 ? _12132 : _12127;
    assign _12134 = _12133[62:0];
    assign _12136 = { _12134,
                      _12135 };
    assign _12137 = _12136 < _22192;
    assign _12138 = ~ _12137;
    assign _12126 = _11683[14:14];
    assign _12123 = _12118 - _22192;
    assign _12124 = _12120 ? _12123 : _12118;
    assign _12125 = _12124[62:0];
    assign _12127 = { _12125,
                      _12126 };
    assign _12128 = _12127 < _22192;
    assign _12129 = ~ _12128;
    assign _12117 = _11683[15:15];
    assign _12114 = _12109 - _22192;
    assign _12115 = _12111 ? _12114 : _12109;
    assign _12116 = _12115[62:0];
    assign _12118 = { _12116,
                      _12117 };
    assign _12119 = _12118 < _22192;
    assign _12120 = ~ _12119;
    assign _12108 = _11683[16:16];
    assign _12105 = _12100 - _22192;
    assign _12106 = _12102 ? _12105 : _12100;
    assign _12107 = _12106[62:0];
    assign _12109 = { _12107,
                      _12108 };
    assign _12110 = _12109 < _22192;
    assign _12111 = ~ _12110;
    assign _12099 = _11683[17:17];
    assign _12096 = _12091 - _22192;
    assign _12097 = _12093 ? _12096 : _12091;
    assign _12098 = _12097[62:0];
    assign _12100 = { _12098,
                      _12099 };
    assign _12101 = _12100 < _22192;
    assign _12102 = ~ _12101;
    assign _12090 = _11683[18:18];
    assign _12087 = _12082 - _22192;
    assign _12088 = _12084 ? _12087 : _12082;
    assign _12089 = _12088[62:0];
    assign _12091 = { _12089,
                      _12090 };
    assign _12092 = _12091 < _22192;
    assign _12093 = ~ _12092;
    assign _12081 = _11683[19:19];
    assign _12078 = _12073 - _22192;
    assign _12079 = _12075 ? _12078 : _12073;
    assign _12080 = _12079[62:0];
    assign _12082 = { _12080,
                      _12081 };
    assign _12083 = _12082 < _22192;
    assign _12084 = ~ _12083;
    assign _12072 = _11683[20:20];
    assign _12069 = _12064 - _22192;
    assign _12070 = _12066 ? _12069 : _12064;
    assign _12071 = _12070[62:0];
    assign _12073 = { _12071,
                      _12072 };
    assign _12074 = _12073 < _22192;
    assign _12075 = ~ _12074;
    assign _12063 = _11683[21:21];
    assign _12060 = _12055 - _22192;
    assign _12061 = _12057 ? _12060 : _12055;
    assign _12062 = _12061[62:0];
    assign _12064 = { _12062,
                      _12063 };
    assign _12065 = _12064 < _22192;
    assign _12066 = ~ _12065;
    assign _12054 = _11683[22:22];
    assign _12051 = _12046 - _22192;
    assign _12052 = _12048 ? _12051 : _12046;
    assign _12053 = _12052[62:0];
    assign _12055 = { _12053,
                      _12054 };
    assign _12056 = _12055 < _22192;
    assign _12057 = ~ _12056;
    assign _12045 = _11683[23:23];
    assign _12042 = _12037 - _22192;
    assign _12043 = _12039 ? _12042 : _12037;
    assign _12044 = _12043[62:0];
    assign _12046 = { _12044,
                      _12045 };
    assign _12047 = _12046 < _22192;
    assign _12048 = ~ _12047;
    assign _12036 = _11683[24:24];
    assign _12033 = _12028 - _22192;
    assign _12034 = _12030 ? _12033 : _12028;
    assign _12035 = _12034[62:0];
    assign _12037 = { _12035,
                      _12036 };
    assign _12038 = _12037 < _22192;
    assign _12039 = ~ _12038;
    assign _12027 = _11683[25:25];
    assign _12024 = _12019 - _22192;
    assign _12025 = _12021 ? _12024 : _12019;
    assign _12026 = _12025[62:0];
    assign _12028 = { _12026,
                      _12027 };
    assign _12029 = _12028 < _22192;
    assign _12030 = ~ _12029;
    assign _12018 = _11683[26:26];
    assign _12015 = _12010 - _22192;
    assign _12016 = _12012 ? _12015 : _12010;
    assign _12017 = _12016[62:0];
    assign _12019 = { _12017,
                      _12018 };
    assign _12020 = _12019 < _22192;
    assign _12021 = ~ _12020;
    assign _12009 = _11683[27:27];
    assign _12006 = _12001 - _22192;
    assign _12007 = _12003 ? _12006 : _12001;
    assign _12008 = _12007[62:0];
    assign _12010 = { _12008,
                      _12009 };
    assign _12011 = _12010 < _22192;
    assign _12012 = ~ _12011;
    assign _12000 = _11683[28:28];
    assign _11997 = _11992 - _22192;
    assign _11998 = _11994 ? _11997 : _11992;
    assign _11999 = _11998[62:0];
    assign _12001 = { _11999,
                      _12000 };
    assign _12002 = _12001 < _22192;
    assign _12003 = ~ _12002;
    assign _11991 = _11683[29:29];
    assign _11988 = _11983 - _22192;
    assign _11989 = _11985 ? _11988 : _11983;
    assign _11990 = _11989[62:0];
    assign _11992 = { _11990,
                      _11991 };
    assign _11993 = _11992 < _22192;
    assign _11994 = ~ _11993;
    assign _11982 = _11683[30:30];
    assign _11979 = _11974 - _22192;
    assign _11980 = _11976 ? _11979 : _11974;
    assign _11981 = _11980[62:0];
    assign _11983 = { _11981,
                      _11982 };
    assign _11984 = _11983 < _22192;
    assign _11985 = ~ _11984;
    assign _11973 = _11683[31:31];
    assign _11970 = _11965 - _22192;
    assign _11971 = _11967 ? _11970 : _11965;
    assign _11972 = _11971[62:0];
    assign _11974 = { _11972,
                      _11973 };
    assign _11975 = _11974 < _22192;
    assign _11976 = ~ _11975;
    assign _11964 = _11683[32:32];
    assign _11961 = _11956 - _22192;
    assign _11962 = _11958 ? _11961 : _11956;
    assign _11963 = _11962[62:0];
    assign _11965 = { _11963,
                      _11964 };
    assign _11966 = _11965 < _22192;
    assign _11967 = ~ _11966;
    assign _11955 = _11683[33:33];
    assign _11952 = _11947 - _22192;
    assign _11953 = _11949 ? _11952 : _11947;
    assign _11954 = _11953[62:0];
    assign _11956 = { _11954,
                      _11955 };
    assign _11957 = _11956 < _22192;
    assign _11958 = ~ _11957;
    assign _11946 = _11683[34:34];
    assign _11943 = _11938 - _22192;
    assign _11944 = _11940 ? _11943 : _11938;
    assign _11945 = _11944[62:0];
    assign _11947 = { _11945,
                      _11946 };
    assign _11948 = _11947 < _22192;
    assign _11949 = ~ _11948;
    assign _11937 = _11683[35:35];
    assign _11934 = _11929 - _22192;
    assign _11935 = _11931 ? _11934 : _11929;
    assign _11936 = _11935[62:0];
    assign _11938 = { _11936,
                      _11937 };
    assign _11939 = _11938 < _22192;
    assign _11940 = ~ _11939;
    assign _11928 = _11683[36:36];
    assign _11925 = _11920 - _22192;
    assign _11926 = _11922 ? _11925 : _11920;
    assign _11927 = _11926[62:0];
    assign _11929 = { _11927,
                      _11928 };
    assign _11930 = _11929 < _22192;
    assign _11931 = ~ _11930;
    assign _11919 = _11683[37:37];
    assign _11916 = _11911 - _22192;
    assign _11917 = _11913 ? _11916 : _11911;
    assign _11918 = _11917[62:0];
    assign _11920 = { _11918,
                      _11919 };
    assign _11921 = _11920 < _22192;
    assign _11922 = ~ _11921;
    assign _11910 = _11683[38:38];
    assign _11907 = _11902 - _22192;
    assign _11908 = _11904 ? _11907 : _11902;
    assign _11909 = _11908[62:0];
    assign _11911 = { _11909,
                      _11910 };
    assign _11912 = _11911 < _22192;
    assign _11913 = ~ _11912;
    assign _11901 = _11683[39:39];
    assign _11898 = _11893 - _22192;
    assign _11899 = _11895 ? _11898 : _11893;
    assign _11900 = _11899[62:0];
    assign _11902 = { _11900,
                      _11901 };
    assign _11903 = _11902 < _22192;
    assign _11904 = ~ _11903;
    assign _11892 = _11683[40:40];
    assign _11889 = _11884 - _22192;
    assign _11890 = _11886 ? _11889 : _11884;
    assign _11891 = _11890[62:0];
    assign _11893 = { _11891,
                      _11892 };
    assign _11894 = _11893 < _22192;
    assign _11895 = ~ _11894;
    assign _11883 = _11683[41:41];
    assign _11880 = _11875 - _22192;
    assign _11881 = _11877 ? _11880 : _11875;
    assign _11882 = _11881[62:0];
    assign _11884 = { _11882,
                      _11883 };
    assign _11885 = _11884 < _22192;
    assign _11886 = ~ _11885;
    assign _11874 = _11683[42:42];
    assign _11871 = _11866 - _22192;
    assign _11872 = _11868 ? _11871 : _11866;
    assign _11873 = _11872[62:0];
    assign _11875 = { _11873,
                      _11874 };
    assign _11876 = _11875 < _22192;
    assign _11877 = ~ _11876;
    assign _11865 = _11683[43:43];
    assign _11862 = _11857 - _22192;
    assign _11863 = _11859 ? _11862 : _11857;
    assign _11864 = _11863[62:0];
    assign _11866 = { _11864,
                      _11865 };
    assign _11867 = _11866 < _22192;
    assign _11868 = ~ _11867;
    assign _11856 = _11683[44:44];
    assign _11853 = _11848 - _22192;
    assign _11854 = _11850 ? _11853 : _11848;
    assign _11855 = _11854[62:0];
    assign _11857 = { _11855,
                      _11856 };
    assign _11858 = _11857 < _22192;
    assign _11859 = ~ _11858;
    assign _11847 = _11683[45:45];
    assign _11844 = _11839 - _22192;
    assign _11845 = _11841 ? _11844 : _11839;
    assign _11846 = _11845[62:0];
    assign _11848 = { _11846,
                      _11847 };
    assign _11849 = _11848 < _22192;
    assign _11850 = ~ _11849;
    assign _11838 = _11683[46:46];
    assign _11835 = _11830 - _22192;
    assign _11836 = _11832 ? _11835 : _11830;
    assign _11837 = _11836[62:0];
    assign _11839 = { _11837,
                      _11838 };
    assign _11840 = _11839 < _22192;
    assign _11841 = ~ _11840;
    assign _11829 = _11683[47:47];
    assign _11826 = _11821 - _22192;
    assign _11827 = _11823 ? _11826 : _11821;
    assign _11828 = _11827[62:0];
    assign _11830 = { _11828,
                      _11829 };
    assign _11831 = _11830 < _22192;
    assign _11832 = ~ _11831;
    assign _11820 = _11683[48:48];
    assign _11817 = _11812 - _22192;
    assign _11818 = _11814 ? _11817 : _11812;
    assign _11819 = _11818[62:0];
    assign _11821 = { _11819,
                      _11820 };
    assign _11822 = _11821 < _22192;
    assign _11823 = ~ _11822;
    assign _11811 = _11683[49:49];
    assign _11808 = _11803 - _22192;
    assign _11809 = _11805 ? _11808 : _11803;
    assign _11810 = _11809[62:0];
    assign _11812 = { _11810,
                      _11811 };
    assign _11813 = _11812 < _22192;
    assign _11814 = ~ _11813;
    assign _11802 = _11683[50:50];
    assign _11799 = _11794 - _22192;
    assign _11800 = _11796 ? _11799 : _11794;
    assign _11801 = _11800[62:0];
    assign _11803 = { _11801,
                      _11802 };
    assign _11804 = _11803 < _22192;
    assign _11805 = ~ _11804;
    assign _11793 = _11683[51:51];
    assign _11790 = _11785 - _22192;
    assign _11791 = _11787 ? _11790 : _11785;
    assign _11792 = _11791[62:0];
    assign _11794 = { _11792,
                      _11793 };
    assign _11795 = _11794 < _22192;
    assign _11796 = ~ _11795;
    assign _11784 = _11683[52:52];
    assign _11781 = _11776 - _22192;
    assign _11782 = _11778 ? _11781 : _11776;
    assign _11783 = _11782[62:0];
    assign _11785 = { _11783,
                      _11784 };
    assign _11786 = _11785 < _22192;
    assign _11787 = ~ _11786;
    assign _11775 = _11683[53:53];
    assign _11772 = _11767 - _22192;
    assign _11773 = _11769 ? _11772 : _11767;
    assign _11774 = _11773[62:0];
    assign _11776 = { _11774,
                      _11775 };
    assign _11777 = _11776 < _22192;
    assign _11778 = ~ _11777;
    assign _11766 = _11683[54:54];
    assign _11763 = _11758 - _22192;
    assign _11764 = _11760 ? _11763 : _11758;
    assign _11765 = _11764[62:0];
    assign _11767 = { _11765,
                      _11766 };
    assign _11768 = _11767 < _22192;
    assign _11769 = ~ _11768;
    assign _11757 = _11683[55:55];
    assign _11754 = _11749 - _22192;
    assign _11755 = _11751 ? _11754 : _11749;
    assign _11756 = _11755[62:0];
    assign _11758 = { _11756,
                      _11757 };
    assign _11759 = _11758 < _22192;
    assign _11760 = ~ _11759;
    assign _11748 = _11683[56:56];
    assign _11745 = _11740 - _22192;
    assign _11746 = _11742 ? _11745 : _11740;
    assign _11747 = _11746[62:0];
    assign _11749 = { _11747,
                      _11748 };
    assign _11750 = _11749 < _22192;
    assign _11751 = ~ _11750;
    assign _11739 = _11683[57:57];
    assign _11736 = _11731 - _22192;
    assign _11737 = _11733 ? _11736 : _11731;
    assign _11738 = _11737[62:0];
    assign _11740 = { _11738,
                      _11739 };
    assign _11741 = _11740 < _22192;
    assign _11742 = ~ _11741;
    assign _11730 = _11683[58:58];
    assign _11727 = _11722 - _22192;
    assign _11728 = _11724 ? _11727 : _11722;
    assign _11729 = _11728[62:0];
    assign _11731 = { _11729,
                      _11730 };
    assign _11732 = _11731 < _22192;
    assign _11733 = ~ _11732;
    assign _11721 = _11683[59:59];
    assign _11718 = _11713 - _22192;
    assign _11719 = _11715 ? _11718 : _11713;
    assign _11720 = _11719[62:0];
    assign _11722 = { _11720,
                      _11721 };
    assign _11723 = _11722 < _22192;
    assign _11724 = ~ _11723;
    assign _11712 = _11683[60:60];
    assign _11709 = _11704 - _22192;
    assign _11710 = _11706 ? _11709 : _11704;
    assign _11711 = _11710[62:0];
    assign _11713 = { _11711,
                      _11712 };
    assign _11714 = _11713 < _22192;
    assign _11715 = ~ _11714;
    assign _11703 = _11683[61:61];
    assign _11700 = _11695 - _22192;
    assign _11701 = _11697 ? _11700 : _11695;
    assign _11702 = _11701[62:0];
    assign _11704 = { _11702,
                      _11703 };
    assign _11705 = _11704 < _22192;
    assign _11706 = ~ _11705;
    assign _11694 = _11683[62:62];
    assign _11691 = _11685 - _22192;
    assign _11692 = _11688 ? _11691 : _11685;
    assign _11693 = _11692[62:0];
    assign _11695 = { _11693,
                      _11694 };
    assign _11696 = _11695 < _22192;
    assign _11697 = ~ _11696;
    assign _11681 = _11673 + _22186;
    assign _11682 = _11673 * _11681;
    assign _11683 = _11682[63:0];
    assign _11684 = _11683[63:63];
    assign _11685 = { _22185,
                      _11684 };
    assign _11687 = _11685 < _22192;
    assign _11688 = ~ _11687;
    assign _11689 = { _22185,
                      _11688 };
    assign _11690 = _11689[62:0];
    assign _11698 = { _11690,
                      _11697 };
    assign _11699 = _11698[62:0];
    assign _11707 = { _11699,
                      _11706 };
    assign _11708 = _11707[62:0];
    assign _11716 = { _11708,
                      _11715 };
    assign _11717 = _11716[62:0];
    assign _11725 = { _11717,
                      _11724 };
    assign _11726 = _11725[62:0];
    assign _11734 = { _11726,
                      _11733 };
    assign _11735 = _11734[62:0];
    assign _11743 = { _11735,
                      _11742 };
    assign _11744 = _11743[62:0];
    assign _11752 = { _11744,
                      _11751 };
    assign _11753 = _11752[62:0];
    assign _11761 = { _11753,
                      _11760 };
    assign _11762 = _11761[62:0];
    assign _11770 = { _11762,
                      _11769 };
    assign _11771 = _11770[62:0];
    assign _11779 = { _11771,
                      _11778 };
    assign _11780 = _11779[62:0];
    assign _11788 = { _11780,
                      _11787 };
    assign _11789 = _11788[62:0];
    assign _11797 = { _11789,
                      _11796 };
    assign _11798 = _11797[62:0];
    assign _11806 = { _11798,
                      _11805 };
    assign _11807 = _11806[62:0];
    assign _11815 = { _11807,
                      _11814 };
    assign _11816 = _11815[62:0];
    assign _11824 = { _11816,
                      _11823 };
    assign _11825 = _11824[62:0];
    assign _11833 = { _11825,
                      _11832 };
    assign _11834 = _11833[62:0];
    assign _11842 = { _11834,
                      _11841 };
    assign _11843 = _11842[62:0];
    assign _11851 = { _11843,
                      _11850 };
    assign _11852 = _11851[62:0];
    assign _11860 = { _11852,
                      _11859 };
    assign _11861 = _11860[62:0];
    assign _11869 = { _11861,
                      _11868 };
    assign _11870 = _11869[62:0];
    assign _11878 = { _11870,
                      _11877 };
    assign _11879 = _11878[62:0];
    assign _11887 = { _11879,
                      _11886 };
    assign _11888 = _11887[62:0];
    assign _11896 = { _11888,
                      _11895 };
    assign _11897 = _11896[62:0];
    assign _11905 = { _11897,
                      _11904 };
    assign _11906 = _11905[62:0];
    assign _11914 = { _11906,
                      _11913 };
    assign _11915 = _11914[62:0];
    assign _11923 = { _11915,
                      _11922 };
    assign _11924 = _11923[62:0];
    assign _11932 = { _11924,
                      _11931 };
    assign _11933 = _11932[62:0];
    assign _11941 = { _11933,
                      _11940 };
    assign _11942 = _11941[62:0];
    assign _11950 = { _11942,
                      _11949 };
    assign _11951 = _11950[62:0];
    assign _11959 = { _11951,
                      _11958 };
    assign _11960 = _11959[62:0];
    assign _11968 = { _11960,
                      _11967 };
    assign _11969 = _11968[62:0];
    assign _11977 = { _11969,
                      _11976 };
    assign _11978 = _11977[62:0];
    assign _11986 = { _11978,
                      _11985 };
    assign _11987 = _11986[62:0];
    assign _11995 = { _11987,
                      _11994 };
    assign _11996 = _11995[62:0];
    assign _12004 = { _11996,
                      _12003 };
    assign _12005 = _12004[62:0];
    assign _12013 = { _12005,
                      _12012 };
    assign _12014 = _12013[62:0];
    assign _12022 = { _12014,
                      _12021 };
    assign _12023 = _12022[62:0];
    assign _12031 = { _12023,
                      _12030 };
    assign _12032 = _12031[62:0];
    assign _12040 = { _12032,
                      _12039 };
    assign _12041 = _12040[62:0];
    assign _12049 = { _12041,
                      _12048 };
    assign _12050 = _12049[62:0];
    assign _12058 = { _12050,
                      _12057 };
    assign _12059 = _12058[62:0];
    assign _12067 = { _12059,
                      _12066 };
    assign _12068 = _12067[62:0];
    assign _12076 = { _12068,
                      _12075 };
    assign _12077 = _12076[62:0];
    assign _12085 = { _12077,
                      _12084 };
    assign _12086 = _12085[62:0];
    assign _12094 = { _12086,
                      _12093 };
    assign _12095 = _12094[62:0];
    assign _12103 = { _12095,
                      _12102 };
    assign _12104 = _12103[62:0];
    assign _12112 = { _12104,
                      _12111 };
    assign _12113 = _12112[62:0];
    assign _12121 = { _12113,
                      _12120 };
    assign _12122 = _12121[62:0];
    assign _12130 = { _12122,
                      _12129 };
    assign _12131 = _12130[62:0];
    assign _12139 = { _12131,
                      _12138 };
    assign _12140 = _12139[62:0];
    assign _12148 = { _12140,
                      _12147 };
    assign _12149 = _12148[62:0];
    assign _12157 = { _12149,
                      _12156 };
    assign _12158 = _12157[62:0];
    assign _12166 = { _12158,
                      _12165 };
    assign _12167 = _12166[62:0];
    assign _12175 = { _12167,
                      _12174 };
    assign _12176 = _12175[62:0];
    assign _12184 = { _12176,
                      _12183 };
    assign _12185 = _12184[62:0];
    assign _12193 = { _12185,
                      _12192 };
    assign _12194 = _12193[62:0];
    assign _12202 = { _12194,
                      _12201 };
    assign _12203 = _12202[62:0];
    assign _12211 = { _12203,
                      _12210 };
    assign _12212 = _12211[62:0];
    assign _12220 = { _12212,
                      _12219 };
    assign _12221 = _12220[62:0];
    assign _12229 = { _12221,
                      _12228 };
    assign _12230 = _12229[62:0];
    assign _12238 = { _12230,
                      _12237 };
    assign _12239 = _12238[62:0];
    assign _12247 = { _12239,
                      _12246 };
    assign _12248 = _12247[62:0];
    assign _12256 = { _12248,
                      _12255 };
    assign _12257 = _10521 * _12256;
    assign _12258 = _12257[63:0];
    assign _11669 = _11101[0:0];
    assign _11666 = _11661 - _10521;
    assign _11667 = _11663 ? _11666 : _11661;
    assign _11668 = _11667[62:0];
    assign _11670 = { _11668,
                      _11669 };
    assign _11671 = _11670 < _10521;
    assign _11672 = ~ _11671;
    assign _11660 = _11101[1:1];
    assign _11657 = _11652 - _10521;
    assign _11658 = _11654 ? _11657 : _11652;
    assign _11659 = _11658[62:0];
    assign _11661 = { _11659,
                      _11660 };
    assign _11662 = _11661 < _10521;
    assign _11663 = ~ _11662;
    assign _11651 = _11101[2:2];
    assign _11648 = _11643 - _10521;
    assign _11649 = _11645 ? _11648 : _11643;
    assign _11650 = _11649[62:0];
    assign _11652 = { _11650,
                      _11651 };
    assign _11653 = _11652 < _10521;
    assign _11654 = ~ _11653;
    assign _11642 = _11101[3:3];
    assign _11639 = _11634 - _10521;
    assign _11640 = _11636 ? _11639 : _11634;
    assign _11641 = _11640[62:0];
    assign _11643 = { _11641,
                      _11642 };
    assign _11644 = _11643 < _10521;
    assign _11645 = ~ _11644;
    assign _11633 = _11101[4:4];
    assign _11630 = _11625 - _10521;
    assign _11631 = _11627 ? _11630 : _11625;
    assign _11632 = _11631[62:0];
    assign _11634 = { _11632,
                      _11633 };
    assign _11635 = _11634 < _10521;
    assign _11636 = ~ _11635;
    assign _11624 = _11101[5:5];
    assign _11621 = _11616 - _10521;
    assign _11622 = _11618 ? _11621 : _11616;
    assign _11623 = _11622[62:0];
    assign _11625 = { _11623,
                      _11624 };
    assign _11626 = _11625 < _10521;
    assign _11627 = ~ _11626;
    assign _11615 = _11101[6:6];
    assign _11612 = _11607 - _10521;
    assign _11613 = _11609 ? _11612 : _11607;
    assign _11614 = _11613[62:0];
    assign _11616 = { _11614,
                      _11615 };
    assign _11617 = _11616 < _10521;
    assign _11618 = ~ _11617;
    assign _11606 = _11101[7:7];
    assign _11603 = _11598 - _10521;
    assign _11604 = _11600 ? _11603 : _11598;
    assign _11605 = _11604[62:0];
    assign _11607 = { _11605,
                      _11606 };
    assign _11608 = _11607 < _10521;
    assign _11609 = ~ _11608;
    assign _11597 = _11101[8:8];
    assign _11594 = _11589 - _10521;
    assign _11595 = _11591 ? _11594 : _11589;
    assign _11596 = _11595[62:0];
    assign _11598 = { _11596,
                      _11597 };
    assign _11599 = _11598 < _10521;
    assign _11600 = ~ _11599;
    assign _11588 = _11101[9:9];
    assign _11585 = _11580 - _10521;
    assign _11586 = _11582 ? _11585 : _11580;
    assign _11587 = _11586[62:0];
    assign _11589 = { _11587,
                      _11588 };
    assign _11590 = _11589 < _10521;
    assign _11591 = ~ _11590;
    assign _11579 = _11101[10:10];
    assign _11576 = _11571 - _10521;
    assign _11577 = _11573 ? _11576 : _11571;
    assign _11578 = _11577[62:0];
    assign _11580 = { _11578,
                      _11579 };
    assign _11581 = _11580 < _10521;
    assign _11582 = ~ _11581;
    assign _11570 = _11101[11:11];
    assign _11567 = _11562 - _10521;
    assign _11568 = _11564 ? _11567 : _11562;
    assign _11569 = _11568[62:0];
    assign _11571 = { _11569,
                      _11570 };
    assign _11572 = _11571 < _10521;
    assign _11573 = ~ _11572;
    assign _11561 = _11101[12:12];
    assign _11558 = _11553 - _10521;
    assign _11559 = _11555 ? _11558 : _11553;
    assign _11560 = _11559[62:0];
    assign _11562 = { _11560,
                      _11561 };
    assign _11563 = _11562 < _10521;
    assign _11564 = ~ _11563;
    assign _11552 = _11101[13:13];
    assign _11549 = _11544 - _10521;
    assign _11550 = _11546 ? _11549 : _11544;
    assign _11551 = _11550[62:0];
    assign _11553 = { _11551,
                      _11552 };
    assign _11554 = _11553 < _10521;
    assign _11555 = ~ _11554;
    assign _11543 = _11101[14:14];
    assign _11540 = _11535 - _10521;
    assign _11541 = _11537 ? _11540 : _11535;
    assign _11542 = _11541[62:0];
    assign _11544 = { _11542,
                      _11543 };
    assign _11545 = _11544 < _10521;
    assign _11546 = ~ _11545;
    assign _11534 = _11101[15:15];
    assign _11531 = _11526 - _10521;
    assign _11532 = _11528 ? _11531 : _11526;
    assign _11533 = _11532[62:0];
    assign _11535 = { _11533,
                      _11534 };
    assign _11536 = _11535 < _10521;
    assign _11537 = ~ _11536;
    assign _11525 = _11101[16:16];
    assign _11522 = _11517 - _10521;
    assign _11523 = _11519 ? _11522 : _11517;
    assign _11524 = _11523[62:0];
    assign _11526 = { _11524,
                      _11525 };
    assign _11527 = _11526 < _10521;
    assign _11528 = ~ _11527;
    assign _11516 = _11101[17:17];
    assign _11513 = _11508 - _10521;
    assign _11514 = _11510 ? _11513 : _11508;
    assign _11515 = _11514[62:0];
    assign _11517 = { _11515,
                      _11516 };
    assign _11518 = _11517 < _10521;
    assign _11519 = ~ _11518;
    assign _11507 = _11101[18:18];
    assign _11504 = _11499 - _10521;
    assign _11505 = _11501 ? _11504 : _11499;
    assign _11506 = _11505[62:0];
    assign _11508 = { _11506,
                      _11507 };
    assign _11509 = _11508 < _10521;
    assign _11510 = ~ _11509;
    assign _11498 = _11101[19:19];
    assign _11495 = _11490 - _10521;
    assign _11496 = _11492 ? _11495 : _11490;
    assign _11497 = _11496[62:0];
    assign _11499 = { _11497,
                      _11498 };
    assign _11500 = _11499 < _10521;
    assign _11501 = ~ _11500;
    assign _11489 = _11101[20:20];
    assign _11486 = _11481 - _10521;
    assign _11487 = _11483 ? _11486 : _11481;
    assign _11488 = _11487[62:0];
    assign _11490 = { _11488,
                      _11489 };
    assign _11491 = _11490 < _10521;
    assign _11492 = ~ _11491;
    assign _11480 = _11101[21:21];
    assign _11477 = _11472 - _10521;
    assign _11478 = _11474 ? _11477 : _11472;
    assign _11479 = _11478[62:0];
    assign _11481 = { _11479,
                      _11480 };
    assign _11482 = _11481 < _10521;
    assign _11483 = ~ _11482;
    assign _11471 = _11101[22:22];
    assign _11468 = _11463 - _10521;
    assign _11469 = _11465 ? _11468 : _11463;
    assign _11470 = _11469[62:0];
    assign _11472 = { _11470,
                      _11471 };
    assign _11473 = _11472 < _10521;
    assign _11474 = ~ _11473;
    assign _11462 = _11101[23:23];
    assign _11459 = _11454 - _10521;
    assign _11460 = _11456 ? _11459 : _11454;
    assign _11461 = _11460[62:0];
    assign _11463 = { _11461,
                      _11462 };
    assign _11464 = _11463 < _10521;
    assign _11465 = ~ _11464;
    assign _11453 = _11101[24:24];
    assign _11450 = _11445 - _10521;
    assign _11451 = _11447 ? _11450 : _11445;
    assign _11452 = _11451[62:0];
    assign _11454 = { _11452,
                      _11453 };
    assign _11455 = _11454 < _10521;
    assign _11456 = ~ _11455;
    assign _11444 = _11101[25:25];
    assign _11441 = _11436 - _10521;
    assign _11442 = _11438 ? _11441 : _11436;
    assign _11443 = _11442[62:0];
    assign _11445 = { _11443,
                      _11444 };
    assign _11446 = _11445 < _10521;
    assign _11447 = ~ _11446;
    assign _11435 = _11101[26:26];
    assign _11432 = _11427 - _10521;
    assign _11433 = _11429 ? _11432 : _11427;
    assign _11434 = _11433[62:0];
    assign _11436 = { _11434,
                      _11435 };
    assign _11437 = _11436 < _10521;
    assign _11438 = ~ _11437;
    assign _11426 = _11101[27:27];
    assign _11423 = _11418 - _10521;
    assign _11424 = _11420 ? _11423 : _11418;
    assign _11425 = _11424[62:0];
    assign _11427 = { _11425,
                      _11426 };
    assign _11428 = _11427 < _10521;
    assign _11429 = ~ _11428;
    assign _11417 = _11101[28:28];
    assign _11414 = _11409 - _10521;
    assign _11415 = _11411 ? _11414 : _11409;
    assign _11416 = _11415[62:0];
    assign _11418 = { _11416,
                      _11417 };
    assign _11419 = _11418 < _10521;
    assign _11420 = ~ _11419;
    assign _11408 = _11101[29:29];
    assign _11405 = _11400 - _10521;
    assign _11406 = _11402 ? _11405 : _11400;
    assign _11407 = _11406[62:0];
    assign _11409 = { _11407,
                      _11408 };
    assign _11410 = _11409 < _10521;
    assign _11411 = ~ _11410;
    assign _11399 = _11101[30:30];
    assign _11396 = _11391 - _10521;
    assign _11397 = _11393 ? _11396 : _11391;
    assign _11398 = _11397[62:0];
    assign _11400 = { _11398,
                      _11399 };
    assign _11401 = _11400 < _10521;
    assign _11402 = ~ _11401;
    assign _11390 = _11101[31:31];
    assign _11387 = _11382 - _10521;
    assign _11388 = _11384 ? _11387 : _11382;
    assign _11389 = _11388[62:0];
    assign _11391 = { _11389,
                      _11390 };
    assign _11392 = _11391 < _10521;
    assign _11393 = ~ _11392;
    assign _11381 = _11101[32:32];
    assign _11378 = _11373 - _10521;
    assign _11379 = _11375 ? _11378 : _11373;
    assign _11380 = _11379[62:0];
    assign _11382 = { _11380,
                      _11381 };
    assign _11383 = _11382 < _10521;
    assign _11384 = ~ _11383;
    assign _11372 = _11101[33:33];
    assign _11369 = _11364 - _10521;
    assign _11370 = _11366 ? _11369 : _11364;
    assign _11371 = _11370[62:0];
    assign _11373 = { _11371,
                      _11372 };
    assign _11374 = _11373 < _10521;
    assign _11375 = ~ _11374;
    assign _11363 = _11101[34:34];
    assign _11360 = _11355 - _10521;
    assign _11361 = _11357 ? _11360 : _11355;
    assign _11362 = _11361[62:0];
    assign _11364 = { _11362,
                      _11363 };
    assign _11365 = _11364 < _10521;
    assign _11366 = ~ _11365;
    assign _11354 = _11101[35:35];
    assign _11351 = _11346 - _10521;
    assign _11352 = _11348 ? _11351 : _11346;
    assign _11353 = _11352[62:0];
    assign _11355 = { _11353,
                      _11354 };
    assign _11356 = _11355 < _10521;
    assign _11357 = ~ _11356;
    assign _11345 = _11101[36:36];
    assign _11342 = _11337 - _10521;
    assign _11343 = _11339 ? _11342 : _11337;
    assign _11344 = _11343[62:0];
    assign _11346 = { _11344,
                      _11345 };
    assign _11347 = _11346 < _10521;
    assign _11348 = ~ _11347;
    assign _11336 = _11101[37:37];
    assign _11333 = _11328 - _10521;
    assign _11334 = _11330 ? _11333 : _11328;
    assign _11335 = _11334[62:0];
    assign _11337 = { _11335,
                      _11336 };
    assign _11338 = _11337 < _10521;
    assign _11339 = ~ _11338;
    assign _11327 = _11101[38:38];
    assign _11324 = _11319 - _10521;
    assign _11325 = _11321 ? _11324 : _11319;
    assign _11326 = _11325[62:0];
    assign _11328 = { _11326,
                      _11327 };
    assign _11329 = _11328 < _10521;
    assign _11330 = ~ _11329;
    assign _11318 = _11101[39:39];
    assign _11315 = _11310 - _10521;
    assign _11316 = _11312 ? _11315 : _11310;
    assign _11317 = _11316[62:0];
    assign _11319 = { _11317,
                      _11318 };
    assign _11320 = _11319 < _10521;
    assign _11321 = ~ _11320;
    assign _11309 = _11101[40:40];
    assign _11306 = _11301 - _10521;
    assign _11307 = _11303 ? _11306 : _11301;
    assign _11308 = _11307[62:0];
    assign _11310 = { _11308,
                      _11309 };
    assign _11311 = _11310 < _10521;
    assign _11312 = ~ _11311;
    assign _11300 = _11101[41:41];
    assign _11297 = _11292 - _10521;
    assign _11298 = _11294 ? _11297 : _11292;
    assign _11299 = _11298[62:0];
    assign _11301 = { _11299,
                      _11300 };
    assign _11302 = _11301 < _10521;
    assign _11303 = ~ _11302;
    assign _11291 = _11101[42:42];
    assign _11288 = _11283 - _10521;
    assign _11289 = _11285 ? _11288 : _11283;
    assign _11290 = _11289[62:0];
    assign _11292 = { _11290,
                      _11291 };
    assign _11293 = _11292 < _10521;
    assign _11294 = ~ _11293;
    assign _11282 = _11101[43:43];
    assign _11279 = _11274 - _10521;
    assign _11280 = _11276 ? _11279 : _11274;
    assign _11281 = _11280[62:0];
    assign _11283 = { _11281,
                      _11282 };
    assign _11284 = _11283 < _10521;
    assign _11285 = ~ _11284;
    assign _11273 = _11101[44:44];
    assign _11270 = _11265 - _10521;
    assign _11271 = _11267 ? _11270 : _11265;
    assign _11272 = _11271[62:0];
    assign _11274 = { _11272,
                      _11273 };
    assign _11275 = _11274 < _10521;
    assign _11276 = ~ _11275;
    assign _11264 = _11101[45:45];
    assign _11261 = _11256 - _10521;
    assign _11262 = _11258 ? _11261 : _11256;
    assign _11263 = _11262[62:0];
    assign _11265 = { _11263,
                      _11264 };
    assign _11266 = _11265 < _10521;
    assign _11267 = ~ _11266;
    assign _11255 = _11101[46:46];
    assign _11252 = _11247 - _10521;
    assign _11253 = _11249 ? _11252 : _11247;
    assign _11254 = _11253[62:0];
    assign _11256 = { _11254,
                      _11255 };
    assign _11257 = _11256 < _10521;
    assign _11258 = ~ _11257;
    assign _11246 = _11101[47:47];
    assign _11243 = _11238 - _10521;
    assign _11244 = _11240 ? _11243 : _11238;
    assign _11245 = _11244[62:0];
    assign _11247 = { _11245,
                      _11246 };
    assign _11248 = _11247 < _10521;
    assign _11249 = ~ _11248;
    assign _11237 = _11101[48:48];
    assign _11234 = _11229 - _10521;
    assign _11235 = _11231 ? _11234 : _11229;
    assign _11236 = _11235[62:0];
    assign _11238 = { _11236,
                      _11237 };
    assign _11239 = _11238 < _10521;
    assign _11240 = ~ _11239;
    assign _11228 = _11101[49:49];
    assign _11225 = _11220 - _10521;
    assign _11226 = _11222 ? _11225 : _11220;
    assign _11227 = _11226[62:0];
    assign _11229 = { _11227,
                      _11228 };
    assign _11230 = _11229 < _10521;
    assign _11231 = ~ _11230;
    assign _11219 = _11101[50:50];
    assign _11216 = _11211 - _10521;
    assign _11217 = _11213 ? _11216 : _11211;
    assign _11218 = _11217[62:0];
    assign _11220 = { _11218,
                      _11219 };
    assign _11221 = _11220 < _10521;
    assign _11222 = ~ _11221;
    assign _11210 = _11101[51:51];
    assign _11207 = _11202 - _10521;
    assign _11208 = _11204 ? _11207 : _11202;
    assign _11209 = _11208[62:0];
    assign _11211 = { _11209,
                      _11210 };
    assign _11212 = _11211 < _10521;
    assign _11213 = ~ _11212;
    assign _11201 = _11101[52:52];
    assign _11198 = _11193 - _10521;
    assign _11199 = _11195 ? _11198 : _11193;
    assign _11200 = _11199[62:0];
    assign _11202 = { _11200,
                      _11201 };
    assign _11203 = _11202 < _10521;
    assign _11204 = ~ _11203;
    assign _11192 = _11101[53:53];
    assign _11189 = _11184 - _10521;
    assign _11190 = _11186 ? _11189 : _11184;
    assign _11191 = _11190[62:0];
    assign _11193 = { _11191,
                      _11192 };
    assign _11194 = _11193 < _10521;
    assign _11195 = ~ _11194;
    assign _11183 = _11101[54:54];
    assign _11180 = _11175 - _10521;
    assign _11181 = _11177 ? _11180 : _11175;
    assign _11182 = _11181[62:0];
    assign _11184 = { _11182,
                      _11183 };
    assign _11185 = _11184 < _10521;
    assign _11186 = ~ _11185;
    assign _11174 = _11101[55:55];
    assign _11171 = _11166 - _10521;
    assign _11172 = _11168 ? _11171 : _11166;
    assign _11173 = _11172[62:0];
    assign _11175 = { _11173,
                      _11174 };
    assign _11176 = _11175 < _10521;
    assign _11177 = ~ _11176;
    assign _11165 = _11101[56:56];
    assign _11162 = _11157 - _10521;
    assign _11163 = _11159 ? _11162 : _11157;
    assign _11164 = _11163[62:0];
    assign _11166 = { _11164,
                      _11165 };
    assign _11167 = _11166 < _10521;
    assign _11168 = ~ _11167;
    assign _11156 = _11101[57:57];
    assign _11153 = _11148 - _10521;
    assign _11154 = _11150 ? _11153 : _11148;
    assign _11155 = _11154[62:0];
    assign _11157 = { _11155,
                      _11156 };
    assign _11158 = _11157 < _10521;
    assign _11159 = ~ _11158;
    assign _11147 = _11101[58:58];
    assign _11144 = _11139 - _10521;
    assign _11145 = _11141 ? _11144 : _11139;
    assign _11146 = _11145[62:0];
    assign _11148 = { _11146,
                      _11147 };
    assign _11149 = _11148 < _10521;
    assign _11150 = ~ _11149;
    assign _11138 = _11101[59:59];
    assign _11135 = _11130 - _10521;
    assign _11136 = _11132 ? _11135 : _11130;
    assign _11137 = _11136[62:0];
    assign _11139 = { _11137,
                      _11138 };
    assign _11140 = _11139 < _10521;
    assign _11141 = ~ _11140;
    assign _11129 = _11101[60:60];
    assign _11126 = _11121 - _10521;
    assign _11127 = _11123 ? _11126 : _11121;
    assign _11128 = _11127[62:0];
    assign _11130 = { _11128,
                      _11129 };
    assign _11131 = _11130 < _10521;
    assign _11132 = ~ _11131;
    assign _11120 = _11101[61:61];
    assign _11117 = _11112 - _10521;
    assign _11118 = _11114 ? _11117 : _11112;
    assign _11119 = _11118[62:0];
    assign _11121 = { _11119,
                      _11120 };
    assign _11122 = _11121 < _10521;
    assign _11123 = ~ _11122;
    assign _11111 = _11101[62:62];
    assign _11108 = _11103 - _10521;
    assign _11109 = _11105 ? _11108 : _11103;
    assign _11110 = _11109[62:0];
    assign _11112 = { _11110,
                      _11111 };
    assign _11113 = _11112 < _10521;
    assign _11114 = ~ _11113;
    assign _11101 = _10513 - _11095;
    assign _11102 = _11101[63:63];
    assign _11103 = { _22185,
                      _11102 };
    assign _11104 = _11103 < _10521;
    assign _11105 = ~ _11104;
    assign _11106 = { _22185,
                      _11105 };
    assign _11107 = _11106[62:0];
    assign _11115 = { _11107,
                      _11114 };
    assign _11116 = _11115[62:0];
    assign _11124 = { _11116,
                      _11123 };
    assign _11125 = _11124[62:0];
    assign _11133 = { _11125,
                      _11132 };
    assign _11134 = _11133[62:0];
    assign _11142 = { _11134,
                      _11141 };
    assign _11143 = _11142[62:0];
    assign _11151 = { _11143,
                      _11150 };
    assign _11152 = _11151[62:0];
    assign _11160 = { _11152,
                      _11159 };
    assign _11161 = _11160[62:0];
    assign _11169 = { _11161,
                      _11168 };
    assign _11170 = _11169[62:0];
    assign _11178 = { _11170,
                      _11177 };
    assign _11179 = _11178[62:0];
    assign _11187 = { _11179,
                      _11186 };
    assign _11188 = _11187[62:0];
    assign _11196 = { _11188,
                      _11195 };
    assign _11197 = _11196[62:0];
    assign _11205 = { _11197,
                      _11204 };
    assign _11206 = _11205[62:0];
    assign _11214 = { _11206,
                      _11213 };
    assign _11215 = _11214[62:0];
    assign _11223 = { _11215,
                      _11222 };
    assign _11224 = _11223[62:0];
    assign _11232 = { _11224,
                      _11231 };
    assign _11233 = _11232[62:0];
    assign _11241 = { _11233,
                      _11240 };
    assign _11242 = _11241[62:0];
    assign _11250 = { _11242,
                      _11249 };
    assign _11251 = _11250[62:0];
    assign _11259 = { _11251,
                      _11258 };
    assign _11260 = _11259[62:0];
    assign _11268 = { _11260,
                      _11267 };
    assign _11269 = _11268[62:0];
    assign _11277 = { _11269,
                      _11276 };
    assign _11278 = _11277[62:0];
    assign _11286 = { _11278,
                      _11285 };
    assign _11287 = _11286[62:0];
    assign _11295 = { _11287,
                      _11294 };
    assign _11296 = _11295[62:0];
    assign _11304 = { _11296,
                      _11303 };
    assign _11305 = _11304[62:0];
    assign _11313 = { _11305,
                      _11312 };
    assign _11314 = _11313[62:0];
    assign _11322 = { _11314,
                      _11321 };
    assign _11323 = _11322[62:0];
    assign _11331 = { _11323,
                      _11330 };
    assign _11332 = _11331[62:0];
    assign _11340 = { _11332,
                      _11339 };
    assign _11341 = _11340[62:0];
    assign _11349 = { _11341,
                      _11348 };
    assign _11350 = _11349[62:0];
    assign _11358 = { _11350,
                      _11357 };
    assign _11359 = _11358[62:0];
    assign _11367 = { _11359,
                      _11366 };
    assign _11368 = _11367[62:0];
    assign _11376 = { _11368,
                      _11375 };
    assign _11377 = _11376[62:0];
    assign _11385 = { _11377,
                      _11384 };
    assign _11386 = _11385[62:0];
    assign _11394 = { _11386,
                      _11393 };
    assign _11395 = _11394[62:0];
    assign _11403 = { _11395,
                      _11402 };
    assign _11404 = _11403[62:0];
    assign _11412 = { _11404,
                      _11411 };
    assign _11413 = _11412[62:0];
    assign _11421 = { _11413,
                      _11420 };
    assign _11422 = _11421[62:0];
    assign _11430 = { _11422,
                      _11429 };
    assign _11431 = _11430[62:0];
    assign _11439 = { _11431,
                      _11438 };
    assign _11440 = _11439[62:0];
    assign _11448 = { _11440,
                      _11447 };
    assign _11449 = _11448[62:0];
    assign _11457 = { _11449,
                      _11456 };
    assign _11458 = _11457[62:0];
    assign _11466 = { _11458,
                      _11465 };
    assign _11467 = _11466[62:0];
    assign _11475 = { _11467,
                      _11474 };
    assign _11476 = _11475[62:0];
    assign _11484 = { _11476,
                      _11483 };
    assign _11485 = _11484[62:0];
    assign _11493 = { _11485,
                      _11492 };
    assign _11494 = _11493[62:0];
    assign _11502 = { _11494,
                      _11501 };
    assign _11503 = _11502[62:0];
    assign _11511 = { _11503,
                      _11510 };
    assign _11512 = _11511[62:0];
    assign _11520 = { _11512,
                      _11519 };
    assign _11521 = _11520[62:0];
    assign _11529 = { _11521,
                      _11528 };
    assign _11530 = _11529[62:0];
    assign _11538 = { _11530,
                      _11537 };
    assign _11539 = _11538[62:0];
    assign _11547 = { _11539,
                      _11546 };
    assign _11548 = _11547[62:0];
    assign _11556 = { _11548,
                      _11555 };
    assign _11557 = _11556[62:0];
    assign _11565 = { _11557,
                      _11564 };
    assign _11566 = _11565[62:0];
    assign _11574 = { _11566,
                      _11573 };
    assign _11575 = _11574[62:0];
    assign _11583 = { _11575,
                      _11582 };
    assign _11584 = _11583[62:0];
    assign _11592 = { _11584,
                      _11591 };
    assign _11593 = _11592[62:0];
    assign _11601 = { _11593,
                      _11600 };
    assign _11602 = _11601[62:0];
    assign _11610 = { _11602,
                      _11609 };
    assign _11611 = _11610[62:0];
    assign _11619 = { _11611,
                      _11618 };
    assign _11620 = _11619[62:0];
    assign _11628 = { _11620,
                      _11627 };
    assign _11629 = _11628[62:0];
    assign _11637 = { _11629,
                      _11636 };
    assign _11638 = _11637[62:0];
    assign _11646 = { _11638,
                      _11645 };
    assign _11647 = _11646[62:0];
    assign _11655 = { _11647,
                      _11654 };
    assign _11656 = _11655[62:0];
    assign _11664 = { _11656,
                      _11663 };
    assign _11665 = _11664[62:0];
    assign _11673 = { _11665,
                      _11672 };
    assign _11675 = _11673 + _22186;
    assign _11676 = _11675 * _11095;
    assign _11677 = _11676[63:0];
    assign _12259 = _11677 + _12258;
    assign _11087 = _10518[0:0];
    assign _11084 = _11079 - _10521;
    assign _11085 = _11081 ? _11084 : _11079;
    assign _11086 = _11085[62:0];
    assign _11088 = { _11086,
                      _11087 };
    assign _11089 = _11088 < _10521;
    assign _11090 = ~ _11089;
    assign _11078 = _10518[1:1];
    assign _11075 = _11070 - _10521;
    assign _11076 = _11072 ? _11075 : _11070;
    assign _11077 = _11076[62:0];
    assign _11079 = { _11077,
                      _11078 };
    assign _11080 = _11079 < _10521;
    assign _11081 = ~ _11080;
    assign _11069 = _10518[2:2];
    assign _11066 = _11061 - _10521;
    assign _11067 = _11063 ? _11066 : _11061;
    assign _11068 = _11067[62:0];
    assign _11070 = { _11068,
                      _11069 };
    assign _11071 = _11070 < _10521;
    assign _11072 = ~ _11071;
    assign _11060 = _10518[3:3];
    assign _11057 = _11052 - _10521;
    assign _11058 = _11054 ? _11057 : _11052;
    assign _11059 = _11058[62:0];
    assign _11061 = { _11059,
                      _11060 };
    assign _11062 = _11061 < _10521;
    assign _11063 = ~ _11062;
    assign _11051 = _10518[4:4];
    assign _11048 = _11043 - _10521;
    assign _11049 = _11045 ? _11048 : _11043;
    assign _11050 = _11049[62:0];
    assign _11052 = { _11050,
                      _11051 };
    assign _11053 = _11052 < _10521;
    assign _11054 = ~ _11053;
    assign _11042 = _10518[5:5];
    assign _11039 = _11034 - _10521;
    assign _11040 = _11036 ? _11039 : _11034;
    assign _11041 = _11040[62:0];
    assign _11043 = { _11041,
                      _11042 };
    assign _11044 = _11043 < _10521;
    assign _11045 = ~ _11044;
    assign _11033 = _10518[6:6];
    assign _11030 = _11025 - _10521;
    assign _11031 = _11027 ? _11030 : _11025;
    assign _11032 = _11031[62:0];
    assign _11034 = { _11032,
                      _11033 };
    assign _11035 = _11034 < _10521;
    assign _11036 = ~ _11035;
    assign _11024 = _10518[7:7];
    assign _11021 = _11016 - _10521;
    assign _11022 = _11018 ? _11021 : _11016;
    assign _11023 = _11022[62:0];
    assign _11025 = { _11023,
                      _11024 };
    assign _11026 = _11025 < _10521;
    assign _11027 = ~ _11026;
    assign _11015 = _10518[8:8];
    assign _11012 = _11007 - _10521;
    assign _11013 = _11009 ? _11012 : _11007;
    assign _11014 = _11013[62:0];
    assign _11016 = { _11014,
                      _11015 };
    assign _11017 = _11016 < _10521;
    assign _11018 = ~ _11017;
    assign _11006 = _10518[9:9];
    assign _11003 = _10998 - _10521;
    assign _11004 = _11000 ? _11003 : _10998;
    assign _11005 = _11004[62:0];
    assign _11007 = { _11005,
                      _11006 };
    assign _11008 = _11007 < _10521;
    assign _11009 = ~ _11008;
    assign _10997 = _10518[10:10];
    assign _10994 = _10989 - _10521;
    assign _10995 = _10991 ? _10994 : _10989;
    assign _10996 = _10995[62:0];
    assign _10998 = { _10996,
                      _10997 };
    assign _10999 = _10998 < _10521;
    assign _11000 = ~ _10999;
    assign _10988 = _10518[11:11];
    assign _10985 = _10980 - _10521;
    assign _10986 = _10982 ? _10985 : _10980;
    assign _10987 = _10986[62:0];
    assign _10989 = { _10987,
                      _10988 };
    assign _10990 = _10989 < _10521;
    assign _10991 = ~ _10990;
    assign _10979 = _10518[12:12];
    assign _10976 = _10971 - _10521;
    assign _10977 = _10973 ? _10976 : _10971;
    assign _10978 = _10977[62:0];
    assign _10980 = { _10978,
                      _10979 };
    assign _10981 = _10980 < _10521;
    assign _10982 = ~ _10981;
    assign _10970 = _10518[13:13];
    assign _10967 = _10962 - _10521;
    assign _10968 = _10964 ? _10967 : _10962;
    assign _10969 = _10968[62:0];
    assign _10971 = { _10969,
                      _10970 };
    assign _10972 = _10971 < _10521;
    assign _10973 = ~ _10972;
    assign _10961 = _10518[14:14];
    assign _10958 = _10953 - _10521;
    assign _10959 = _10955 ? _10958 : _10953;
    assign _10960 = _10959[62:0];
    assign _10962 = { _10960,
                      _10961 };
    assign _10963 = _10962 < _10521;
    assign _10964 = ~ _10963;
    assign _10952 = _10518[15:15];
    assign _10949 = _10944 - _10521;
    assign _10950 = _10946 ? _10949 : _10944;
    assign _10951 = _10950[62:0];
    assign _10953 = { _10951,
                      _10952 };
    assign _10954 = _10953 < _10521;
    assign _10955 = ~ _10954;
    assign _10943 = _10518[16:16];
    assign _10940 = _10935 - _10521;
    assign _10941 = _10937 ? _10940 : _10935;
    assign _10942 = _10941[62:0];
    assign _10944 = { _10942,
                      _10943 };
    assign _10945 = _10944 < _10521;
    assign _10946 = ~ _10945;
    assign _10934 = _10518[17:17];
    assign _10931 = _10926 - _10521;
    assign _10932 = _10928 ? _10931 : _10926;
    assign _10933 = _10932[62:0];
    assign _10935 = { _10933,
                      _10934 };
    assign _10936 = _10935 < _10521;
    assign _10937 = ~ _10936;
    assign _10925 = _10518[18:18];
    assign _10922 = _10917 - _10521;
    assign _10923 = _10919 ? _10922 : _10917;
    assign _10924 = _10923[62:0];
    assign _10926 = { _10924,
                      _10925 };
    assign _10927 = _10926 < _10521;
    assign _10928 = ~ _10927;
    assign _10916 = _10518[19:19];
    assign _10913 = _10908 - _10521;
    assign _10914 = _10910 ? _10913 : _10908;
    assign _10915 = _10914[62:0];
    assign _10917 = { _10915,
                      _10916 };
    assign _10918 = _10917 < _10521;
    assign _10919 = ~ _10918;
    assign _10907 = _10518[20:20];
    assign _10904 = _10899 - _10521;
    assign _10905 = _10901 ? _10904 : _10899;
    assign _10906 = _10905[62:0];
    assign _10908 = { _10906,
                      _10907 };
    assign _10909 = _10908 < _10521;
    assign _10910 = ~ _10909;
    assign _10898 = _10518[21:21];
    assign _10895 = _10890 - _10521;
    assign _10896 = _10892 ? _10895 : _10890;
    assign _10897 = _10896[62:0];
    assign _10899 = { _10897,
                      _10898 };
    assign _10900 = _10899 < _10521;
    assign _10901 = ~ _10900;
    assign _10889 = _10518[22:22];
    assign _10886 = _10881 - _10521;
    assign _10887 = _10883 ? _10886 : _10881;
    assign _10888 = _10887[62:0];
    assign _10890 = { _10888,
                      _10889 };
    assign _10891 = _10890 < _10521;
    assign _10892 = ~ _10891;
    assign _10880 = _10518[23:23];
    assign _10877 = _10872 - _10521;
    assign _10878 = _10874 ? _10877 : _10872;
    assign _10879 = _10878[62:0];
    assign _10881 = { _10879,
                      _10880 };
    assign _10882 = _10881 < _10521;
    assign _10883 = ~ _10882;
    assign _10871 = _10518[24:24];
    assign _10868 = _10863 - _10521;
    assign _10869 = _10865 ? _10868 : _10863;
    assign _10870 = _10869[62:0];
    assign _10872 = { _10870,
                      _10871 };
    assign _10873 = _10872 < _10521;
    assign _10874 = ~ _10873;
    assign _10862 = _10518[25:25];
    assign _10859 = _10854 - _10521;
    assign _10860 = _10856 ? _10859 : _10854;
    assign _10861 = _10860[62:0];
    assign _10863 = { _10861,
                      _10862 };
    assign _10864 = _10863 < _10521;
    assign _10865 = ~ _10864;
    assign _10853 = _10518[26:26];
    assign _10850 = _10845 - _10521;
    assign _10851 = _10847 ? _10850 : _10845;
    assign _10852 = _10851[62:0];
    assign _10854 = { _10852,
                      _10853 };
    assign _10855 = _10854 < _10521;
    assign _10856 = ~ _10855;
    assign _10844 = _10518[27:27];
    assign _10841 = _10836 - _10521;
    assign _10842 = _10838 ? _10841 : _10836;
    assign _10843 = _10842[62:0];
    assign _10845 = { _10843,
                      _10844 };
    assign _10846 = _10845 < _10521;
    assign _10847 = ~ _10846;
    assign _10835 = _10518[28:28];
    assign _10832 = _10827 - _10521;
    assign _10833 = _10829 ? _10832 : _10827;
    assign _10834 = _10833[62:0];
    assign _10836 = { _10834,
                      _10835 };
    assign _10837 = _10836 < _10521;
    assign _10838 = ~ _10837;
    assign _10826 = _10518[29:29];
    assign _10823 = _10818 - _10521;
    assign _10824 = _10820 ? _10823 : _10818;
    assign _10825 = _10824[62:0];
    assign _10827 = { _10825,
                      _10826 };
    assign _10828 = _10827 < _10521;
    assign _10829 = ~ _10828;
    assign _10817 = _10518[30:30];
    assign _10814 = _10809 - _10521;
    assign _10815 = _10811 ? _10814 : _10809;
    assign _10816 = _10815[62:0];
    assign _10818 = { _10816,
                      _10817 };
    assign _10819 = _10818 < _10521;
    assign _10820 = ~ _10819;
    assign _10808 = _10518[31:31];
    assign _10805 = _10800 - _10521;
    assign _10806 = _10802 ? _10805 : _10800;
    assign _10807 = _10806[62:0];
    assign _10809 = { _10807,
                      _10808 };
    assign _10810 = _10809 < _10521;
    assign _10811 = ~ _10810;
    assign _10799 = _10518[32:32];
    assign _10796 = _10791 - _10521;
    assign _10797 = _10793 ? _10796 : _10791;
    assign _10798 = _10797[62:0];
    assign _10800 = { _10798,
                      _10799 };
    assign _10801 = _10800 < _10521;
    assign _10802 = ~ _10801;
    assign _10790 = _10518[33:33];
    assign _10787 = _10782 - _10521;
    assign _10788 = _10784 ? _10787 : _10782;
    assign _10789 = _10788[62:0];
    assign _10791 = { _10789,
                      _10790 };
    assign _10792 = _10791 < _10521;
    assign _10793 = ~ _10792;
    assign _10781 = _10518[34:34];
    assign _10778 = _10773 - _10521;
    assign _10779 = _10775 ? _10778 : _10773;
    assign _10780 = _10779[62:0];
    assign _10782 = { _10780,
                      _10781 };
    assign _10783 = _10782 < _10521;
    assign _10784 = ~ _10783;
    assign _10772 = _10518[35:35];
    assign _10769 = _10764 - _10521;
    assign _10770 = _10766 ? _10769 : _10764;
    assign _10771 = _10770[62:0];
    assign _10773 = { _10771,
                      _10772 };
    assign _10774 = _10773 < _10521;
    assign _10775 = ~ _10774;
    assign _10763 = _10518[36:36];
    assign _10760 = _10755 - _10521;
    assign _10761 = _10757 ? _10760 : _10755;
    assign _10762 = _10761[62:0];
    assign _10764 = { _10762,
                      _10763 };
    assign _10765 = _10764 < _10521;
    assign _10766 = ~ _10765;
    assign _10754 = _10518[37:37];
    assign _10751 = _10746 - _10521;
    assign _10752 = _10748 ? _10751 : _10746;
    assign _10753 = _10752[62:0];
    assign _10755 = { _10753,
                      _10754 };
    assign _10756 = _10755 < _10521;
    assign _10757 = ~ _10756;
    assign _10745 = _10518[38:38];
    assign _10742 = _10737 - _10521;
    assign _10743 = _10739 ? _10742 : _10737;
    assign _10744 = _10743[62:0];
    assign _10746 = { _10744,
                      _10745 };
    assign _10747 = _10746 < _10521;
    assign _10748 = ~ _10747;
    assign _10736 = _10518[39:39];
    assign _10733 = _10728 - _10521;
    assign _10734 = _10730 ? _10733 : _10728;
    assign _10735 = _10734[62:0];
    assign _10737 = { _10735,
                      _10736 };
    assign _10738 = _10737 < _10521;
    assign _10739 = ~ _10738;
    assign _10727 = _10518[40:40];
    assign _10724 = _10719 - _10521;
    assign _10725 = _10721 ? _10724 : _10719;
    assign _10726 = _10725[62:0];
    assign _10728 = { _10726,
                      _10727 };
    assign _10729 = _10728 < _10521;
    assign _10730 = ~ _10729;
    assign _10718 = _10518[41:41];
    assign _10715 = _10710 - _10521;
    assign _10716 = _10712 ? _10715 : _10710;
    assign _10717 = _10716[62:0];
    assign _10719 = { _10717,
                      _10718 };
    assign _10720 = _10719 < _10521;
    assign _10721 = ~ _10720;
    assign _10709 = _10518[42:42];
    assign _10706 = _10701 - _10521;
    assign _10707 = _10703 ? _10706 : _10701;
    assign _10708 = _10707[62:0];
    assign _10710 = { _10708,
                      _10709 };
    assign _10711 = _10710 < _10521;
    assign _10712 = ~ _10711;
    assign _10700 = _10518[43:43];
    assign _10697 = _10692 - _10521;
    assign _10698 = _10694 ? _10697 : _10692;
    assign _10699 = _10698[62:0];
    assign _10701 = { _10699,
                      _10700 };
    assign _10702 = _10701 < _10521;
    assign _10703 = ~ _10702;
    assign _10691 = _10518[44:44];
    assign _10688 = _10683 - _10521;
    assign _10689 = _10685 ? _10688 : _10683;
    assign _10690 = _10689[62:0];
    assign _10692 = { _10690,
                      _10691 };
    assign _10693 = _10692 < _10521;
    assign _10694 = ~ _10693;
    assign _10682 = _10518[45:45];
    assign _10679 = _10674 - _10521;
    assign _10680 = _10676 ? _10679 : _10674;
    assign _10681 = _10680[62:0];
    assign _10683 = { _10681,
                      _10682 };
    assign _10684 = _10683 < _10521;
    assign _10685 = ~ _10684;
    assign _10673 = _10518[46:46];
    assign _10670 = _10665 - _10521;
    assign _10671 = _10667 ? _10670 : _10665;
    assign _10672 = _10671[62:0];
    assign _10674 = { _10672,
                      _10673 };
    assign _10675 = _10674 < _10521;
    assign _10676 = ~ _10675;
    assign _10664 = _10518[47:47];
    assign _10661 = _10656 - _10521;
    assign _10662 = _10658 ? _10661 : _10656;
    assign _10663 = _10662[62:0];
    assign _10665 = { _10663,
                      _10664 };
    assign _10666 = _10665 < _10521;
    assign _10667 = ~ _10666;
    assign _10655 = _10518[48:48];
    assign _10652 = _10647 - _10521;
    assign _10653 = _10649 ? _10652 : _10647;
    assign _10654 = _10653[62:0];
    assign _10656 = { _10654,
                      _10655 };
    assign _10657 = _10656 < _10521;
    assign _10658 = ~ _10657;
    assign _10646 = _10518[49:49];
    assign _10643 = _10638 - _10521;
    assign _10644 = _10640 ? _10643 : _10638;
    assign _10645 = _10644[62:0];
    assign _10647 = { _10645,
                      _10646 };
    assign _10648 = _10647 < _10521;
    assign _10649 = ~ _10648;
    assign _10637 = _10518[50:50];
    assign _10634 = _10629 - _10521;
    assign _10635 = _10631 ? _10634 : _10629;
    assign _10636 = _10635[62:0];
    assign _10638 = { _10636,
                      _10637 };
    assign _10639 = _10638 < _10521;
    assign _10640 = ~ _10639;
    assign _10628 = _10518[51:51];
    assign _10625 = _10620 - _10521;
    assign _10626 = _10622 ? _10625 : _10620;
    assign _10627 = _10626[62:0];
    assign _10629 = { _10627,
                      _10628 };
    assign _10630 = _10629 < _10521;
    assign _10631 = ~ _10630;
    assign _10619 = _10518[52:52];
    assign _10616 = _10611 - _10521;
    assign _10617 = _10613 ? _10616 : _10611;
    assign _10618 = _10617[62:0];
    assign _10620 = { _10618,
                      _10619 };
    assign _10621 = _10620 < _10521;
    assign _10622 = ~ _10621;
    assign _10610 = _10518[53:53];
    assign _10607 = _10602 - _10521;
    assign _10608 = _10604 ? _10607 : _10602;
    assign _10609 = _10608[62:0];
    assign _10611 = { _10609,
                      _10610 };
    assign _10612 = _10611 < _10521;
    assign _10613 = ~ _10612;
    assign _10601 = _10518[54:54];
    assign _10598 = _10593 - _10521;
    assign _10599 = _10595 ? _10598 : _10593;
    assign _10600 = _10599[62:0];
    assign _10602 = { _10600,
                      _10601 };
    assign _10603 = _10602 < _10521;
    assign _10604 = ~ _10603;
    assign _10592 = _10518[55:55];
    assign _10589 = _10584 - _10521;
    assign _10590 = _10586 ? _10589 : _10584;
    assign _10591 = _10590[62:0];
    assign _10593 = { _10591,
                      _10592 };
    assign _10594 = _10593 < _10521;
    assign _10595 = ~ _10594;
    assign _10583 = _10518[56:56];
    assign _10580 = _10575 - _10521;
    assign _10581 = _10577 ? _10580 : _10575;
    assign _10582 = _10581[62:0];
    assign _10584 = { _10582,
                      _10583 };
    assign _10585 = _10584 < _10521;
    assign _10586 = ~ _10585;
    assign _10574 = _10518[57:57];
    assign _10571 = _10566 - _10521;
    assign _10572 = _10568 ? _10571 : _10566;
    assign _10573 = _10572[62:0];
    assign _10575 = { _10573,
                      _10574 };
    assign _10576 = _10575 < _10521;
    assign _10577 = ~ _10576;
    assign _10565 = _10518[58:58];
    assign _10562 = _10557 - _10521;
    assign _10563 = _10559 ? _10562 : _10557;
    assign _10564 = _10563[62:0];
    assign _10566 = { _10564,
                      _10565 };
    assign _10567 = _10566 < _10521;
    assign _10568 = ~ _10567;
    assign _10556 = _10518[59:59];
    assign _10553 = _10548 - _10521;
    assign _10554 = _10550 ? _10553 : _10548;
    assign _10555 = _10554[62:0];
    assign _10557 = { _10555,
                      _10556 };
    assign _10558 = _10557 < _10521;
    assign _10559 = ~ _10558;
    assign _10547 = _10518[60:60];
    assign _10544 = _10539 - _10521;
    assign _10545 = _10541 ? _10544 : _10539;
    assign _10546 = _10545[62:0];
    assign _10548 = { _10546,
                      _10547 };
    assign _10549 = _10548 < _10521;
    assign _10550 = ~ _10549;
    assign _10538 = _10518[61:61];
    assign _10535 = _10530 - _10521;
    assign _10536 = _10532 ? _10535 : _10530;
    assign _10537 = _10536[62:0];
    assign _10539 = { _10537,
                      _10538 };
    assign _10540 = _10539 < _10521;
    assign _10541 = ~ _10540;
    assign _10529 = _10518[62:62];
    assign _10526 = _10520 - _10521;
    assign _10527 = _10523 ? _10526 : _10520;
    assign _10528 = _10527[62:0];
    assign _10530 = { _10528,
                      _10529 };
    assign _10531 = _10530 < _10521;
    assign _10532 = ~ _10531;
    assign _10521 = 64'b0000000000000000000000000000000000000000000000000010101101100111;
    assign _10517 = 64'b0000000000000000000000000000000000000000000000000010101101100110;
    assign _10518 = _3 + _10517;
    assign _10519 = _10518[63:63];
    assign _10520 = { _22185,
                      _10519 };
    assign _10522 = _10520 < _10521;
    assign _10523 = ~ _10522;
    assign _10524 = { _22185,
                      _10523 };
    assign _10525 = _10524[62:0];
    assign _10533 = { _10525,
                      _10532 };
    assign _10534 = _10533[62:0];
    assign _10542 = { _10534,
                      _10541 };
    assign _10543 = _10542[62:0];
    assign _10551 = { _10543,
                      _10550 };
    assign _10552 = _10551[62:0];
    assign _10560 = { _10552,
                      _10559 };
    assign _10561 = _10560[62:0];
    assign _10569 = { _10561,
                      _10568 };
    assign _10570 = _10569[62:0];
    assign _10578 = { _10570,
                      _10577 };
    assign _10579 = _10578[62:0];
    assign _10587 = { _10579,
                      _10586 };
    assign _10588 = _10587[62:0];
    assign _10596 = { _10588,
                      _10595 };
    assign _10597 = _10596[62:0];
    assign _10605 = { _10597,
                      _10604 };
    assign _10606 = _10605[62:0];
    assign _10614 = { _10606,
                      _10613 };
    assign _10615 = _10614[62:0];
    assign _10623 = { _10615,
                      _10622 };
    assign _10624 = _10623[62:0];
    assign _10632 = { _10624,
                      _10631 };
    assign _10633 = _10632[62:0];
    assign _10641 = { _10633,
                      _10640 };
    assign _10642 = _10641[62:0];
    assign _10650 = { _10642,
                      _10649 };
    assign _10651 = _10650[62:0];
    assign _10659 = { _10651,
                      _10658 };
    assign _10660 = _10659[62:0];
    assign _10668 = { _10660,
                      _10667 };
    assign _10669 = _10668[62:0];
    assign _10677 = { _10669,
                      _10676 };
    assign _10678 = _10677[62:0];
    assign _10686 = { _10678,
                      _10685 };
    assign _10687 = _10686[62:0];
    assign _10695 = { _10687,
                      _10694 };
    assign _10696 = _10695[62:0];
    assign _10704 = { _10696,
                      _10703 };
    assign _10705 = _10704[62:0];
    assign _10713 = { _10705,
                      _10712 };
    assign _10714 = _10713[62:0];
    assign _10722 = { _10714,
                      _10721 };
    assign _10723 = _10722[62:0];
    assign _10731 = { _10723,
                      _10730 };
    assign _10732 = _10731[62:0];
    assign _10740 = { _10732,
                      _10739 };
    assign _10741 = _10740[62:0];
    assign _10749 = { _10741,
                      _10748 };
    assign _10750 = _10749[62:0];
    assign _10758 = { _10750,
                      _10757 };
    assign _10759 = _10758[62:0];
    assign _10767 = { _10759,
                      _10766 };
    assign _10768 = _10767[62:0];
    assign _10776 = { _10768,
                      _10775 };
    assign _10777 = _10776[62:0];
    assign _10785 = { _10777,
                      _10784 };
    assign _10786 = _10785[62:0];
    assign _10794 = { _10786,
                      _10793 };
    assign _10795 = _10794[62:0];
    assign _10803 = { _10795,
                      _10802 };
    assign _10804 = _10803[62:0];
    assign _10812 = { _10804,
                      _10811 };
    assign _10813 = _10812[62:0];
    assign _10821 = { _10813,
                      _10820 };
    assign _10822 = _10821[62:0];
    assign _10830 = { _10822,
                      _10829 };
    assign _10831 = _10830[62:0];
    assign _10839 = { _10831,
                      _10838 };
    assign _10840 = _10839[62:0];
    assign _10848 = { _10840,
                      _10847 };
    assign _10849 = _10848[62:0];
    assign _10857 = { _10849,
                      _10856 };
    assign _10858 = _10857[62:0];
    assign _10866 = { _10858,
                      _10865 };
    assign _10867 = _10866[62:0];
    assign _10875 = { _10867,
                      _10874 };
    assign _10876 = _10875[62:0];
    assign _10884 = { _10876,
                      _10883 };
    assign _10885 = _10884[62:0];
    assign _10893 = { _10885,
                      _10892 };
    assign _10894 = _10893[62:0];
    assign _10902 = { _10894,
                      _10901 };
    assign _10903 = _10902[62:0];
    assign _10911 = { _10903,
                      _10910 };
    assign _10912 = _10911[62:0];
    assign _10920 = { _10912,
                      _10919 };
    assign _10921 = _10920[62:0];
    assign _10929 = { _10921,
                      _10928 };
    assign _10930 = _10929[62:0];
    assign _10938 = { _10930,
                      _10937 };
    assign _10939 = _10938[62:0];
    assign _10947 = { _10939,
                      _10946 };
    assign _10948 = _10947[62:0];
    assign _10956 = { _10948,
                      _10955 };
    assign _10957 = _10956[62:0];
    assign _10965 = { _10957,
                      _10964 };
    assign _10966 = _10965[62:0];
    assign _10974 = { _10966,
                      _10973 };
    assign _10975 = _10974[62:0];
    assign _10983 = { _10975,
                      _10982 };
    assign _10984 = _10983[62:0];
    assign _10992 = { _10984,
                      _10991 };
    assign _10993 = _10992[62:0];
    assign _11001 = { _10993,
                      _11000 };
    assign _11002 = _11001[62:0];
    assign _11010 = { _11002,
                      _11009 };
    assign _11011 = _11010[62:0];
    assign _11019 = { _11011,
                      _11018 };
    assign _11020 = _11019[62:0];
    assign _11028 = { _11020,
                      _11027 };
    assign _11029 = _11028[62:0];
    assign _11037 = { _11029,
                      _11036 };
    assign _11038 = _11037[62:0];
    assign _11046 = { _11038,
                      _11045 };
    assign _11047 = _11046[62:0];
    assign _11055 = { _11047,
                      _11054 };
    assign _11056 = _11055[62:0];
    assign _11064 = { _11056,
                      _11063 };
    assign _11065 = _11064[62:0];
    assign _11073 = { _11065,
                      _11072 };
    assign _11074 = _11073[62:0];
    assign _11082 = { _11074,
                      _11081 };
    assign _11083 = _11082[62:0];
    assign _11091 = { _11083,
                      _11090 };
    assign _11092 = _11091 * _10521;
    assign _11093 = _11092[63:0];
    assign _11094 = _10521 < _11093;
    assign _11095 = _11094 ? _11093 : _10521;
    assign _10511 = 64'b0000000000000000000000000000000000000000000000011000011010011111;
    assign _10512 = _5 < _10511;
    assign _10513 = _10512 ? _5 : _10511;
    assign _11096 = _10513 < _11095;
    assign _11097 = ~ _11096;
    assign _12260 = _11097 ? _12259 : _21604;
    assign _10502 = _9933[0:0];
    assign _10499 = _10494 - _22192;
    assign _10500 = _10496 ? _10499 : _10494;
    assign _10501 = _10500[62:0];
    assign _10503 = { _10501,
                      _10502 };
    assign _10504 = _10503 < _22192;
    assign _10505 = ~ _10504;
    assign _10493 = _9933[1:1];
    assign _10490 = _10485 - _22192;
    assign _10491 = _10487 ? _10490 : _10485;
    assign _10492 = _10491[62:0];
    assign _10494 = { _10492,
                      _10493 };
    assign _10495 = _10494 < _22192;
    assign _10496 = ~ _10495;
    assign _10484 = _9933[2:2];
    assign _10481 = _10476 - _22192;
    assign _10482 = _10478 ? _10481 : _10476;
    assign _10483 = _10482[62:0];
    assign _10485 = { _10483,
                      _10484 };
    assign _10486 = _10485 < _22192;
    assign _10487 = ~ _10486;
    assign _10475 = _9933[3:3];
    assign _10472 = _10467 - _22192;
    assign _10473 = _10469 ? _10472 : _10467;
    assign _10474 = _10473[62:0];
    assign _10476 = { _10474,
                      _10475 };
    assign _10477 = _10476 < _22192;
    assign _10478 = ~ _10477;
    assign _10466 = _9933[4:4];
    assign _10463 = _10458 - _22192;
    assign _10464 = _10460 ? _10463 : _10458;
    assign _10465 = _10464[62:0];
    assign _10467 = { _10465,
                      _10466 };
    assign _10468 = _10467 < _22192;
    assign _10469 = ~ _10468;
    assign _10457 = _9933[5:5];
    assign _10454 = _10449 - _22192;
    assign _10455 = _10451 ? _10454 : _10449;
    assign _10456 = _10455[62:0];
    assign _10458 = { _10456,
                      _10457 };
    assign _10459 = _10458 < _22192;
    assign _10460 = ~ _10459;
    assign _10448 = _9933[6:6];
    assign _10445 = _10440 - _22192;
    assign _10446 = _10442 ? _10445 : _10440;
    assign _10447 = _10446[62:0];
    assign _10449 = { _10447,
                      _10448 };
    assign _10450 = _10449 < _22192;
    assign _10451 = ~ _10450;
    assign _10439 = _9933[7:7];
    assign _10436 = _10431 - _22192;
    assign _10437 = _10433 ? _10436 : _10431;
    assign _10438 = _10437[62:0];
    assign _10440 = { _10438,
                      _10439 };
    assign _10441 = _10440 < _22192;
    assign _10442 = ~ _10441;
    assign _10430 = _9933[8:8];
    assign _10427 = _10422 - _22192;
    assign _10428 = _10424 ? _10427 : _10422;
    assign _10429 = _10428[62:0];
    assign _10431 = { _10429,
                      _10430 };
    assign _10432 = _10431 < _22192;
    assign _10433 = ~ _10432;
    assign _10421 = _9933[9:9];
    assign _10418 = _10413 - _22192;
    assign _10419 = _10415 ? _10418 : _10413;
    assign _10420 = _10419[62:0];
    assign _10422 = { _10420,
                      _10421 };
    assign _10423 = _10422 < _22192;
    assign _10424 = ~ _10423;
    assign _10412 = _9933[10:10];
    assign _10409 = _10404 - _22192;
    assign _10410 = _10406 ? _10409 : _10404;
    assign _10411 = _10410[62:0];
    assign _10413 = { _10411,
                      _10412 };
    assign _10414 = _10413 < _22192;
    assign _10415 = ~ _10414;
    assign _10403 = _9933[11:11];
    assign _10400 = _10395 - _22192;
    assign _10401 = _10397 ? _10400 : _10395;
    assign _10402 = _10401[62:0];
    assign _10404 = { _10402,
                      _10403 };
    assign _10405 = _10404 < _22192;
    assign _10406 = ~ _10405;
    assign _10394 = _9933[12:12];
    assign _10391 = _10386 - _22192;
    assign _10392 = _10388 ? _10391 : _10386;
    assign _10393 = _10392[62:0];
    assign _10395 = { _10393,
                      _10394 };
    assign _10396 = _10395 < _22192;
    assign _10397 = ~ _10396;
    assign _10385 = _9933[13:13];
    assign _10382 = _10377 - _22192;
    assign _10383 = _10379 ? _10382 : _10377;
    assign _10384 = _10383[62:0];
    assign _10386 = { _10384,
                      _10385 };
    assign _10387 = _10386 < _22192;
    assign _10388 = ~ _10387;
    assign _10376 = _9933[14:14];
    assign _10373 = _10368 - _22192;
    assign _10374 = _10370 ? _10373 : _10368;
    assign _10375 = _10374[62:0];
    assign _10377 = { _10375,
                      _10376 };
    assign _10378 = _10377 < _22192;
    assign _10379 = ~ _10378;
    assign _10367 = _9933[15:15];
    assign _10364 = _10359 - _22192;
    assign _10365 = _10361 ? _10364 : _10359;
    assign _10366 = _10365[62:0];
    assign _10368 = { _10366,
                      _10367 };
    assign _10369 = _10368 < _22192;
    assign _10370 = ~ _10369;
    assign _10358 = _9933[16:16];
    assign _10355 = _10350 - _22192;
    assign _10356 = _10352 ? _10355 : _10350;
    assign _10357 = _10356[62:0];
    assign _10359 = { _10357,
                      _10358 };
    assign _10360 = _10359 < _22192;
    assign _10361 = ~ _10360;
    assign _10349 = _9933[17:17];
    assign _10346 = _10341 - _22192;
    assign _10347 = _10343 ? _10346 : _10341;
    assign _10348 = _10347[62:0];
    assign _10350 = { _10348,
                      _10349 };
    assign _10351 = _10350 < _22192;
    assign _10352 = ~ _10351;
    assign _10340 = _9933[18:18];
    assign _10337 = _10332 - _22192;
    assign _10338 = _10334 ? _10337 : _10332;
    assign _10339 = _10338[62:0];
    assign _10341 = { _10339,
                      _10340 };
    assign _10342 = _10341 < _22192;
    assign _10343 = ~ _10342;
    assign _10331 = _9933[19:19];
    assign _10328 = _10323 - _22192;
    assign _10329 = _10325 ? _10328 : _10323;
    assign _10330 = _10329[62:0];
    assign _10332 = { _10330,
                      _10331 };
    assign _10333 = _10332 < _22192;
    assign _10334 = ~ _10333;
    assign _10322 = _9933[20:20];
    assign _10319 = _10314 - _22192;
    assign _10320 = _10316 ? _10319 : _10314;
    assign _10321 = _10320[62:0];
    assign _10323 = { _10321,
                      _10322 };
    assign _10324 = _10323 < _22192;
    assign _10325 = ~ _10324;
    assign _10313 = _9933[21:21];
    assign _10310 = _10305 - _22192;
    assign _10311 = _10307 ? _10310 : _10305;
    assign _10312 = _10311[62:0];
    assign _10314 = { _10312,
                      _10313 };
    assign _10315 = _10314 < _22192;
    assign _10316 = ~ _10315;
    assign _10304 = _9933[22:22];
    assign _10301 = _10296 - _22192;
    assign _10302 = _10298 ? _10301 : _10296;
    assign _10303 = _10302[62:0];
    assign _10305 = { _10303,
                      _10304 };
    assign _10306 = _10305 < _22192;
    assign _10307 = ~ _10306;
    assign _10295 = _9933[23:23];
    assign _10292 = _10287 - _22192;
    assign _10293 = _10289 ? _10292 : _10287;
    assign _10294 = _10293[62:0];
    assign _10296 = { _10294,
                      _10295 };
    assign _10297 = _10296 < _22192;
    assign _10298 = ~ _10297;
    assign _10286 = _9933[24:24];
    assign _10283 = _10278 - _22192;
    assign _10284 = _10280 ? _10283 : _10278;
    assign _10285 = _10284[62:0];
    assign _10287 = { _10285,
                      _10286 };
    assign _10288 = _10287 < _22192;
    assign _10289 = ~ _10288;
    assign _10277 = _9933[25:25];
    assign _10274 = _10269 - _22192;
    assign _10275 = _10271 ? _10274 : _10269;
    assign _10276 = _10275[62:0];
    assign _10278 = { _10276,
                      _10277 };
    assign _10279 = _10278 < _22192;
    assign _10280 = ~ _10279;
    assign _10268 = _9933[26:26];
    assign _10265 = _10260 - _22192;
    assign _10266 = _10262 ? _10265 : _10260;
    assign _10267 = _10266[62:0];
    assign _10269 = { _10267,
                      _10268 };
    assign _10270 = _10269 < _22192;
    assign _10271 = ~ _10270;
    assign _10259 = _9933[27:27];
    assign _10256 = _10251 - _22192;
    assign _10257 = _10253 ? _10256 : _10251;
    assign _10258 = _10257[62:0];
    assign _10260 = { _10258,
                      _10259 };
    assign _10261 = _10260 < _22192;
    assign _10262 = ~ _10261;
    assign _10250 = _9933[28:28];
    assign _10247 = _10242 - _22192;
    assign _10248 = _10244 ? _10247 : _10242;
    assign _10249 = _10248[62:0];
    assign _10251 = { _10249,
                      _10250 };
    assign _10252 = _10251 < _22192;
    assign _10253 = ~ _10252;
    assign _10241 = _9933[29:29];
    assign _10238 = _10233 - _22192;
    assign _10239 = _10235 ? _10238 : _10233;
    assign _10240 = _10239[62:0];
    assign _10242 = { _10240,
                      _10241 };
    assign _10243 = _10242 < _22192;
    assign _10244 = ~ _10243;
    assign _10232 = _9933[30:30];
    assign _10229 = _10224 - _22192;
    assign _10230 = _10226 ? _10229 : _10224;
    assign _10231 = _10230[62:0];
    assign _10233 = { _10231,
                      _10232 };
    assign _10234 = _10233 < _22192;
    assign _10235 = ~ _10234;
    assign _10223 = _9933[31:31];
    assign _10220 = _10215 - _22192;
    assign _10221 = _10217 ? _10220 : _10215;
    assign _10222 = _10221[62:0];
    assign _10224 = { _10222,
                      _10223 };
    assign _10225 = _10224 < _22192;
    assign _10226 = ~ _10225;
    assign _10214 = _9933[32:32];
    assign _10211 = _10206 - _22192;
    assign _10212 = _10208 ? _10211 : _10206;
    assign _10213 = _10212[62:0];
    assign _10215 = { _10213,
                      _10214 };
    assign _10216 = _10215 < _22192;
    assign _10217 = ~ _10216;
    assign _10205 = _9933[33:33];
    assign _10202 = _10197 - _22192;
    assign _10203 = _10199 ? _10202 : _10197;
    assign _10204 = _10203[62:0];
    assign _10206 = { _10204,
                      _10205 };
    assign _10207 = _10206 < _22192;
    assign _10208 = ~ _10207;
    assign _10196 = _9933[34:34];
    assign _10193 = _10188 - _22192;
    assign _10194 = _10190 ? _10193 : _10188;
    assign _10195 = _10194[62:0];
    assign _10197 = { _10195,
                      _10196 };
    assign _10198 = _10197 < _22192;
    assign _10199 = ~ _10198;
    assign _10187 = _9933[35:35];
    assign _10184 = _10179 - _22192;
    assign _10185 = _10181 ? _10184 : _10179;
    assign _10186 = _10185[62:0];
    assign _10188 = { _10186,
                      _10187 };
    assign _10189 = _10188 < _22192;
    assign _10190 = ~ _10189;
    assign _10178 = _9933[36:36];
    assign _10175 = _10170 - _22192;
    assign _10176 = _10172 ? _10175 : _10170;
    assign _10177 = _10176[62:0];
    assign _10179 = { _10177,
                      _10178 };
    assign _10180 = _10179 < _22192;
    assign _10181 = ~ _10180;
    assign _10169 = _9933[37:37];
    assign _10166 = _10161 - _22192;
    assign _10167 = _10163 ? _10166 : _10161;
    assign _10168 = _10167[62:0];
    assign _10170 = { _10168,
                      _10169 };
    assign _10171 = _10170 < _22192;
    assign _10172 = ~ _10171;
    assign _10160 = _9933[38:38];
    assign _10157 = _10152 - _22192;
    assign _10158 = _10154 ? _10157 : _10152;
    assign _10159 = _10158[62:0];
    assign _10161 = { _10159,
                      _10160 };
    assign _10162 = _10161 < _22192;
    assign _10163 = ~ _10162;
    assign _10151 = _9933[39:39];
    assign _10148 = _10143 - _22192;
    assign _10149 = _10145 ? _10148 : _10143;
    assign _10150 = _10149[62:0];
    assign _10152 = { _10150,
                      _10151 };
    assign _10153 = _10152 < _22192;
    assign _10154 = ~ _10153;
    assign _10142 = _9933[40:40];
    assign _10139 = _10134 - _22192;
    assign _10140 = _10136 ? _10139 : _10134;
    assign _10141 = _10140[62:0];
    assign _10143 = { _10141,
                      _10142 };
    assign _10144 = _10143 < _22192;
    assign _10145 = ~ _10144;
    assign _10133 = _9933[41:41];
    assign _10130 = _10125 - _22192;
    assign _10131 = _10127 ? _10130 : _10125;
    assign _10132 = _10131[62:0];
    assign _10134 = { _10132,
                      _10133 };
    assign _10135 = _10134 < _22192;
    assign _10136 = ~ _10135;
    assign _10124 = _9933[42:42];
    assign _10121 = _10116 - _22192;
    assign _10122 = _10118 ? _10121 : _10116;
    assign _10123 = _10122[62:0];
    assign _10125 = { _10123,
                      _10124 };
    assign _10126 = _10125 < _22192;
    assign _10127 = ~ _10126;
    assign _10115 = _9933[43:43];
    assign _10112 = _10107 - _22192;
    assign _10113 = _10109 ? _10112 : _10107;
    assign _10114 = _10113[62:0];
    assign _10116 = { _10114,
                      _10115 };
    assign _10117 = _10116 < _22192;
    assign _10118 = ~ _10117;
    assign _10106 = _9933[44:44];
    assign _10103 = _10098 - _22192;
    assign _10104 = _10100 ? _10103 : _10098;
    assign _10105 = _10104[62:0];
    assign _10107 = { _10105,
                      _10106 };
    assign _10108 = _10107 < _22192;
    assign _10109 = ~ _10108;
    assign _10097 = _9933[45:45];
    assign _10094 = _10089 - _22192;
    assign _10095 = _10091 ? _10094 : _10089;
    assign _10096 = _10095[62:0];
    assign _10098 = { _10096,
                      _10097 };
    assign _10099 = _10098 < _22192;
    assign _10100 = ~ _10099;
    assign _10088 = _9933[46:46];
    assign _10085 = _10080 - _22192;
    assign _10086 = _10082 ? _10085 : _10080;
    assign _10087 = _10086[62:0];
    assign _10089 = { _10087,
                      _10088 };
    assign _10090 = _10089 < _22192;
    assign _10091 = ~ _10090;
    assign _10079 = _9933[47:47];
    assign _10076 = _10071 - _22192;
    assign _10077 = _10073 ? _10076 : _10071;
    assign _10078 = _10077[62:0];
    assign _10080 = { _10078,
                      _10079 };
    assign _10081 = _10080 < _22192;
    assign _10082 = ~ _10081;
    assign _10070 = _9933[48:48];
    assign _10067 = _10062 - _22192;
    assign _10068 = _10064 ? _10067 : _10062;
    assign _10069 = _10068[62:0];
    assign _10071 = { _10069,
                      _10070 };
    assign _10072 = _10071 < _22192;
    assign _10073 = ~ _10072;
    assign _10061 = _9933[49:49];
    assign _10058 = _10053 - _22192;
    assign _10059 = _10055 ? _10058 : _10053;
    assign _10060 = _10059[62:0];
    assign _10062 = { _10060,
                      _10061 };
    assign _10063 = _10062 < _22192;
    assign _10064 = ~ _10063;
    assign _10052 = _9933[50:50];
    assign _10049 = _10044 - _22192;
    assign _10050 = _10046 ? _10049 : _10044;
    assign _10051 = _10050[62:0];
    assign _10053 = { _10051,
                      _10052 };
    assign _10054 = _10053 < _22192;
    assign _10055 = ~ _10054;
    assign _10043 = _9933[51:51];
    assign _10040 = _10035 - _22192;
    assign _10041 = _10037 ? _10040 : _10035;
    assign _10042 = _10041[62:0];
    assign _10044 = { _10042,
                      _10043 };
    assign _10045 = _10044 < _22192;
    assign _10046 = ~ _10045;
    assign _10034 = _9933[52:52];
    assign _10031 = _10026 - _22192;
    assign _10032 = _10028 ? _10031 : _10026;
    assign _10033 = _10032[62:0];
    assign _10035 = { _10033,
                      _10034 };
    assign _10036 = _10035 < _22192;
    assign _10037 = ~ _10036;
    assign _10025 = _9933[53:53];
    assign _10022 = _10017 - _22192;
    assign _10023 = _10019 ? _10022 : _10017;
    assign _10024 = _10023[62:0];
    assign _10026 = { _10024,
                      _10025 };
    assign _10027 = _10026 < _22192;
    assign _10028 = ~ _10027;
    assign _10016 = _9933[54:54];
    assign _10013 = _10008 - _22192;
    assign _10014 = _10010 ? _10013 : _10008;
    assign _10015 = _10014[62:0];
    assign _10017 = { _10015,
                      _10016 };
    assign _10018 = _10017 < _22192;
    assign _10019 = ~ _10018;
    assign _10007 = _9933[55:55];
    assign _10004 = _9999 - _22192;
    assign _10005 = _10001 ? _10004 : _9999;
    assign _10006 = _10005[62:0];
    assign _10008 = { _10006,
                      _10007 };
    assign _10009 = _10008 < _22192;
    assign _10010 = ~ _10009;
    assign _9998 = _9933[56:56];
    assign _9995 = _9990 - _22192;
    assign _9996 = _9992 ? _9995 : _9990;
    assign _9997 = _9996[62:0];
    assign _9999 = { _9997,
                     _9998 };
    assign _10000 = _9999 < _22192;
    assign _10001 = ~ _10000;
    assign _9989 = _9933[57:57];
    assign _9986 = _9981 - _22192;
    assign _9987 = _9983 ? _9986 : _9981;
    assign _9988 = _9987[62:0];
    assign _9990 = { _9988,
                     _9989 };
    assign _9991 = _9990 < _22192;
    assign _9992 = ~ _9991;
    assign _9980 = _9933[58:58];
    assign _9977 = _9972 - _22192;
    assign _9978 = _9974 ? _9977 : _9972;
    assign _9979 = _9978[62:0];
    assign _9981 = { _9979,
                     _9980 };
    assign _9982 = _9981 < _22192;
    assign _9983 = ~ _9982;
    assign _9971 = _9933[59:59];
    assign _9968 = _9963 - _22192;
    assign _9969 = _9965 ? _9968 : _9963;
    assign _9970 = _9969[62:0];
    assign _9972 = { _9970,
                     _9971 };
    assign _9973 = _9972 < _22192;
    assign _9974 = ~ _9973;
    assign _9962 = _9933[60:60];
    assign _9959 = _9954 - _22192;
    assign _9960 = _9956 ? _9959 : _9954;
    assign _9961 = _9960[62:0];
    assign _9963 = { _9961,
                     _9962 };
    assign _9964 = _9963 < _22192;
    assign _9965 = ~ _9964;
    assign _9953 = _9933[61:61];
    assign _9950 = _9945 - _22192;
    assign _9951 = _9947 ? _9950 : _9945;
    assign _9952 = _9951[62:0];
    assign _9954 = { _9952,
                     _9953 };
    assign _9955 = _9954 < _22192;
    assign _9956 = ~ _9955;
    assign _9944 = _9933[62:62];
    assign _9941 = _9935 - _22192;
    assign _9942 = _9938 ? _9941 : _9935;
    assign _9943 = _9942[62:0];
    assign _9945 = { _9943,
                     _9944 };
    assign _9946 = _9945 < _22192;
    assign _9947 = ~ _9946;
    assign _9931 = _9923 + _22186;
    assign _9932 = _9923 * _9931;
    assign _9933 = _9932[63:0];
    assign _9934 = _9933[63:63];
    assign _9935 = { _22185,
                     _9934 };
    assign _9937 = _9935 < _22192;
    assign _9938 = ~ _9937;
    assign _9939 = { _22185,
                     _9938 };
    assign _9940 = _9939[62:0];
    assign _9948 = { _9940,
                     _9947 };
    assign _9949 = _9948[62:0];
    assign _9957 = { _9949,
                     _9956 };
    assign _9958 = _9957[62:0];
    assign _9966 = { _9958,
                     _9965 };
    assign _9967 = _9966[62:0];
    assign _9975 = { _9967,
                     _9974 };
    assign _9976 = _9975[62:0];
    assign _9984 = { _9976,
                     _9983 };
    assign _9985 = _9984[62:0];
    assign _9993 = { _9985,
                     _9992 };
    assign _9994 = _9993[62:0];
    assign _10002 = { _9994,
                      _10001 };
    assign _10003 = _10002[62:0];
    assign _10011 = { _10003,
                      _10010 };
    assign _10012 = _10011[62:0];
    assign _10020 = { _10012,
                      _10019 };
    assign _10021 = _10020[62:0];
    assign _10029 = { _10021,
                      _10028 };
    assign _10030 = _10029[62:0];
    assign _10038 = { _10030,
                      _10037 };
    assign _10039 = _10038[62:0];
    assign _10047 = { _10039,
                      _10046 };
    assign _10048 = _10047[62:0];
    assign _10056 = { _10048,
                      _10055 };
    assign _10057 = _10056[62:0];
    assign _10065 = { _10057,
                      _10064 };
    assign _10066 = _10065[62:0];
    assign _10074 = { _10066,
                      _10073 };
    assign _10075 = _10074[62:0];
    assign _10083 = { _10075,
                      _10082 };
    assign _10084 = _10083[62:0];
    assign _10092 = { _10084,
                      _10091 };
    assign _10093 = _10092[62:0];
    assign _10101 = { _10093,
                      _10100 };
    assign _10102 = _10101[62:0];
    assign _10110 = { _10102,
                      _10109 };
    assign _10111 = _10110[62:0];
    assign _10119 = { _10111,
                      _10118 };
    assign _10120 = _10119[62:0];
    assign _10128 = { _10120,
                      _10127 };
    assign _10129 = _10128[62:0];
    assign _10137 = { _10129,
                      _10136 };
    assign _10138 = _10137[62:0];
    assign _10146 = { _10138,
                      _10145 };
    assign _10147 = _10146[62:0];
    assign _10155 = { _10147,
                      _10154 };
    assign _10156 = _10155[62:0];
    assign _10164 = { _10156,
                      _10163 };
    assign _10165 = _10164[62:0];
    assign _10173 = { _10165,
                      _10172 };
    assign _10174 = _10173[62:0];
    assign _10182 = { _10174,
                      _10181 };
    assign _10183 = _10182[62:0];
    assign _10191 = { _10183,
                      _10190 };
    assign _10192 = _10191[62:0];
    assign _10200 = { _10192,
                      _10199 };
    assign _10201 = _10200[62:0];
    assign _10209 = { _10201,
                      _10208 };
    assign _10210 = _10209[62:0];
    assign _10218 = { _10210,
                      _10217 };
    assign _10219 = _10218[62:0];
    assign _10227 = { _10219,
                      _10226 };
    assign _10228 = _10227[62:0];
    assign _10236 = { _10228,
                      _10235 };
    assign _10237 = _10236[62:0];
    assign _10245 = { _10237,
                      _10244 };
    assign _10246 = _10245[62:0];
    assign _10254 = { _10246,
                      _10253 };
    assign _10255 = _10254[62:0];
    assign _10263 = { _10255,
                      _10262 };
    assign _10264 = _10263[62:0];
    assign _10272 = { _10264,
                      _10271 };
    assign _10273 = _10272[62:0];
    assign _10281 = { _10273,
                      _10280 };
    assign _10282 = _10281[62:0];
    assign _10290 = { _10282,
                      _10289 };
    assign _10291 = _10290[62:0];
    assign _10299 = { _10291,
                      _10298 };
    assign _10300 = _10299[62:0];
    assign _10308 = { _10300,
                      _10307 };
    assign _10309 = _10308[62:0];
    assign _10317 = { _10309,
                      _10316 };
    assign _10318 = _10317[62:0];
    assign _10326 = { _10318,
                      _10325 };
    assign _10327 = _10326[62:0];
    assign _10335 = { _10327,
                      _10334 };
    assign _10336 = _10335[62:0];
    assign _10344 = { _10336,
                      _10343 };
    assign _10345 = _10344[62:0];
    assign _10353 = { _10345,
                      _10352 };
    assign _10354 = _10353[62:0];
    assign _10362 = { _10354,
                      _10361 };
    assign _10363 = _10362[62:0];
    assign _10371 = { _10363,
                      _10370 };
    assign _10372 = _10371[62:0];
    assign _10380 = { _10372,
                      _10379 };
    assign _10381 = _10380[62:0];
    assign _10389 = { _10381,
                      _10388 };
    assign _10390 = _10389[62:0];
    assign _10398 = { _10390,
                      _10397 };
    assign _10399 = _10398[62:0];
    assign _10407 = { _10399,
                      _10406 };
    assign _10408 = _10407[62:0];
    assign _10416 = { _10408,
                      _10415 };
    assign _10417 = _10416[62:0];
    assign _10425 = { _10417,
                      _10424 };
    assign _10426 = _10425[62:0];
    assign _10434 = { _10426,
                      _10433 };
    assign _10435 = _10434[62:0];
    assign _10443 = { _10435,
                      _10442 };
    assign _10444 = _10443[62:0];
    assign _10452 = { _10444,
                      _10451 };
    assign _10453 = _10452[62:0];
    assign _10461 = { _10453,
                      _10460 };
    assign _10462 = _10461[62:0];
    assign _10470 = { _10462,
                      _10469 };
    assign _10471 = _10470[62:0];
    assign _10479 = { _10471,
                      _10478 };
    assign _10480 = _10479[62:0];
    assign _10488 = { _10480,
                      _10487 };
    assign _10489 = _10488[62:0];
    assign _10497 = { _10489,
                      _10496 };
    assign _10498 = _10497[62:0];
    assign _10506 = { _10498,
                      _10505 };
    assign _10507 = _8771 * _10506;
    assign _10508 = _10507[63:0];
    assign _9919 = _9351[0:0];
    assign _9916 = _9911 - _8771;
    assign _9917 = _9913 ? _9916 : _9911;
    assign _9918 = _9917[62:0];
    assign _9920 = { _9918,
                     _9919 };
    assign _9921 = _9920 < _8771;
    assign _9922 = ~ _9921;
    assign _9910 = _9351[1:1];
    assign _9907 = _9902 - _8771;
    assign _9908 = _9904 ? _9907 : _9902;
    assign _9909 = _9908[62:0];
    assign _9911 = { _9909,
                     _9910 };
    assign _9912 = _9911 < _8771;
    assign _9913 = ~ _9912;
    assign _9901 = _9351[2:2];
    assign _9898 = _9893 - _8771;
    assign _9899 = _9895 ? _9898 : _9893;
    assign _9900 = _9899[62:0];
    assign _9902 = { _9900,
                     _9901 };
    assign _9903 = _9902 < _8771;
    assign _9904 = ~ _9903;
    assign _9892 = _9351[3:3];
    assign _9889 = _9884 - _8771;
    assign _9890 = _9886 ? _9889 : _9884;
    assign _9891 = _9890[62:0];
    assign _9893 = { _9891,
                     _9892 };
    assign _9894 = _9893 < _8771;
    assign _9895 = ~ _9894;
    assign _9883 = _9351[4:4];
    assign _9880 = _9875 - _8771;
    assign _9881 = _9877 ? _9880 : _9875;
    assign _9882 = _9881[62:0];
    assign _9884 = { _9882,
                     _9883 };
    assign _9885 = _9884 < _8771;
    assign _9886 = ~ _9885;
    assign _9874 = _9351[5:5];
    assign _9871 = _9866 - _8771;
    assign _9872 = _9868 ? _9871 : _9866;
    assign _9873 = _9872[62:0];
    assign _9875 = { _9873,
                     _9874 };
    assign _9876 = _9875 < _8771;
    assign _9877 = ~ _9876;
    assign _9865 = _9351[6:6];
    assign _9862 = _9857 - _8771;
    assign _9863 = _9859 ? _9862 : _9857;
    assign _9864 = _9863[62:0];
    assign _9866 = { _9864,
                     _9865 };
    assign _9867 = _9866 < _8771;
    assign _9868 = ~ _9867;
    assign _9856 = _9351[7:7];
    assign _9853 = _9848 - _8771;
    assign _9854 = _9850 ? _9853 : _9848;
    assign _9855 = _9854[62:0];
    assign _9857 = { _9855,
                     _9856 };
    assign _9858 = _9857 < _8771;
    assign _9859 = ~ _9858;
    assign _9847 = _9351[8:8];
    assign _9844 = _9839 - _8771;
    assign _9845 = _9841 ? _9844 : _9839;
    assign _9846 = _9845[62:0];
    assign _9848 = { _9846,
                     _9847 };
    assign _9849 = _9848 < _8771;
    assign _9850 = ~ _9849;
    assign _9838 = _9351[9:9];
    assign _9835 = _9830 - _8771;
    assign _9836 = _9832 ? _9835 : _9830;
    assign _9837 = _9836[62:0];
    assign _9839 = { _9837,
                     _9838 };
    assign _9840 = _9839 < _8771;
    assign _9841 = ~ _9840;
    assign _9829 = _9351[10:10];
    assign _9826 = _9821 - _8771;
    assign _9827 = _9823 ? _9826 : _9821;
    assign _9828 = _9827[62:0];
    assign _9830 = { _9828,
                     _9829 };
    assign _9831 = _9830 < _8771;
    assign _9832 = ~ _9831;
    assign _9820 = _9351[11:11];
    assign _9817 = _9812 - _8771;
    assign _9818 = _9814 ? _9817 : _9812;
    assign _9819 = _9818[62:0];
    assign _9821 = { _9819,
                     _9820 };
    assign _9822 = _9821 < _8771;
    assign _9823 = ~ _9822;
    assign _9811 = _9351[12:12];
    assign _9808 = _9803 - _8771;
    assign _9809 = _9805 ? _9808 : _9803;
    assign _9810 = _9809[62:0];
    assign _9812 = { _9810,
                     _9811 };
    assign _9813 = _9812 < _8771;
    assign _9814 = ~ _9813;
    assign _9802 = _9351[13:13];
    assign _9799 = _9794 - _8771;
    assign _9800 = _9796 ? _9799 : _9794;
    assign _9801 = _9800[62:0];
    assign _9803 = { _9801,
                     _9802 };
    assign _9804 = _9803 < _8771;
    assign _9805 = ~ _9804;
    assign _9793 = _9351[14:14];
    assign _9790 = _9785 - _8771;
    assign _9791 = _9787 ? _9790 : _9785;
    assign _9792 = _9791[62:0];
    assign _9794 = { _9792,
                     _9793 };
    assign _9795 = _9794 < _8771;
    assign _9796 = ~ _9795;
    assign _9784 = _9351[15:15];
    assign _9781 = _9776 - _8771;
    assign _9782 = _9778 ? _9781 : _9776;
    assign _9783 = _9782[62:0];
    assign _9785 = { _9783,
                     _9784 };
    assign _9786 = _9785 < _8771;
    assign _9787 = ~ _9786;
    assign _9775 = _9351[16:16];
    assign _9772 = _9767 - _8771;
    assign _9773 = _9769 ? _9772 : _9767;
    assign _9774 = _9773[62:0];
    assign _9776 = { _9774,
                     _9775 };
    assign _9777 = _9776 < _8771;
    assign _9778 = ~ _9777;
    assign _9766 = _9351[17:17];
    assign _9763 = _9758 - _8771;
    assign _9764 = _9760 ? _9763 : _9758;
    assign _9765 = _9764[62:0];
    assign _9767 = { _9765,
                     _9766 };
    assign _9768 = _9767 < _8771;
    assign _9769 = ~ _9768;
    assign _9757 = _9351[18:18];
    assign _9754 = _9749 - _8771;
    assign _9755 = _9751 ? _9754 : _9749;
    assign _9756 = _9755[62:0];
    assign _9758 = { _9756,
                     _9757 };
    assign _9759 = _9758 < _8771;
    assign _9760 = ~ _9759;
    assign _9748 = _9351[19:19];
    assign _9745 = _9740 - _8771;
    assign _9746 = _9742 ? _9745 : _9740;
    assign _9747 = _9746[62:0];
    assign _9749 = { _9747,
                     _9748 };
    assign _9750 = _9749 < _8771;
    assign _9751 = ~ _9750;
    assign _9739 = _9351[20:20];
    assign _9736 = _9731 - _8771;
    assign _9737 = _9733 ? _9736 : _9731;
    assign _9738 = _9737[62:0];
    assign _9740 = { _9738,
                     _9739 };
    assign _9741 = _9740 < _8771;
    assign _9742 = ~ _9741;
    assign _9730 = _9351[21:21];
    assign _9727 = _9722 - _8771;
    assign _9728 = _9724 ? _9727 : _9722;
    assign _9729 = _9728[62:0];
    assign _9731 = { _9729,
                     _9730 };
    assign _9732 = _9731 < _8771;
    assign _9733 = ~ _9732;
    assign _9721 = _9351[22:22];
    assign _9718 = _9713 - _8771;
    assign _9719 = _9715 ? _9718 : _9713;
    assign _9720 = _9719[62:0];
    assign _9722 = { _9720,
                     _9721 };
    assign _9723 = _9722 < _8771;
    assign _9724 = ~ _9723;
    assign _9712 = _9351[23:23];
    assign _9709 = _9704 - _8771;
    assign _9710 = _9706 ? _9709 : _9704;
    assign _9711 = _9710[62:0];
    assign _9713 = { _9711,
                     _9712 };
    assign _9714 = _9713 < _8771;
    assign _9715 = ~ _9714;
    assign _9703 = _9351[24:24];
    assign _9700 = _9695 - _8771;
    assign _9701 = _9697 ? _9700 : _9695;
    assign _9702 = _9701[62:0];
    assign _9704 = { _9702,
                     _9703 };
    assign _9705 = _9704 < _8771;
    assign _9706 = ~ _9705;
    assign _9694 = _9351[25:25];
    assign _9691 = _9686 - _8771;
    assign _9692 = _9688 ? _9691 : _9686;
    assign _9693 = _9692[62:0];
    assign _9695 = { _9693,
                     _9694 };
    assign _9696 = _9695 < _8771;
    assign _9697 = ~ _9696;
    assign _9685 = _9351[26:26];
    assign _9682 = _9677 - _8771;
    assign _9683 = _9679 ? _9682 : _9677;
    assign _9684 = _9683[62:0];
    assign _9686 = { _9684,
                     _9685 };
    assign _9687 = _9686 < _8771;
    assign _9688 = ~ _9687;
    assign _9676 = _9351[27:27];
    assign _9673 = _9668 - _8771;
    assign _9674 = _9670 ? _9673 : _9668;
    assign _9675 = _9674[62:0];
    assign _9677 = { _9675,
                     _9676 };
    assign _9678 = _9677 < _8771;
    assign _9679 = ~ _9678;
    assign _9667 = _9351[28:28];
    assign _9664 = _9659 - _8771;
    assign _9665 = _9661 ? _9664 : _9659;
    assign _9666 = _9665[62:0];
    assign _9668 = { _9666,
                     _9667 };
    assign _9669 = _9668 < _8771;
    assign _9670 = ~ _9669;
    assign _9658 = _9351[29:29];
    assign _9655 = _9650 - _8771;
    assign _9656 = _9652 ? _9655 : _9650;
    assign _9657 = _9656[62:0];
    assign _9659 = { _9657,
                     _9658 };
    assign _9660 = _9659 < _8771;
    assign _9661 = ~ _9660;
    assign _9649 = _9351[30:30];
    assign _9646 = _9641 - _8771;
    assign _9647 = _9643 ? _9646 : _9641;
    assign _9648 = _9647[62:0];
    assign _9650 = { _9648,
                     _9649 };
    assign _9651 = _9650 < _8771;
    assign _9652 = ~ _9651;
    assign _9640 = _9351[31:31];
    assign _9637 = _9632 - _8771;
    assign _9638 = _9634 ? _9637 : _9632;
    assign _9639 = _9638[62:0];
    assign _9641 = { _9639,
                     _9640 };
    assign _9642 = _9641 < _8771;
    assign _9643 = ~ _9642;
    assign _9631 = _9351[32:32];
    assign _9628 = _9623 - _8771;
    assign _9629 = _9625 ? _9628 : _9623;
    assign _9630 = _9629[62:0];
    assign _9632 = { _9630,
                     _9631 };
    assign _9633 = _9632 < _8771;
    assign _9634 = ~ _9633;
    assign _9622 = _9351[33:33];
    assign _9619 = _9614 - _8771;
    assign _9620 = _9616 ? _9619 : _9614;
    assign _9621 = _9620[62:0];
    assign _9623 = { _9621,
                     _9622 };
    assign _9624 = _9623 < _8771;
    assign _9625 = ~ _9624;
    assign _9613 = _9351[34:34];
    assign _9610 = _9605 - _8771;
    assign _9611 = _9607 ? _9610 : _9605;
    assign _9612 = _9611[62:0];
    assign _9614 = { _9612,
                     _9613 };
    assign _9615 = _9614 < _8771;
    assign _9616 = ~ _9615;
    assign _9604 = _9351[35:35];
    assign _9601 = _9596 - _8771;
    assign _9602 = _9598 ? _9601 : _9596;
    assign _9603 = _9602[62:0];
    assign _9605 = { _9603,
                     _9604 };
    assign _9606 = _9605 < _8771;
    assign _9607 = ~ _9606;
    assign _9595 = _9351[36:36];
    assign _9592 = _9587 - _8771;
    assign _9593 = _9589 ? _9592 : _9587;
    assign _9594 = _9593[62:0];
    assign _9596 = { _9594,
                     _9595 };
    assign _9597 = _9596 < _8771;
    assign _9598 = ~ _9597;
    assign _9586 = _9351[37:37];
    assign _9583 = _9578 - _8771;
    assign _9584 = _9580 ? _9583 : _9578;
    assign _9585 = _9584[62:0];
    assign _9587 = { _9585,
                     _9586 };
    assign _9588 = _9587 < _8771;
    assign _9589 = ~ _9588;
    assign _9577 = _9351[38:38];
    assign _9574 = _9569 - _8771;
    assign _9575 = _9571 ? _9574 : _9569;
    assign _9576 = _9575[62:0];
    assign _9578 = { _9576,
                     _9577 };
    assign _9579 = _9578 < _8771;
    assign _9580 = ~ _9579;
    assign _9568 = _9351[39:39];
    assign _9565 = _9560 - _8771;
    assign _9566 = _9562 ? _9565 : _9560;
    assign _9567 = _9566[62:0];
    assign _9569 = { _9567,
                     _9568 };
    assign _9570 = _9569 < _8771;
    assign _9571 = ~ _9570;
    assign _9559 = _9351[40:40];
    assign _9556 = _9551 - _8771;
    assign _9557 = _9553 ? _9556 : _9551;
    assign _9558 = _9557[62:0];
    assign _9560 = { _9558,
                     _9559 };
    assign _9561 = _9560 < _8771;
    assign _9562 = ~ _9561;
    assign _9550 = _9351[41:41];
    assign _9547 = _9542 - _8771;
    assign _9548 = _9544 ? _9547 : _9542;
    assign _9549 = _9548[62:0];
    assign _9551 = { _9549,
                     _9550 };
    assign _9552 = _9551 < _8771;
    assign _9553 = ~ _9552;
    assign _9541 = _9351[42:42];
    assign _9538 = _9533 - _8771;
    assign _9539 = _9535 ? _9538 : _9533;
    assign _9540 = _9539[62:0];
    assign _9542 = { _9540,
                     _9541 };
    assign _9543 = _9542 < _8771;
    assign _9544 = ~ _9543;
    assign _9532 = _9351[43:43];
    assign _9529 = _9524 - _8771;
    assign _9530 = _9526 ? _9529 : _9524;
    assign _9531 = _9530[62:0];
    assign _9533 = { _9531,
                     _9532 };
    assign _9534 = _9533 < _8771;
    assign _9535 = ~ _9534;
    assign _9523 = _9351[44:44];
    assign _9520 = _9515 - _8771;
    assign _9521 = _9517 ? _9520 : _9515;
    assign _9522 = _9521[62:0];
    assign _9524 = { _9522,
                     _9523 };
    assign _9525 = _9524 < _8771;
    assign _9526 = ~ _9525;
    assign _9514 = _9351[45:45];
    assign _9511 = _9506 - _8771;
    assign _9512 = _9508 ? _9511 : _9506;
    assign _9513 = _9512[62:0];
    assign _9515 = { _9513,
                     _9514 };
    assign _9516 = _9515 < _8771;
    assign _9517 = ~ _9516;
    assign _9505 = _9351[46:46];
    assign _9502 = _9497 - _8771;
    assign _9503 = _9499 ? _9502 : _9497;
    assign _9504 = _9503[62:0];
    assign _9506 = { _9504,
                     _9505 };
    assign _9507 = _9506 < _8771;
    assign _9508 = ~ _9507;
    assign _9496 = _9351[47:47];
    assign _9493 = _9488 - _8771;
    assign _9494 = _9490 ? _9493 : _9488;
    assign _9495 = _9494[62:0];
    assign _9497 = { _9495,
                     _9496 };
    assign _9498 = _9497 < _8771;
    assign _9499 = ~ _9498;
    assign _9487 = _9351[48:48];
    assign _9484 = _9479 - _8771;
    assign _9485 = _9481 ? _9484 : _9479;
    assign _9486 = _9485[62:0];
    assign _9488 = { _9486,
                     _9487 };
    assign _9489 = _9488 < _8771;
    assign _9490 = ~ _9489;
    assign _9478 = _9351[49:49];
    assign _9475 = _9470 - _8771;
    assign _9476 = _9472 ? _9475 : _9470;
    assign _9477 = _9476[62:0];
    assign _9479 = { _9477,
                     _9478 };
    assign _9480 = _9479 < _8771;
    assign _9481 = ~ _9480;
    assign _9469 = _9351[50:50];
    assign _9466 = _9461 - _8771;
    assign _9467 = _9463 ? _9466 : _9461;
    assign _9468 = _9467[62:0];
    assign _9470 = { _9468,
                     _9469 };
    assign _9471 = _9470 < _8771;
    assign _9472 = ~ _9471;
    assign _9460 = _9351[51:51];
    assign _9457 = _9452 - _8771;
    assign _9458 = _9454 ? _9457 : _9452;
    assign _9459 = _9458[62:0];
    assign _9461 = { _9459,
                     _9460 };
    assign _9462 = _9461 < _8771;
    assign _9463 = ~ _9462;
    assign _9451 = _9351[52:52];
    assign _9448 = _9443 - _8771;
    assign _9449 = _9445 ? _9448 : _9443;
    assign _9450 = _9449[62:0];
    assign _9452 = { _9450,
                     _9451 };
    assign _9453 = _9452 < _8771;
    assign _9454 = ~ _9453;
    assign _9442 = _9351[53:53];
    assign _9439 = _9434 - _8771;
    assign _9440 = _9436 ? _9439 : _9434;
    assign _9441 = _9440[62:0];
    assign _9443 = { _9441,
                     _9442 };
    assign _9444 = _9443 < _8771;
    assign _9445 = ~ _9444;
    assign _9433 = _9351[54:54];
    assign _9430 = _9425 - _8771;
    assign _9431 = _9427 ? _9430 : _9425;
    assign _9432 = _9431[62:0];
    assign _9434 = { _9432,
                     _9433 };
    assign _9435 = _9434 < _8771;
    assign _9436 = ~ _9435;
    assign _9424 = _9351[55:55];
    assign _9421 = _9416 - _8771;
    assign _9422 = _9418 ? _9421 : _9416;
    assign _9423 = _9422[62:0];
    assign _9425 = { _9423,
                     _9424 };
    assign _9426 = _9425 < _8771;
    assign _9427 = ~ _9426;
    assign _9415 = _9351[56:56];
    assign _9412 = _9407 - _8771;
    assign _9413 = _9409 ? _9412 : _9407;
    assign _9414 = _9413[62:0];
    assign _9416 = { _9414,
                     _9415 };
    assign _9417 = _9416 < _8771;
    assign _9418 = ~ _9417;
    assign _9406 = _9351[57:57];
    assign _9403 = _9398 - _8771;
    assign _9404 = _9400 ? _9403 : _9398;
    assign _9405 = _9404[62:0];
    assign _9407 = { _9405,
                     _9406 };
    assign _9408 = _9407 < _8771;
    assign _9409 = ~ _9408;
    assign _9397 = _9351[58:58];
    assign _9394 = _9389 - _8771;
    assign _9395 = _9391 ? _9394 : _9389;
    assign _9396 = _9395[62:0];
    assign _9398 = { _9396,
                     _9397 };
    assign _9399 = _9398 < _8771;
    assign _9400 = ~ _9399;
    assign _9388 = _9351[59:59];
    assign _9385 = _9380 - _8771;
    assign _9386 = _9382 ? _9385 : _9380;
    assign _9387 = _9386[62:0];
    assign _9389 = { _9387,
                     _9388 };
    assign _9390 = _9389 < _8771;
    assign _9391 = ~ _9390;
    assign _9379 = _9351[60:60];
    assign _9376 = _9371 - _8771;
    assign _9377 = _9373 ? _9376 : _9371;
    assign _9378 = _9377[62:0];
    assign _9380 = { _9378,
                     _9379 };
    assign _9381 = _9380 < _8771;
    assign _9382 = ~ _9381;
    assign _9370 = _9351[61:61];
    assign _9367 = _9362 - _8771;
    assign _9368 = _9364 ? _9367 : _9362;
    assign _9369 = _9368[62:0];
    assign _9371 = { _9369,
                     _9370 };
    assign _9372 = _9371 < _8771;
    assign _9373 = ~ _9372;
    assign _9361 = _9351[62:62];
    assign _9358 = _9353 - _8771;
    assign _9359 = _9355 ? _9358 : _9353;
    assign _9360 = _9359[62:0];
    assign _9362 = { _9360,
                     _9361 };
    assign _9363 = _9362 < _8771;
    assign _9364 = ~ _9363;
    assign _9351 = _8763 - _9345;
    assign _9352 = _9351[63:63];
    assign _9353 = { _22185,
                     _9352 };
    assign _9354 = _9353 < _8771;
    assign _9355 = ~ _9354;
    assign _9356 = { _22185,
                     _9355 };
    assign _9357 = _9356[62:0];
    assign _9365 = { _9357,
                     _9364 };
    assign _9366 = _9365[62:0];
    assign _9374 = { _9366,
                     _9373 };
    assign _9375 = _9374[62:0];
    assign _9383 = { _9375,
                     _9382 };
    assign _9384 = _9383[62:0];
    assign _9392 = { _9384,
                     _9391 };
    assign _9393 = _9392[62:0];
    assign _9401 = { _9393,
                     _9400 };
    assign _9402 = _9401[62:0];
    assign _9410 = { _9402,
                     _9409 };
    assign _9411 = _9410[62:0];
    assign _9419 = { _9411,
                     _9418 };
    assign _9420 = _9419[62:0];
    assign _9428 = { _9420,
                     _9427 };
    assign _9429 = _9428[62:0];
    assign _9437 = { _9429,
                     _9436 };
    assign _9438 = _9437[62:0];
    assign _9446 = { _9438,
                     _9445 };
    assign _9447 = _9446[62:0];
    assign _9455 = { _9447,
                     _9454 };
    assign _9456 = _9455[62:0];
    assign _9464 = { _9456,
                     _9463 };
    assign _9465 = _9464[62:0];
    assign _9473 = { _9465,
                     _9472 };
    assign _9474 = _9473[62:0];
    assign _9482 = { _9474,
                     _9481 };
    assign _9483 = _9482[62:0];
    assign _9491 = { _9483,
                     _9490 };
    assign _9492 = _9491[62:0];
    assign _9500 = { _9492,
                     _9499 };
    assign _9501 = _9500[62:0];
    assign _9509 = { _9501,
                     _9508 };
    assign _9510 = _9509[62:0];
    assign _9518 = { _9510,
                     _9517 };
    assign _9519 = _9518[62:0];
    assign _9527 = { _9519,
                     _9526 };
    assign _9528 = _9527[62:0];
    assign _9536 = { _9528,
                     _9535 };
    assign _9537 = _9536[62:0];
    assign _9545 = { _9537,
                     _9544 };
    assign _9546 = _9545[62:0];
    assign _9554 = { _9546,
                     _9553 };
    assign _9555 = _9554[62:0];
    assign _9563 = { _9555,
                     _9562 };
    assign _9564 = _9563[62:0];
    assign _9572 = { _9564,
                     _9571 };
    assign _9573 = _9572[62:0];
    assign _9581 = { _9573,
                     _9580 };
    assign _9582 = _9581[62:0];
    assign _9590 = { _9582,
                     _9589 };
    assign _9591 = _9590[62:0];
    assign _9599 = { _9591,
                     _9598 };
    assign _9600 = _9599[62:0];
    assign _9608 = { _9600,
                     _9607 };
    assign _9609 = _9608[62:0];
    assign _9617 = { _9609,
                     _9616 };
    assign _9618 = _9617[62:0];
    assign _9626 = { _9618,
                     _9625 };
    assign _9627 = _9626[62:0];
    assign _9635 = { _9627,
                     _9634 };
    assign _9636 = _9635[62:0];
    assign _9644 = { _9636,
                     _9643 };
    assign _9645 = _9644[62:0];
    assign _9653 = { _9645,
                     _9652 };
    assign _9654 = _9653[62:0];
    assign _9662 = { _9654,
                     _9661 };
    assign _9663 = _9662[62:0];
    assign _9671 = { _9663,
                     _9670 };
    assign _9672 = _9671[62:0];
    assign _9680 = { _9672,
                     _9679 };
    assign _9681 = _9680[62:0];
    assign _9689 = { _9681,
                     _9688 };
    assign _9690 = _9689[62:0];
    assign _9698 = { _9690,
                     _9697 };
    assign _9699 = _9698[62:0];
    assign _9707 = { _9699,
                     _9706 };
    assign _9708 = _9707[62:0];
    assign _9716 = { _9708,
                     _9715 };
    assign _9717 = _9716[62:0];
    assign _9725 = { _9717,
                     _9724 };
    assign _9726 = _9725[62:0];
    assign _9734 = { _9726,
                     _9733 };
    assign _9735 = _9734[62:0];
    assign _9743 = { _9735,
                     _9742 };
    assign _9744 = _9743[62:0];
    assign _9752 = { _9744,
                     _9751 };
    assign _9753 = _9752[62:0];
    assign _9761 = { _9753,
                     _9760 };
    assign _9762 = _9761[62:0];
    assign _9770 = { _9762,
                     _9769 };
    assign _9771 = _9770[62:0];
    assign _9779 = { _9771,
                     _9778 };
    assign _9780 = _9779[62:0];
    assign _9788 = { _9780,
                     _9787 };
    assign _9789 = _9788[62:0];
    assign _9797 = { _9789,
                     _9796 };
    assign _9798 = _9797[62:0];
    assign _9806 = { _9798,
                     _9805 };
    assign _9807 = _9806[62:0];
    assign _9815 = { _9807,
                     _9814 };
    assign _9816 = _9815[62:0];
    assign _9824 = { _9816,
                     _9823 };
    assign _9825 = _9824[62:0];
    assign _9833 = { _9825,
                     _9832 };
    assign _9834 = _9833[62:0];
    assign _9842 = { _9834,
                     _9841 };
    assign _9843 = _9842[62:0];
    assign _9851 = { _9843,
                     _9850 };
    assign _9852 = _9851[62:0];
    assign _9860 = { _9852,
                     _9859 };
    assign _9861 = _9860[62:0];
    assign _9869 = { _9861,
                     _9868 };
    assign _9870 = _9869[62:0];
    assign _9878 = { _9870,
                     _9877 };
    assign _9879 = _9878[62:0];
    assign _9887 = { _9879,
                     _9886 };
    assign _9888 = _9887[62:0];
    assign _9896 = { _9888,
                     _9895 };
    assign _9897 = _9896[62:0];
    assign _9905 = { _9897,
                     _9904 };
    assign _9906 = _9905[62:0];
    assign _9914 = { _9906,
                     _9913 };
    assign _9915 = _9914[62:0];
    assign _9923 = { _9915,
                     _9922 };
    assign _9925 = _9923 + _22186;
    assign _9926 = _9925 * _9345;
    assign _9927 = _9926[63:0];
    assign _10509 = _9927 + _10508;
    assign _9337 = _8768[0:0];
    assign _9334 = _9329 - _8771;
    assign _9335 = _9331 ? _9334 : _9329;
    assign _9336 = _9335[62:0];
    assign _9338 = { _9336,
                     _9337 };
    assign _9339 = _9338 < _8771;
    assign _9340 = ~ _9339;
    assign _9328 = _8768[1:1];
    assign _9325 = _9320 - _8771;
    assign _9326 = _9322 ? _9325 : _9320;
    assign _9327 = _9326[62:0];
    assign _9329 = { _9327,
                     _9328 };
    assign _9330 = _9329 < _8771;
    assign _9331 = ~ _9330;
    assign _9319 = _8768[2:2];
    assign _9316 = _9311 - _8771;
    assign _9317 = _9313 ? _9316 : _9311;
    assign _9318 = _9317[62:0];
    assign _9320 = { _9318,
                     _9319 };
    assign _9321 = _9320 < _8771;
    assign _9322 = ~ _9321;
    assign _9310 = _8768[3:3];
    assign _9307 = _9302 - _8771;
    assign _9308 = _9304 ? _9307 : _9302;
    assign _9309 = _9308[62:0];
    assign _9311 = { _9309,
                     _9310 };
    assign _9312 = _9311 < _8771;
    assign _9313 = ~ _9312;
    assign _9301 = _8768[4:4];
    assign _9298 = _9293 - _8771;
    assign _9299 = _9295 ? _9298 : _9293;
    assign _9300 = _9299[62:0];
    assign _9302 = { _9300,
                     _9301 };
    assign _9303 = _9302 < _8771;
    assign _9304 = ~ _9303;
    assign _9292 = _8768[5:5];
    assign _9289 = _9284 - _8771;
    assign _9290 = _9286 ? _9289 : _9284;
    assign _9291 = _9290[62:0];
    assign _9293 = { _9291,
                     _9292 };
    assign _9294 = _9293 < _8771;
    assign _9295 = ~ _9294;
    assign _9283 = _8768[6:6];
    assign _9280 = _9275 - _8771;
    assign _9281 = _9277 ? _9280 : _9275;
    assign _9282 = _9281[62:0];
    assign _9284 = { _9282,
                     _9283 };
    assign _9285 = _9284 < _8771;
    assign _9286 = ~ _9285;
    assign _9274 = _8768[7:7];
    assign _9271 = _9266 - _8771;
    assign _9272 = _9268 ? _9271 : _9266;
    assign _9273 = _9272[62:0];
    assign _9275 = { _9273,
                     _9274 };
    assign _9276 = _9275 < _8771;
    assign _9277 = ~ _9276;
    assign _9265 = _8768[8:8];
    assign _9262 = _9257 - _8771;
    assign _9263 = _9259 ? _9262 : _9257;
    assign _9264 = _9263[62:0];
    assign _9266 = { _9264,
                     _9265 };
    assign _9267 = _9266 < _8771;
    assign _9268 = ~ _9267;
    assign _9256 = _8768[9:9];
    assign _9253 = _9248 - _8771;
    assign _9254 = _9250 ? _9253 : _9248;
    assign _9255 = _9254[62:0];
    assign _9257 = { _9255,
                     _9256 };
    assign _9258 = _9257 < _8771;
    assign _9259 = ~ _9258;
    assign _9247 = _8768[10:10];
    assign _9244 = _9239 - _8771;
    assign _9245 = _9241 ? _9244 : _9239;
    assign _9246 = _9245[62:0];
    assign _9248 = { _9246,
                     _9247 };
    assign _9249 = _9248 < _8771;
    assign _9250 = ~ _9249;
    assign _9238 = _8768[11:11];
    assign _9235 = _9230 - _8771;
    assign _9236 = _9232 ? _9235 : _9230;
    assign _9237 = _9236[62:0];
    assign _9239 = { _9237,
                     _9238 };
    assign _9240 = _9239 < _8771;
    assign _9241 = ~ _9240;
    assign _9229 = _8768[12:12];
    assign _9226 = _9221 - _8771;
    assign _9227 = _9223 ? _9226 : _9221;
    assign _9228 = _9227[62:0];
    assign _9230 = { _9228,
                     _9229 };
    assign _9231 = _9230 < _8771;
    assign _9232 = ~ _9231;
    assign _9220 = _8768[13:13];
    assign _9217 = _9212 - _8771;
    assign _9218 = _9214 ? _9217 : _9212;
    assign _9219 = _9218[62:0];
    assign _9221 = { _9219,
                     _9220 };
    assign _9222 = _9221 < _8771;
    assign _9223 = ~ _9222;
    assign _9211 = _8768[14:14];
    assign _9208 = _9203 - _8771;
    assign _9209 = _9205 ? _9208 : _9203;
    assign _9210 = _9209[62:0];
    assign _9212 = { _9210,
                     _9211 };
    assign _9213 = _9212 < _8771;
    assign _9214 = ~ _9213;
    assign _9202 = _8768[15:15];
    assign _9199 = _9194 - _8771;
    assign _9200 = _9196 ? _9199 : _9194;
    assign _9201 = _9200[62:0];
    assign _9203 = { _9201,
                     _9202 };
    assign _9204 = _9203 < _8771;
    assign _9205 = ~ _9204;
    assign _9193 = _8768[16:16];
    assign _9190 = _9185 - _8771;
    assign _9191 = _9187 ? _9190 : _9185;
    assign _9192 = _9191[62:0];
    assign _9194 = { _9192,
                     _9193 };
    assign _9195 = _9194 < _8771;
    assign _9196 = ~ _9195;
    assign _9184 = _8768[17:17];
    assign _9181 = _9176 - _8771;
    assign _9182 = _9178 ? _9181 : _9176;
    assign _9183 = _9182[62:0];
    assign _9185 = { _9183,
                     _9184 };
    assign _9186 = _9185 < _8771;
    assign _9187 = ~ _9186;
    assign _9175 = _8768[18:18];
    assign _9172 = _9167 - _8771;
    assign _9173 = _9169 ? _9172 : _9167;
    assign _9174 = _9173[62:0];
    assign _9176 = { _9174,
                     _9175 };
    assign _9177 = _9176 < _8771;
    assign _9178 = ~ _9177;
    assign _9166 = _8768[19:19];
    assign _9163 = _9158 - _8771;
    assign _9164 = _9160 ? _9163 : _9158;
    assign _9165 = _9164[62:0];
    assign _9167 = { _9165,
                     _9166 };
    assign _9168 = _9167 < _8771;
    assign _9169 = ~ _9168;
    assign _9157 = _8768[20:20];
    assign _9154 = _9149 - _8771;
    assign _9155 = _9151 ? _9154 : _9149;
    assign _9156 = _9155[62:0];
    assign _9158 = { _9156,
                     _9157 };
    assign _9159 = _9158 < _8771;
    assign _9160 = ~ _9159;
    assign _9148 = _8768[21:21];
    assign _9145 = _9140 - _8771;
    assign _9146 = _9142 ? _9145 : _9140;
    assign _9147 = _9146[62:0];
    assign _9149 = { _9147,
                     _9148 };
    assign _9150 = _9149 < _8771;
    assign _9151 = ~ _9150;
    assign _9139 = _8768[22:22];
    assign _9136 = _9131 - _8771;
    assign _9137 = _9133 ? _9136 : _9131;
    assign _9138 = _9137[62:0];
    assign _9140 = { _9138,
                     _9139 };
    assign _9141 = _9140 < _8771;
    assign _9142 = ~ _9141;
    assign _9130 = _8768[23:23];
    assign _9127 = _9122 - _8771;
    assign _9128 = _9124 ? _9127 : _9122;
    assign _9129 = _9128[62:0];
    assign _9131 = { _9129,
                     _9130 };
    assign _9132 = _9131 < _8771;
    assign _9133 = ~ _9132;
    assign _9121 = _8768[24:24];
    assign _9118 = _9113 - _8771;
    assign _9119 = _9115 ? _9118 : _9113;
    assign _9120 = _9119[62:0];
    assign _9122 = { _9120,
                     _9121 };
    assign _9123 = _9122 < _8771;
    assign _9124 = ~ _9123;
    assign _9112 = _8768[25:25];
    assign _9109 = _9104 - _8771;
    assign _9110 = _9106 ? _9109 : _9104;
    assign _9111 = _9110[62:0];
    assign _9113 = { _9111,
                     _9112 };
    assign _9114 = _9113 < _8771;
    assign _9115 = ~ _9114;
    assign _9103 = _8768[26:26];
    assign _9100 = _9095 - _8771;
    assign _9101 = _9097 ? _9100 : _9095;
    assign _9102 = _9101[62:0];
    assign _9104 = { _9102,
                     _9103 };
    assign _9105 = _9104 < _8771;
    assign _9106 = ~ _9105;
    assign _9094 = _8768[27:27];
    assign _9091 = _9086 - _8771;
    assign _9092 = _9088 ? _9091 : _9086;
    assign _9093 = _9092[62:0];
    assign _9095 = { _9093,
                     _9094 };
    assign _9096 = _9095 < _8771;
    assign _9097 = ~ _9096;
    assign _9085 = _8768[28:28];
    assign _9082 = _9077 - _8771;
    assign _9083 = _9079 ? _9082 : _9077;
    assign _9084 = _9083[62:0];
    assign _9086 = { _9084,
                     _9085 };
    assign _9087 = _9086 < _8771;
    assign _9088 = ~ _9087;
    assign _9076 = _8768[29:29];
    assign _9073 = _9068 - _8771;
    assign _9074 = _9070 ? _9073 : _9068;
    assign _9075 = _9074[62:0];
    assign _9077 = { _9075,
                     _9076 };
    assign _9078 = _9077 < _8771;
    assign _9079 = ~ _9078;
    assign _9067 = _8768[30:30];
    assign _9064 = _9059 - _8771;
    assign _9065 = _9061 ? _9064 : _9059;
    assign _9066 = _9065[62:0];
    assign _9068 = { _9066,
                     _9067 };
    assign _9069 = _9068 < _8771;
    assign _9070 = ~ _9069;
    assign _9058 = _8768[31:31];
    assign _9055 = _9050 - _8771;
    assign _9056 = _9052 ? _9055 : _9050;
    assign _9057 = _9056[62:0];
    assign _9059 = { _9057,
                     _9058 };
    assign _9060 = _9059 < _8771;
    assign _9061 = ~ _9060;
    assign _9049 = _8768[32:32];
    assign _9046 = _9041 - _8771;
    assign _9047 = _9043 ? _9046 : _9041;
    assign _9048 = _9047[62:0];
    assign _9050 = { _9048,
                     _9049 };
    assign _9051 = _9050 < _8771;
    assign _9052 = ~ _9051;
    assign _9040 = _8768[33:33];
    assign _9037 = _9032 - _8771;
    assign _9038 = _9034 ? _9037 : _9032;
    assign _9039 = _9038[62:0];
    assign _9041 = { _9039,
                     _9040 };
    assign _9042 = _9041 < _8771;
    assign _9043 = ~ _9042;
    assign _9031 = _8768[34:34];
    assign _9028 = _9023 - _8771;
    assign _9029 = _9025 ? _9028 : _9023;
    assign _9030 = _9029[62:0];
    assign _9032 = { _9030,
                     _9031 };
    assign _9033 = _9032 < _8771;
    assign _9034 = ~ _9033;
    assign _9022 = _8768[35:35];
    assign _9019 = _9014 - _8771;
    assign _9020 = _9016 ? _9019 : _9014;
    assign _9021 = _9020[62:0];
    assign _9023 = { _9021,
                     _9022 };
    assign _9024 = _9023 < _8771;
    assign _9025 = ~ _9024;
    assign _9013 = _8768[36:36];
    assign _9010 = _9005 - _8771;
    assign _9011 = _9007 ? _9010 : _9005;
    assign _9012 = _9011[62:0];
    assign _9014 = { _9012,
                     _9013 };
    assign _9015 = _9014 < _8771;
    assign _9016 = ~ _9015;
    assign _9004 = _8768[37:37];
    assign _9001 = _8996 - _8771;
    assign _9002 = _8998 ? _9001 : _8996;
    assign _9003 = _9002[62:0];
    assign _9005 = { _9003,
                     _9004 };
    assign _9006 = _9005 < _8771;
    assign _9007 = ~ _9006;
    assign _8995 = _8768[38:38];
    assign _8992 = _8987 - _8771;
    assign _8993 = _8989 ? _8992 : _8987;
    assign _8994 = _8993[62:0];
    assign _8996 = { _8994,
                     _8995 };
    assign _8997 = _8996 < _8771;
    assign _8998 = ~ _8997;
    assign _8986 = _8768[39:39];
    assign _8983 = _8978 - _8771;
    assign _8984 = _8980 ? _8983 : _8978;
    assign _8985 = _8984[62:0];
    assign _8987 = { _8985,
                     _8986 };
    assign _8988 = _8987 < _8771;
    assign _8989 = ~ _8988;
    assign _8977 = _8768[40:40];
    assign _8974 = _8969 - _8771;
    assign _8975 = _8971 ? _8974 : _8969;
    assign _8976 = _8975[62:0];
    assign _8978 = { _8976,
                     _8977 };
    assign _8979 = _8978 < _8771;
    assign _8980 = ~ _8979;
    assign _8968 = _8768[41:41];
    assign _8965 = _8960 - _8771;
    assign _8966 = _8962 ? _8965 : _8960;
    assign _8967 = _8966[62:0];
    assign _8969 = { _8967,
                     _8968 };
    assign _8970 = _8969 < _8771;
    assign _8971 = ~ _8970;
    assign _8959 = _8768[42:42];
    assign _8956 = _8951 - _8771;
    assign _8957 = _8953 ? _8956 : _8951;
    assign _8958 = _8957[62:0];
    assign _8960 = { _8958,
                     _8959 };
    assign _8961 = _8960 < _8771;
    assign _8962 = ~ _8961;
    assign _8950 = _8768[43:43];
    assign _8947 = _8942 - _8771;
    assign _8948 = _8944 ? _8947 : _8942;
    assign _8949 = _8948[62:0];
    assign _8951 = { _8949,
                     _8950 };
    assign _8952 = _8951 < _8771;
    assign _8953 = ~ _8952;
    assign _8941 = _8768[44:44];
    assign _8938 = _8933 - _8771;
    assign _8939 = _8935 ? _8938 : _8933;
    assign _8940 = _8939[62:0];
    assign _8942 = { _8940,
                     _8941 };
    assign _8943 = _8942 < _8771;
    assign _8944 = ~ _8943;
    assign _8932 = _8768[45:45];
    assign _8929 = _8924 - _8771;
    assign _8930 = _8926 ? _8929 : _8924;
    assign _8931 = _8930[62:0];
    assign _8933 = { _8931,
                     _8932 };
    assign _8934 = _8933 < _8771;
    assign _8935 = ~ _8934;
    assign _8923 = _8768[46:46];
    assign _8920 = _8915 - _8771;
    assign _8921 = _8917 ? _8920 : _8915;
    assign _8922 = _8921[62:0];
    assign _8924 = { _8922,
                     _8923 };
    assign _8925 = _8924 < _8771;
    assign _8926 = ~ _8925;
    assign _8914 = _8768[47:47];
    assign _8911 = _8906 - _8771;
    assign _8912 = _8908 ? _8911 : _8906;
    assign _8913 = _8912[62:0];
    assign _8915 = { _8913,
                     _8914 };
    assign _8916 = _8915 < _8771;
    assign _8917 = ~ _8916;
    assign _8905 = _8768[48:48];
    assign _8902 = _8897 - _8771;
    assign _8903 = _8899 ? _8902 : _8897;
    assign _8904 = _8903[62:0];
    assign _8906 = { _8904,
                     _8905 };
    assign _8907 = _8906 < _8771;
    assign _8908 = ~ _8907;
    assign _8896 = _8768[49:49];
    assign _8893 = _8888 - _8771;
    assign _8894 = _8890 ? _8893 : _8888;
    assign _8895 = _8894[62:0];
    assign _8897 = { _8895,
                     _8896 };
    assign _8898 = _8897 < _8771;
    assign _8899 = ~ _8898;
    assign _8887 = _8768[50:50];
    assign _8884 = _8879 - _8771;
    assign _8885 = _8881 ? _8884 : _8879;
    assign _8886 = _8885[62:0];
    assign _8888 = { _8886,
                     _8887 };
    assign _8889 = _8888 < _8771;
    assign _8890 = ~ _8889;
    assign _8878 = _8768[51:51];
    assign _8875 = _8870 - _8771;
    assign _8876 = _8872 ? _8875 : _8870;
    assign _8877 = _8876[62:0];
    assign _8879 = { _8877,
                     _8878 };
    assign _8880 = _8879 < _8771;
    assign _8881 = ~ _8880;
    assign _8869 = _8768[52:52];
    assign _8866 = _8861 - _8771;
    assign _8867 = _8863 ? _8866 : _8861;
    assign _8868 = _8867[62:0];
    assign _8870 = { _8868,
                     _8869 };
    assign _8871 = _8870 < _8771;
    assign _8872 = ~ _8871;
    assign _8860 = _8768[53:53];
    assign _8857 = _8852 - _8771;
    assign _8858 = _8854 ? _8857 : _8852;
    assign _8859 = _8858[62:0];
    assign _8861 = { _8859,
                     _8860 };
    assign _8862 = _8861 < _8771;
    assign _8863 = ~ _8862;
    assign _8851 = _8768[54:54];
    assign _8848 = _8843 - _8771;
    assign _8849 = _8845 ? _8848 : _8843;
    assign _8850 = _8849[62:0];
    assign _8852 = { _8850,
                     _8851 };
    assign _8853 = _8852 < _8771;
    assign _8854 = ~ _8853;
    assign _8842 = _8768[55:55];
    assign _8839 = _8834 - _8771;
    assign _8840 = _8836 ? _8839 : _8834;
    assign _8841 = _8840[62:0];
    assign _8843 = { _8841,
                     _8842 };
    assign _8844 = _8843 < _8771;
    assign _8845 = ~ _8844;
    assign _8833 = _8768[56:56];
    assign _8830 = _8825 - _8771;
    assign _8831 = _8827 ? _8830 : _8825;
    assign _8832 = _8831[62:0];
    assign _8834 = { _8832,
                     _8833 };
    assign _8835 = _8834 < _8771;
    assign _8836 = ~ _8835;
    assign _8824 = _8768[57:57];
    assign _8821 = _8816 - _8771;
    assign _8822 = _8818 ? _8821 : _8816;
    assign _8823 = _8822[62:0];
    assign _8825 = { _8823,
                     _8824 };
    assign _8826 = _8825 < _8771;
    assign _8827 = ~ _8826;
    assign _8815 = _8768[58:58];
    assign _8812 = _8807 - _8771;
    assign _8813 = _8809 ? _8812 : _8807;
    assign _8814 = _8813[62:0];
    assign _8816 = { _8814,
                     _8815 };
    assign _8817 = _8816 < _8771;
    assign _8818 = ~ _8817;
    assign _8806 = _8768[59:59];
    assign _8803 = _8798 - _8771;
    assign _8804 = _8800 ? _8803 : _8798;
    assign _8805 = _8804[62:0];
    assign _8807 = { _8805,
                     _8806 };
    assign _8808 = _8807 < _8771;
    assign _8809 = ~ _8808;
    assign _8797 = _8768[60:60];
    assign _8794 = _8789 - _8771;
    assign _8795 = _8791 ? _8794 : _8789;
    assign _8796 = _8795[62:0];
    assign _8798 = { _8796,
                     _8797 };
    assign _8799 = _8798 < _8771;
    assign _8800 = ~ _8799;
    assign _8788 = _8768[61:61];
    assign _8785 = _8780 - _8771;
    assign _8786 = _8782 ? _8785 : _8780;
    assign _8787 = _8786[62:0];
    assign _8789 = { _8787,
                     _8788 };
    assign _8790 = _8789 < _8771;
    assign _8791 = ~ _8790;
    assign _8779 = _8768[62:62];
    assign _8776 = _8770 - _8771;
    assign _8777 = _8773 ? _8776 : _8770;
    assign _8778 = _8777[62:0];
    assign _8780 = { _8778,
                     _8779 };
    assign _8781 = _8780 < _8771;
    assign _8782 = ~ _8781;
    assign _8771 = 64'b0000000000000000000000000000000000000000000000000000000001101111;
    assign _8767 = 64'b0000000000000000000000000000000000000000000000000000000001101110;
    assign _8768 = _3 + _8767;
    assign _8769 = _8768[63:63];
    assign _8770 = { _22185,
                     _8769 };
    assign _8772 = _8770 < _8771;
    assign _8773 = ~ _8772;
    assign _8774 = { _22185,
                     _8773 };
    assign _8775 = _8774[62:0];
    assign _8783 = { _8775,
                     _8782 };
    assign _8784 = _8783[62:0];
    assign _8792 = { _8784,
                     _8791 };
    assign _8793 = _8792[62:0];
    assign _8801 = { _8793,
                     _8800 };
    assign _8802 = _8801[62:0];
    assign _8810 = { _8802,
                     _8809 };
    assign _8811 = _8810[62:0];
    assign _8819 = { _8811,
                     _8818 };
    assign _8820 = _8819[62:0];
    assign _8828 = { _8820,
                     _8827 };
    assign _8829 = _8828[62:0];
    assign _8837 = { _8829,
                     _8836 };
    assign _8838 = _8837[62:0];
    assign _8846 = { _8838,
                     _8845 };
    assign _8847 = _8846[62:0];
    assign _8855 = { _8847,
                     _8854 };
    assign _8856 = _8855[62:0];
    assign _8864 = { _8856,
                     _8863 };
    assign _8865 = _8864[62:0];
    assign _8873 = { _8865,
                     _8872 };
    assign _8874 = _8873[62:0];
    assign _8882 = { _8874,
                     _8881 };
    assign _8883 = _8882[62:0];
    assign _8891 = { _8883,
                     _8890 };
    assign _8892 = _8891[62:0];
    assign _8900 = { _8892,
                     _8899 };
    assign _8901 = _8900[62:0];
    assign _8909 = { _8901,
                     _8908 };
    assign _8910 = _8909[62:0];
    assign _8918 = { _8910,
                     _8917 };
    assign _8919 = _8918[62:0];
    assign _8927 = { _8919,
                     _8926 };
    assign _8928 = _8927[62:0];
    assign _8936 = { _8928,
                     _8935 };
    assign _8937 = _8936[62:0];
    assign _8945 = { _8937,
                     _8944 };
    assign _8946 = _8945[62:0];
    assign _8954 = { _8946,
                     _8953 };
    assign _8955 = _8954[62:0];
    assign _8963 = { _8955,
                     _8962 };
    assign _8964 = _8963[62:0];
    assign _8972 = { _8964,
                     _8971 };
    assign _8973 = _8972[62:0];
    assign _8981 = { _8973,
                     _8980 };
    assign _8982 = _8981[62:0];
    assign _8990 = { _8982,
                     _8989 };
    assign _8991 = _8990[62:0];
    assign _8999 = { _8991,
                     _8998 };
    assign _9000 = _8999[62:0];
    assign _9008 = { _9000,
                     _9007 };
    assign _9009 = _9008[62:0];
    assign _9017 = { _9009,
                     _9016 };
    assign _9018 = _9017[62:0];
    assign _9026 = { _9018,
                     _9025 };
    assign _9027 = _9026[62:0];
    assign _9035 = { _9027,
                     _9034 };
    assign _9036 = _9035[62:0];
    assign _9044 = { _9036,
                     _9043 };
    assign _9045 = _9044[62:0];
    assign _9053 = { _9045,
                     _9052 };
    assign _9054 = _9053[62:0];
    assign _9062 = { _9054,
                     _9061 };
    assign _9063 = _9062[62:0];
    assign _9071 = { _9063,
                     _9070 };
    assign _9072 = _9071[62:0];
    assign _9080 = { _9072,
                     _9079 };
    assign _9081 = _9080[62:0];
    assign _9089 = { _9081,
                     _9088 };
    assign _9090 = _9089[62:0];
    assign _9098 = { _9090,
                     _9097 };
    assign _9099 = _9098[62:0];
    assign _9107 = { _9099,
                     _9106 };
    assign _9108 = _9107[62:0];
    assign _9116 = { _9108,
                     _9115 };
    assign _9117 = _9116[62:0];
    assign _9125 = { _9117,
                     _9124 };
    assign _9126 = _9125[62:0];
    assign _9134 = { _9126,
                     _9133 };
    assign _9135 = _9134[62:0];
    assign _9143 = { _9135,
                     _9142 };
    assign _9144 = _9143[62:0];
    assign _9152 = { _9144,
                     _9151 };
    assign _9153 = _9152[62:0];
    assign _9161 = { _9153,
                     _9160 };
    assign _9162 = _9161[62:0];
    assign _9170 = { _9162,
                     _9169 };
    assign _9171 = _9170[62:0];
    assign _9179 = { _9171,
                     _9178 };
    assign _9180 = _9179[62:0];
    assign _9188 = { _9180,
                     _9187 };
    assign _9189 = _9188[62:0];
    assign _9197 = { _9189,
                     _9196 };
    assign _9198 = _9197[62:0];
    assign _9206 = { _9198,
                     _9205 };
    assign _9207 = _9206[62:0];
    assign _9215 = { _9207,
                     _9214 };
    assign _9216 = _9215[62:0];
    assign _9224 = { _9216,
                     _9223 };
    assign _9225 = _9224[62:0];
    assign _9233 = { _9225,
                     _9232 };
    assign _9234 = _9233[62:0];
    assign _9242 = { _9234,
                     _9241 };
    assign _9243 = _9242[62:0];
    assign _9251 = { _9243,
                     _9250 };
    assign _9252 = _9251[62:0];
    assign _9260 = { _9252,
                     _9259 };
    assign _9261 = _9260[62:0];
    assign _9269 = { _9261,
                     _9268 };
    assign _9270 = _9269[62:0];
    assign _9278 = { _9270,
                     _9277 };
    assign _9279 = _9278[62:0];
    assign _9287 = { _9279,
                     _9286 };
    assign _9288 = _9287[62:0];
    assign _9296 = { _9288,
                     _9295 };
    assign _9297 = _9296[62:0];
    assign _9305 = { _9297,
                     _9304 };
    assign _9306 = _9305[62:0];
    assign _9314 = { _9306,
                     _9313 };
    assign _9315 = _9314[62:0];
    assign _9323 = { _9315,
                     _9322 };
    assign _9324 = _9323[62:0];
    assign _9332 = { _9324,
                     _9331 };
    assign _9333 = _9332[62:0];
    assign _9341 = { _9333,
                     _9340 };
    assign _9342 = _9341 * _8771;
    assign _9343 = _9342[63:0];
    assign _9344 = _8771 < _9343;
    assign _9345 = _9344 ? _9343 : _8771;
    assign _8761 = 64'b0000000000000000000000000000000000000000000000000000001111100111;
    assign _8762 = _5 < _8761;
    assign _8763 = _8762 ? _5 : _8761;
    assign _9346 = _8763 < _9345;
    assign _9347 = ~ _9346;
    assign _10510 = _9347 ? _10509 : _21604;
    assign _12261 = _10510 + _12260;
    assign _14012 = _12261 + _14011;
    assign _15763 = _14012 + _15762;
    assign _17514 = _15763 + _17513;
    assign _19265 = _17514 + _19264;
    assign _19266 = _8760 + _19265;
    assign _22768 = _19266 - _22767;
    assign _8751 = _8182[0:0];
    assign _8748 = _8743 - _22192;
    assign _8749 = _8745 ? _8748 : _8743;
    assign _8750 = _8749[62:0];
    assign _8752 = { _8750,
                     _8751 };
    assign _8753 = _8752 < _22192;
    assign _8754 = ~ _8753;
    assign _8742 = _8182[1:1];
    assign _8739 = _8734 - _22192;
    assign _8740 = _8736 ? _8739 : _8734;
    assign _8741 = _8740[62:0];
    assign _8743 = { _8741,
                     _8742 };
    assign _8744 = _8743 < _22192;
    assign _8745 = ~ _8744;
    assign _8733 = _8182[2:2];
    assign _8730 = _8725 - _22192;
    assign _8731 = _8727 ? _8730 : _8725;
    assign _8732 = _8731[62:0];
    assign _8734 = { _8732,
                     _8733 };
    assign _8735 = _8734 < _22192;
    assign _8736 = ~ _8735;
    assign _8724 = _8182[3:3];
    assign _8721 = _8716 - _22192;
    assign _8722 = _8718 ? _8721 : _8716;
    assign _8723 = _8722[62:0];
    assign _8725 = { _8723,
                     _8724 };
    assign _8726 = _8725 < _22192;
    assign _8727 = ~ _8726;
    assign _8715 = _8182[4:4];
    assign _8712 = _8707 - _22192;
    assign _8713 = _8709 ? _8712 : _8707;
    assign _8714 = _8713[62:0];
    assign _8716 = { _8714,
                     _8715 };
    assign _8717 = _8716 < _22192;
    assign _8718 = ~ _8717;
    assign _8706 = _8182[5:5];
    assign _8703 = _8698 - _22192;
    assign _8704 = _8700 ? _8703 : _8698;
    assign _8705 = _8704[62:0];
    assign _8707 = { _8705,
                     _8706 };
    assign _8708 = _8707 < _22192;
    assign _8709 = ~ _8708;
    assign _8697 = _8182[6:6];
    assign _8694 = _8689 - _22192;
    assign _8695 = _8691 ? _8694 : _8689;
    assign _8696 = _8695[62:0];
    assign _8698 = { _8696,
                     _8697 };
    assign _8699 = _8698 < _22192;
    assign _8700 = ~ _8699;
    assign _8688 = _8182[7:7];
    assign _8685 = _8680 - _22192;
    assign _8686 = _8682 ? _8685 : _8680;
    assign _8687 = _8686[62:0];
    assign _8689 = { _8687,
                     _8688 };
    assign _8690 = _8689 < _22192;
    assign _8691 = ~ _8690;
    assign _8679 = _8182[8:8];
    assign _8676 = _8671 - _22192;
    assign _8677 = _8673 ? _8676 : _8671;
    assign _8678 = _8677[62:0];
    assign _8680 = { _8678,
                     _8679 };
    assign _8681 = _8680 < _22192;
    assign _8682 = ~ _8681;
    assign _8670 = _8182[9:9];
    assign _8667 = _8662 - _22192;
    assign _8668 = _8664 ? _8667 : _8662;
    assign _8669 = _8668[62:0];
    assign _8671 = { _8669,
                     _8670 };
    assign _8672 = _8671 < _22192;
    assign _8673 = ~ _8672;
    assign _8661 = _8182[10:10];
    assign _8658 = _8653 - _22192;
    assign _8659 = _8655 ? _8658 : _8653;
    assign _8660 = _8659[62:0];
    assign _8662 = { _8660,
                     _8661 };
    assign _8663 = _8662 < _22192;
    assign _8664 = ~ _8663;
    assign _8652 = _8182[11:11];
    assign _8649 = _8644 - _22192;
    assign _8650 = _8646 ? _8649 : _8644;
    assign _8651 = _8650[62:0];
    assign _8653 = { _8651,
                     _8652 };
    assign _8654 = _8653 < _22192;
    assign _8655 = ~ _8654;
    assign _8643 = _8182[12:12];
    assign _8640 = _8635 - _22192;
    assign _8641 = _8637 ? _8640 : _8635;
    assign _8642 = _8641[62:0];
    assign _8644 = { _8642,
                     _8643 };
    assign _8645 = _8644 < _22192;
    assign _8646 = ~ _8645;
    assign _8634 = _8182[13:13];
    assign _8631 = _8626 - _22192;
    assign _8632 = _8628 ? _8631 : _8626;
    assign _8633 = _8632[62:0];
    assign _8635 = { _8633,
                     _8634 };
    assign _8636 = _8635 < _22192;
    assign _8637 = ~ _8636;
    assign _8625 = _8182[14:14];
    assign _8622 = _8617 - _22192;
    assign _8623 = _8619 ? _8622 : _8617;
    assign _8624 = _8623[62:0];
    assign _8626 = { _8624,
                     _8625 };
    assign _8627 = _8626 < _22192;
    assign _8628 = ~ _8627;
    assign _8616 = _8182[15:15];
    assign _8613 = _8608 - _22192;
    assign _8614 = _8610 ? _8613 : _8608;
    assign _8615 = _8614[62:0];
    assign _8617 = { _8615,
                     _8616 };
    assign _8618 = _8617 < _22192;
    assign _8619 = ~ _8618;
    assign _8607 = _8182[16:16];
    assign _8604 = _8599 - _22192;
    assign _8605 = _8601 ? _8604 : _8599;
    assign _8606 = _8605[62:0];
    assign _8608 = { _8606,
                     _8607 };
    assign _8609 = _8608 < _22192;
    assign _8610 = ~ _8609;
    assign _8598 = _8182[17:17];
    assign _8595 = _8590 - _22192;
    assign _8596 = _8592 ? _8595 : _8590;
    assign _8597 = _8596[62:0];
    assign _8599 = { _8597,
                     _8598 };
    assign _8600 = _8599 < _22192;
    assign _8601 = ~ _8600;
    assign _8589 = _8182[18:18];
    assign _8586 = _8581 - _22192;
    assign _8587 = _8583 ? _8586 : _8581;
    assign _8588 = _8587[62:0];
    assign _8590 = { _8588,
                     _8589 };
    assign _8591 = _8590 < _22192;
    assign _8592 = ~ _8591;
    assign _8580 = _8182[19:19];
    assign _8577 = _8572 - _22192;
    assign _8578 = _8574 ? _8577 : _8572;
    assign _8579 = _8578[62:0];
    assign _8581 = { _8579,
                     _8580 };
    assign _8582 = _8581 < _22192;
    assign _8583 = ~ _8582;
    assign _8571 = _8182[20:20];
    assign _8568 = _8563 - _22192;
    assign _8569 = _8565 ? _8568 : _8563;
    assign _8570 = _8569[62:0];
    assign _8572 = { _8570,
                     _8571 };
    assign _8573 = _8572 < _22192;
    assign _8574 = ~ _8573;
    assign _8562 = _8182[21:21];
    assign _8559 = _8554 - _22192;
    assign _8560 = _8556 ? _8559 : _8554;
    assign _8561 = _8560[62:0];
    assign _8563 = { _8561,
                     _8562 };
    assign _8564 = _8563 < _22192;
    assign _8565 = ~ _8564;
    assign _8553 = _8182[22:22];
    assign _8550 = _8545 - _22192;
    assign _8551 = _8547 ? _8550 : _8545;
    assign _8552 = _8551[62:0];
    assign _8554 = { _8552,
                     _8553 };
    assign _8555 = _8554 < _22192;
    assign _8556 = ~ _8555;
    assign _8544 = _8182[23:23];
    assign _8541 = _8536 - _22192;
    assign _8542 = _8538 ? _8541 : _8536;
    assign _8543 = _8542[62:0];
    assign _8545 = { _8543,
                     _8544 };
    assign _8546 = _8545 < _22192;
    assign _8547 = ~ _8546;
    assign _8535 = _8182[24:24];
    assign _8532 = _8527 - _22192;
    assign _8533 = _8529 ? _8532 : _8527;
    assign _8534 = _8533[62:0];
    assign _8536 = { _8534,
                     _8535 };
    assign _8537 = _8536 < _22192;
    assign _8538 = ~ _8537;
    assign _8526 = _8182[25:25];
    assign _8523 = _8518 - _22192;
    assign _8524 = _8520 ? _8523 : _8518;
    assign _8525 = _8524[62:0];
    assign _8527 = { _8525,
                     _8526 };
    assign _8528 = _8527 < _22192;
    assign _8529 = ~ _8528;
    assign _8517 = _8182[26:26];
    assign _8514 = _8509 - _22192;
    assign _8515 = _8511 ? _8514 : _8509;
    assign _8516 = _8515[62:0];
    assign _8518 = { _8516,
                     _8517 };
    assign _8519 = _8518 < _22192;
    assign _8520 = ~ _8519;
    assign _8508 = _8182[27:27];
    assign _8505 = _8500 - _22192;
    assign _8506 = _8502 ? _8505 : _8500;
    assign _8507 = _8506[62:0];
    assign _8509 = { _8507,
                     _8508 };
    assign _8510 = _8509 < _22192;
    assign _8511 = ~ _8510;
    assign _8499 = _8182[28:28];
    assign _8496 = _8491 - _22192;
    assign _8497 = _8493 ? _8496 : _8491;
    assign _8498 = _8497[62:0];
    assign _8500 = { _8498,
                     _8499 };
    assign _8501 = _8500 < _22192;
    assign _8502 = ~ _8501;
    assign _8490 = _8182[29:29];
    assign _8487 = _8482 - _22192;
    assign _8488 = _8484 ? _8487 : _8482;
    assign _8489 = _8488[62:0];
    assign _8491 = { _8489,
                     _8490 };
    assign _8492 = _8491 < _22192;
    assign _8493 = ~ _8492;
    assign _8481 = _8182[30:30];
    assign _8478 = _8473 - _22192;
    assign _8479 = _8475 ? _8478 : _8473;
    assign _8480 = _8479[62:0];
    assign _8482 = { _8480,
                     _8481 };
    assign _8483 = _8482 < _22192;
    assign _8484 = ~ _8483;
    assign _8472 = _8182[31:31];
    assign _8469 = _8464 - _22192;
    assign _8470 = _8466 ? _8469 : _8464;
    assign _8471 = _8470[62:0];
    assign _8473 = { _8471,
                     _8472 };
    assign _8474 = _8473 < _22192;
    assign _8475 = ~ _8474;
    assign _8463 = _8182[32:32];
    assign _8460 = _8455 - _22192;
    assign _8461 = _8457 ? _8460 : _8455;
    assign _8462 = _8461[62:0];
    assign _8464 = { _8462,
                     _8463 };
    assign _8465 = _8464 < _22192;
    assign _8466 = ~ _8465;
    assign _8454 = _8182[33:33];
    assign _8451 = _8446 - _22192;
    assign _8452 = _8448 ? _8451 : _8446;
    assign _8453 = _8452[62:0];
    assign _8455 = { _8453,
                     _8454 };
    assign _8456 = _8455 < _22192;
    assign _8457 = ~ _8456;
    assign _8445 = _8182[34:34];
    assign _8442 = _8437 - _22192;
    assign _8443 = _8439 ? _8442 : _8437;
    assign _8444 = _8443[62:0];
    assign _8446 = { _8444,
                     _8445 };
    assign _8447 = _8446 < _22192;
    assign _8448 = ~ _8447;
    assign _8436 = _8182[35:35];
    assign _8433 = _8428 - _22192;
    assign _8434 = _8430 ? _8433 : _8428;
    assign _8435 = _8434[62:0];
    assign _8437 = { _8435,
                     _8436 };
    assign _8438 = _8437 < _22192;
    assign _8439 = ~ _8438;
    assign _8427 = _8182[36:36];
    assign _8424 = _8419 - _22192;
    assign _8425 = _8421 ? _8424 : _8419;
    assign _8426 = _8425[62:0];
    assign _8428 = { _8426,
                     _8427 };
    assign _8429 = _8428 < _22192;
    assign _8430 = ~ _8429;
    assign _8418 = _8182[37:37];
    assign _8415 = _8410 - _22192;
    assign _8416 = _8412 ? _8415 : _8410;
    assign _8417 = _8416[62:0];
    assign _8419 = { _8417,
                     _8418 };
    assign _8420 = _8419 < _22192;
    assign _8421 = ~ _8420;
    assign _8409 = _8182[38:38];
    assign _8406 = _8401 - _22192;
    assign _8407 = _8403 ? _8406 : _8401;
    assign _8408 = _8407[62:0];
    assign _8410 = { _8408,
                     _8409 };
    assign _8411 = _8410 < _22192;
    assign _8412 = ~ _8411;
    assign _8400 = _8182[39:39];
    assign _8397 = _8392 - _22192;
    assign _8398 = _8394 ? _8397 : _8392;
    assign _8399 = _8398[62:0];
    assign _8401 = { _8399,
                     _8400 };
    assign _8402 = _8401 < _22192;
    assign _8403 = ~ _8402;
    assign _8391 = _8182[40:40];
    assign _8388 = _8383 - _22192;
    assign _8389 = _8385 ? _8388 : _8383;
    assign _8390 = _8389[62:0];
    assign _8392 = { _8390,
                     _8391 };
    assign _8393 = _8392 < _22192;
    assign _8394 = ~ _8393;
    assign _8382 = _8182[41:41];
    assign _8379 = _8374 - _22192;
    assign _8380 = _8376 ? _8379 : _8374;
    assign _8381 = _8380[62:0];
    assign _8383 = { _8381,
                     _8382 };
    assign _8384 = _8383 < _22192;
    assign _8385 = ~ _8384;
    assign _8373 = _8182[42:42];
    assign _8370 = _8365 - _22192;
    assign _8371 = _8367 ? _8370 : _8365;
    assign _8372 = _8371[62:0];
    assign _8374 = { _8372,
                     _8373 };
    assign _8375 = _8374 < _22192;
    assign _8376 = ~ _8375;
    assign _8364 = _8182[43:43];
    assign _8361 = _8356 - _22192;
    assign _8362 = _8358 ? _8361 : _8356;
    assign _8363 = _8362[62:0];
    assign _8365 = { _8363,
                     _8364 };
    assign _8366 = _8365 < _22192;
    assign _8367 = ~ _8366;
    assign _8355 = _8182[44:44];
    assign _8352 = _8347 - _22192;
    assign _8353 = _8349 ? _8352 : _8347;
    assign _8354 = _8353[62:0];
    assign _8356 = { _8354,
                     _8355 };
    assign _8357 = _8356 < _22192;
    assign _8358 = ~ _8357;
    assign _8346 = _8182[45:45];
    assign _8343 = _8338 - _22192;
    assign _8344 = _8340 ? _8343 : _8338;
    assign _8345 = _8344[62:0];
    assign _8347 = { _8345,
                     _8346 };
    assign _8348 = _8347 < _22192;
    assign _8349 = ~ _8348;
    assign _8337 = _8182[46:46];
    assign _8334 = _8329 - _22192;
    assign _8335 = _8331 ? _8334 : _8329;
    assign _8336 = _8335[62:0];
    assign _8338 = { _8336,
                     _8337 };
    assign _8339 = _8338 < _22192;
    assign _8340 = ~ _8339;
    assign _8328 = _8182[47:47];
    assign _8325 = _8320 - _22192;
    assign _8326 = _8322 ? _8325 : _8320;
    assign _8327 = _8326[62:0];
    assign _8329 = { _8327,
                     _8328 };
    assign _8330 = _8329 < _22192;
    assign _8331 = ~ _8330;
    assign _8319 = _8182[48:48];
    assign _8316 = _8311 - _22192;
    assign _8317 = _8313 ? _8316 : _8311;
    assign _8318 = _8317[62:0];
    assign _8320 = { _8318,
                     _8319 };
    assign _8321 = _8320 < _22192;
    assign _8322 = ~ _8321;
    assign _8310 = _8182[49:49];
    assign _8307 = _8302 - _22192;
    assign _8308 = _8304 ? _8307 : _8302;
    assign _8309 = _8308[62:0];
    assign _8311 = { _8309,
                     _8310 };
    assign _8312 = _8311 < _22192;
    assign _8313 = ~ _8312;
    assign _8301 = _8182[50:50];
    assign _8298 = _8293 - _22192;
    assign _8299 = _8295 ? _8298 : _8293;
    assign _8300 = _8299[62:0];
    assign _8302 = { _8300,
                     _8301 };
    assign _8303 = _8302 < _22192;
    assign _8304 = ~ _8303;
    assign _8292 = _8182[51:51];
    assign _8289 = _8284 - _22192;
    assign _8290 = _8286 ? _8289 : _8284;
    assign _8291 = _8290[62:0];
    assign _8293 = { _8291,
                     _8292 };
    assign _8294 = _8293 < _22192;
    assign _8295 = ~ _8294;
    assign _8283 = _8182[52:52];
    assign _8280 = _8275 - _22192;
    assign _8281 = _8277 ? _8280 : _8275;
    assign _8282 = _8281[62:0];
    assign _8284 = { _8282,
                     _8283 };
    assign _8285 = _8284 < _22192;
    assign _8286 = ~ _8285;
    assign _8274 = _8182[53:53];
    assign _8271 = _8266 - _22192;
    assign _8272 = _8268 ? _8271 : _8266;
    assign _8273 = _8272[62:0];
    assign _8275 = { _8273,
                     _8274 };
    assign _8276 = _8275 < _22192;
    assign _8277 = ~ _8276;
    assign _8265 = _8182[54:54];
    assign _8262 = _8257 - _22192;
    assign _8263 = _8259 ? _8262 : _8257;
    assign _8264 = _8263[62:0];
    assign _8266 = { _8264,
                     _8265 };
    assign _8267 = _8266 < _22192;
    assign _8268 = ~ _8267;
    assign _8256 = _8182[55:55];
    assign _8253 = _8248 - _22192;
    assign _8254 = _8250 ? _8253 : _8248;
    assign _8255 = _8254[62:0];
    assign _8257 = { _8255,
                     _8256 };
    assign _8258 = _8257 < _22192;
    assign _8259 = ~ _8258;
    assign _8247 = _8182[56:56];
    assign _8244 = _8239 - _22192;
    assign _8245 = _8241 ? _8244 : _8239;
    assign _8246 = _8245[62:0];
    assign _8248 = { _8246,
                     _8247 };
    assign _8249 = _8248 < _22192;
    assign _8250 = ~ _8249;
    assign _8238 = _8182[57:57];
    assign _8235 = _8230 - _22192;
    assign _8236 = _8232 ? _8235 : _8230;
    assign _8237 = _8236[62:0];
    assign _8239 = { _8237,
                     _8238 };
    assign _8240 = _8239 < _22192;
    assign _8241 = ~ _8240;
    assign _8229 = _8182[58:58];
    assign _8226 = _8221 - _22192;
    assign _8227 = _8223 ? _8226 : _8221;
    assign _8228 = _8227[62:0];
    assign _8230 = { _8228,
                     _8229 };
    assign _8231 = _8230 < _22192;
    assign _8232 = ~ _8231;
    assign _8220 = _8182[59:59];
    assign _8217 = _8212 - _22192;
    assign _8218 = _8214 ? _8217 : _8212;
    assign _8219 = _8218[62:0];
    assign _8221 = { _8219,
                     _8220 };
    assign _8222 = _8221 < _22192;
    assign _8223 = ~ _8222;
    assign _8211 = _8182[60:60];
    assign _8208 = _8203 - _22192;
    assign _8209 = _8205 ? _8208 : _8203;
    assign _8210 = _8209[62:0];
    assign _8212 = { _8210,
                     _8211 };
    assign _8213 = _8212 < _22192;
    assign _8214 = ~ _8213;
    assign _8202 = _8182[61:61];
    assign _8199 = _8194 - _22192;
    assign _8200 = _8196 ? _8199 : _8194;
    assign _8201 = _8200[62:0];
    assign _8203 = { _8201,
                     _8202 };
    assign _8204 = _8203 < _22192;
    assign _8205 = ~ _8204;
    assign _8193 = _8182[62:62];
    assign _8190 = _8184 - _22192;
    assign _8191 = _8187 ? _8190 : _8184;
    assign _8192 = _8191[62:0];
    assign _8194 = { _8192,
                     _8193 };
    assign _8195 = _8194 < _22192;
    assign _8196 = ~ _8195;
    assign _8180 = _8172 + _22186;
    assign _8181 = _8172 * _8180;
    assign _8182 = _8181[63:0];
    assign _8183 = _8182[63:63];
    assign _8184 = { _22185,
                     _8183 };
    assign _8186 = _8184 < _22192;
    assign _8187 = ~ _8186;
    assign _8188 = { _22185,
                     _8187 };
    assign _8189 = _8188[62:0];
    assign _8197 = { _8189,
                     _8196 };
    assign _8198 = _8197[62:0];
    assign _8206 = { _8198,
                     _8205 };
    assign _8207 = _8206[62:0];
    assign _8215 = { _8207,
                     _8214 };
    assign _8216 = _8215[62:0];
    assign _8224 = { _8216,
                     _8223 };
    assign _8225 = _8224[62:0];
    assign _8233 = { _8225,
                     _8232 };
    assign _8234 = _8233[62:0];
    assign _8242 = { _8234,
                     _8241 };
    assign _8243 = _8242[62:0];
    assign _8251 = { _8243,
                     _8250 };
    assign _8252 = _8251[62:0];
    assign _8260 = { _8252,
                     _8259 };
    assign _8261 = _8260[62:0];
    assign _8269 = { _8261,
                     _8268 };
    assign _8270 = _8269[62:0];
    assign _8278 = { _8270,
                     _8277 };
    assign _8279 = _8278[62:0];
    assign _8287 = { _8279,
                     _8286 };
    assign _8288 = _8287[62:0];
    assign _8296 = { _8288,
                     _8295 };
    assign _8297 = _8296[62:0];
    assign _8305 = { _8297,
                     _8304 };
    assign _8306 = _8305[62:0];
    assign _8314 = { _8306,
                     _8313 };
    assign _8315 = _8314[62:0];
    assign _8323 = { _8315,
                     _8322 };
    assign _8324 = _8323[62:0];
    assign _8332 = { _8324,
                     _8331 };
    assign _8333 = _8332[62:0];
    assign _8341 = { _8333,
                     _8340 };
    assign _8342 = _8341[62:0];
    assign _8350 = { _8342,
                     _8349 };
    assign _8351 = _8350[62:0];
    assign _8359 = { _8351,
                     _8358 };
    assign _8360 = _8359[62:0];
    assign _8368 = { _8360,
                     _8367 };
    assign _8369 = _8368[62:0];
    assign _8377 = { _8369,
                     _8376 };
    assign _8378 = _8377[62:0];
    assign _8386 = { _8378,
                     _8385 };
    assign _8387 = _8386[62:0];
    assign _8395 = { _8387,
                     _8394 };
    assign _8396 = _8395[62:0];
    assign _8404 = { _8396,
                     _8403 };
    assign _8405 = _8404[62:0];
    assign _8413 = { _8405,
                     _8412 };
    assign _8414 = _8413[62:0];
    assign _8422 = { _8414,
                     _8421 };
    assign _8423 = _8422[62:0];
    assign _8431 = { _8423,
                     _8430 };
    assign _8432 = _8431[62:0];
    assign _8440 = { _8432,
                     _8439 };
    assign _8441 = _8440[62:0];
    assign _8449 = { _8441,
                     _8448 };
    assign _8450 = _8449[62:0];
    assign _8458 = { _8450,
                     _8457 };
    assign _8459 = _8458[62:0];
    assign _8467 = { _8459,
                     _8466 };
    assign _8468 = _8467[62:0];
    assign _8476 = { _8468,
                     _8475 };
    assign _8477 = _8476[62:0];
    assign _8485 = { _8477,
                     _8484 };
    assign _8486 = _8485[62:0];
    assign _8494 = { _8486,
                     _8493 };
    assign _8495 = _8494[62:0];
    assign _8503 = { _8495,
                     _8502 };
    assign _8504 = _8503[62:0];
    assign _8512 = { _8504,
                     _8511 };
    assign _8513 = _8512[62:0];
    assign _8521 = { _8513,
                     _8520 };
    assign _8522 = _8521[62:0];
    assign _8530 = { _8522,
                     _8529 };
    assign _8531 = _8530[62:0];
    assign _8539 = { _8531,
                     _8538 };
    assign _8540 = _8539[62:0];
    assign _8548 = { _8540,
                     _8547 };
    assign _8549 = _8548[62:0];
    assign _8557 = { _8549,
                     _8556 };
    assign _8558 = _8557[62:0];
    assign _8566 = { _8558,
                     _8565 };
    assign _8567 = _8566[62:0];
    assign _8575 = { _8567,
                     _8574 };
    assign _8576 = _8575[62:0];
    assign _8584 = { _8576,
                     _8583 };
    assign _8585 = _8584[62:0];
    assign _8593 = { _8585,
                     _8592 };
    assign _8594 = _8593[62:0];
    assign _8602 = { _8594,
                     _8601 };
    assign _8603 = _8602[62:0];
    assign _8611 = { _8603,
                     _8610 };
    assign _8612 = _8611[62:0];
    assign _8620 = { _8612,
                     _8619 };
    assign _8621 = _8620[62:0];
    assign _8629 = { _8621,
                     _8628 };
    assign _8630 = _8629[62:0];
    assign _8638 = { _8630,
                     _8637 };
    assign _8639 = _8638[62:0];
    assign _8647 = { _8639,
                     _8646 };
    assign _8648 = _8647[62:0];
    assign _8656 = { _8648,
                     _8655 };
    assign _8657 = _8656[62:0];
    assign _8665 = { _8657,
                     _8664 };
    assign _8666 = _8665[62:0];
    assign _8674 = { _8666,
                     _8673 };
    assign _8675 = _8674[62:0];
    assign _8683 = { _8675,
                     _8682 };
    assign _8684 = _8683[62:0];
    assign _8692 = { _8684,
                     _8691 };
    assign _8693 = _8692[62:0];
    assign _8701 = { _8693,
                     _8700 };
    assign _8702 = _8701[62:0];
    assign _8710 = { _8702,
                     _8709 };
    assign _8711 = _8710[62:0];
    assign _8719 = { _8711,
                     _8718 };
    assign _8720 = _8719[62:0];
    assign _8728 = { _8720,
                     _8727 };
    assign _8729 = _8728[62:0];
    assign _8737 = { _8729,
                     _8736 };
    assign _8738 = _8737[62:0];
    assign _8746 = { _8738,
                     _8745 };
    assign _8747 = _8746[62:0];
    assign _8755 = { _8747,
                     _8754 };
    assign _8756 = _7020 * _8755;
    assign _8757 = _8756[63:0];
    assign _8168 = _7600[0:0];
    assign _8165 = _8160 - _7020;
    assign _8166 = _8162 ? _8165 : _8160;
    assign _8167 = _8166[62:0];
    assign _8169 = { _8167,
                     _8168 };
    assign _8170 = _8169 < _7020;
    assign _8171 = ~ _8170;
    assign _8159 = _7600[1:1];
    assign _8156 = _8151 - _7020;
    assign _8157 = _8153 ? _8156 : _8151;
    assign _8158 = _8157[62:0];
    assign _8160 = { _8158,
                     _8159 };
    assign _8161 = _8160 < _7020;
    assign _8162 = ~ _8161;
    assign _8150 = _7600[2:2];
    assign _8147 = _8142 - _7020;
    assign _8148 = _8144 ? _8147 : _8142;
    assign _8149 = _8148[62:0];
    assign _8151 = { _8149,
                     _8150 };
    assign _8152 = _8151 < _7020;
    assign _8153 = ~ _8152;
    assign _8141 = _7600[3:3];
    assign _8138 = _8133 - _7020;
    assign _8139 = _8135 ? _8138 : _8133;
    assign _8140 = _8139[62:0];
    assign _8142 = { _8140,
                     _8141 };
    assign _8143 = _8142 < _7020;
    assign _8144 = ~ _8143;
    assign _8132 = _7600[4:4];
    assign _8129 = _8124 - _7020;
    assign _8130 = _8126 ? _8129 : _8124;
    assign _8131 = _8130[62:0];
    assign _8133 = { _8131,
                     _8132 };
    assign _8134 = _8133 < _7020;
    assign _8135 = ~ _8134;
    assign _8123 = _7600[5:5];
    assign _8120 = _8115 - _7020;
    assign _8121 = _8117 ? _8120 : _8115;
    assign _8122 = _8121[62:0];
    assign _8124 = { _8122,
                     _8123 };
    assign _8125 = _8124 < _7020;
    assign _8126 = ~ _8125;
    assign _8114 = _7600[6:6];
    assign _8111 = _8106 - _7020;
    assign _8112 = _8108 ? _8111 : _8106;
    assign _8113 = _8112[62:0];
    assign _8115 = { _8113,
                     _8114 };
    assign _8116 = _8115 < _7020;
    assign _8117 = ~ _8116;
    assign _8105 = _7600[7:7];
    assign _8102 = _8097 - _7020;
    assign _8103 = _8099 ? _8102 : _8097;
    assign _8104 = _8103[62:0];
    assign _8106 = { _8104,
                     _8105 };
    assign _8107 = _8106 < _7020;
    assign _8108 = ~ _8107;
    assign _8096 = _7600[8:8];
    assign _8093 = _8088 - _7020;
    assign _8094 = _8090 ? _8093 : _8088;
    assign _8095 = _8094[62:0];
    assign _8097 = { _8095,
                     _8096 };
    assign _8098 = _8097 < _7020;
    assign _8099 = ~ _8098;
    assign _8087 = _7600[9:9];
    assign _8084 = _8079 - _7020;
    assign _8085 = _8081 ? _8084 : _8079;
    assign _8086 = _8085[62:0];
    assign _8088 = { _8086,
                     _8087 };
    assign _8089 = _8088 < _7020;
    assign _8090 = ~ _8089;
    assign _8078 = _7600[10:10];
    assign _8075 = _8070 - _7020;
    assign _8076 = _8072 ? _8075 : _8070;
    assign _8077 = _8076[62:0];
    assign _8079 = { _8077,
                     _8078 };
    assign _8080 = _8079 < _7020;
    assign _8081 = ~ _8080;
    assign _8069 = _7600[11:11];
    assign _8066 = _8061 - _7020;
    assign _8067 = _8063 ? _8066 : _8061;
    assign _8068 = _8067[62:0];
    assign _8070 = { _8068,
                     _8069 };
    assign _8071 = _8070 < _7020;
    assign _8072 = ~ _8071;
    assign _8060 = _7600[12:12];
    assign _8057 = _8052 - _7020;
    assign _8058 = _8054 ? _8057 : _8052;
    assign _8059 = _8058[62:0];
    assign _8061 = { _8059,
                     _8060 };
    assign _8062 = _8061 < _7020;
    assign _8063 = ~ _8062;
    assign _8051 = _7600[13:13];
    assign _8048 = _8043 - _7020;
    assign _8049 = _8045 ? _8048 : _8043;
    assign _8050 = _8049[62:0];
    assign _8052 = { _8050,
                     _8051 };
    assign _8053 = _8052 < _7020;
    assign _8054 = ~ _8053;
    assign _8042 = _7600[14:14];
    assign _8039 = _8034 - _7020;
    assign _8040 = _8036 ? _8039 : _8034;
    assign _8041 = _8040[62:0];
    assign _8043 = { _8041,
                     _8042 };
    assign _8044 = _8043 < _7020;
    assign _8045 = ~ _8044;
    assign _8033 = _7600[15:15];
    assign _8030 = _8025 - _7020;
    assign _8031 = _8027 ? _8030 : _8025;
    assign _8032 = _8031[62:0];
    assign _8034 = { _8032,
                     _8033 };
    assign _8035 = _8034 < _7020;
    assign _8036 = ~ _8035;
    assign _8024 = _7600[16:16];
    assign _8021 = _8016 - _7020;
    assign _8022 = _8018 ? _8021 : _8016;
    assign _8023 = _8022[62:0];
    assign _8025 = { _8023,
                     _8024 };
    assign _8026 = _8025 < _7020;
    assign _8027 = ~ _8026;
    assign _8015 = _7600[17:17];
    assign _8012 = _8007 - _7020;
    assign _8013 = _8009 ? _8012 : _8007;
    assign _8014 = _8013[62:0];
    assign _8016 = { _8014,
                     _8015 };
    assign _8017 = _8016 < _7020;
    assign _8018 = ~ _8017;
    assign _8006 = _7600[18:18];
    assign _8003 = _7998 - _7020;
    assign _8004 = _8000 ? _8003 : _7998;
    assign _8005 = _8004[62:0];
    assign _8007 = { _8005,
                     _8006 };
    assign _8008 = _8007 < _7020;
    assign _8009 = ~ _8008;
    assign _7997 = _7600[19:19];
    assign _7994 = _7989 - _7020;
    assign _7995 = _7991 ? _7994 : _7989;
    assign _7996 = _7995[62:0];
    assign _7998 = { _7996,
                     _7997 };
    assign _7999 = _7998 < _7020;
    assign _8000 = ~ _7999;
    assign _7988 = _7600[20:20];
    assign _7985 = _7980 - _7020;
    assign _7986 = _7982 ? _7985 : _7980;
    assign _7987 = _7986[62:0];
    assign _7989 = { _7987,
                     _7988 };
    assign _7990 = _7989 < _7020;
    assign _7991 = ~ _7990;
    assign _7979 = _7600[21:21];
    assign _7976 = _7971 - _7020;
    assign _7977 = _7973 ? _7976 : _7971;
    assign _7978 = _7977[62:0];
    assign _7980 = { _7978,
                     _7979 };
    assign _7981 = _7980 < _7020;
    assign _7982 = ~ _7981;
    assign _7970 = _7600[22:22];
    assign _7967 = _7962 - _7020;
    assign _7968 = _7964 ? _7967 : _7962;
    assign _7969 = _7968[62:0];
    assign _7971 = { _7969,
                     _7970 };
    assign _7972 = _7971 < _7020;
    assign _7973 = ~ _7972;
    assign _7961 = _7600[23:23];
    assign _7958 = _7953 - _7020;
    assign _7959 = _7955 ? _7958 : _7953;
    assign _7960 = _7959[62:0];
    assign _7962 = { _7960,
                     _7961 };
    assign _7963 = _7962 < _7020;
    assign _7964 = ~ _7963;
    assign _7952 = _7600[24:24];
    assign _7949 = _7944 - _7020;
    assign _7950 = _7946 ? _7949 : _7944;
    assign _7951 = _7950[62:0];
    assign _7953 = { _7951,
                     _7952 };
    assign _7954 = _7953 < _7020;
    assign _7955 = ~ _7954;
    assign _7943 = _7600[25:25];
    assign _7940 = _7935 - _7020;
    assign _7941 = _7937 ? _7940 : _7935;
    assign _7942 = _7941[62:0];
    assign _7944 = { _7942,
                     _7943 };
    assign _7945 = _7944 < _7020;
    assign _7946 = ~ _7945;
    assign _7934 = _7600[26:26];
    assign _7931 = _7926 - _7020;
    assign _7932 = _7928 ? _7931 : _7926;
    assign _7933 = _7932[62:0];
    assign _7935 = { _7933,
                     _7934 };
    assign _7936 = _7935 < _7020;
    assign _7937 = ~ _7936;
    assign _7925 = _7600[27:27];
    assign _7922 = _7917 - _7020;
    assign _7923 = _7919 ? _7922 : _7917;
    assign _7924 = _7923[62:0];
    assign _7926 = { _7924,
                     _7925 };
    assign _7927 = _7926 < _7020;
    assign _7928 = ~ _7927;
    assign _7916 = _7600[28:28];
    assign _7913 = _7908 - _7020;
    assign _7914 = _7910 ? _7913 : _7908;
    assign _7915 = _7914[62:0];
    assign _7917 = { _7915,
                     _7916 };
    assign _7918 = _7917 < _7020;
    assign _7919 = ~ _7918;
    assign _7907 = _7600[29:29];
    assign _7904 = _7899 - _7020;
    assign _7905 = _7901 ? _7904 : _7899;
    assign _7906 = _7905[62:0];
    assign _7908 = { _7906,
                     _7907 };
    assign _7909 = _7908 < _7020;
    assign _7910 = ~ _7909;
    assign _7898 = _7600[30:30];
    assign _7895 = _7890 - _7020;
    assign _7896 = _7892 ? _7895 : _7890;
    assign _7897 = _7896[62:0];
    assign _7899 = { _7897,
                     _7898 };
    assign _7900 = _7899 < _7020;
    assign _7901 = ~ _7900;
    assign _7889 = _7600[31:31];
    assign _7886 = _7881 - _7020;
    assign _7887 = _7883 ? _7886 : _7881;
    assign _7888 = _7887[62:0];
    assign _7890 = { _7888,
                     _7889 };
    assign _7891 = _7890 < _7020;
    assign _7892 = ~ _7891;
    assign _7880 = _7600[32:32];
    assign _7877 = _7872 - _7020;
    assign _7878 = _7874 ? _7877 : _7872;
    assign _7879 = _7878[62:0];
    assign _7881 = { _7879,
                     _7880 };
    assign _7882 = _7881 < _7020;
    assign _7883 = ~ _7882;
    assign _7871 = _7600[33:33];
    assign _7868 = _7863 - _7020;
    assign _7869 = _7865 ? _7868 : _7863;
    assign _7870 = _7869[62:0];
    assign _7872 = { _7870,
                     _7871 };
    assign _7873 = _7872 < _7020;
    assign _7874 = ~ _7873;
    assign _7862 = _7600[34:34];
    assign _7859 = _7854 - _7020;
    assign _7860 = _7856 ? _7859 : _7854;
    assign _7861 = _7860[62:0];
    assign _7863 = { _7861,
                     _7862 };
    assign _7864 = _7863 < _7020;
    assign _7865 = ~ _7864;
    assign _7853 = _7600[35:35];
    assign _7850 = _7845 - _7020;
    assign _7851 = _7847 ? _7850 : _7845;
    assign _7852 = _7851[62:0];
    assign _7854 = { _7852,
                     _7853 };
    assign _7855 = _7854 < _7020;
    assign _7856 = ~ _7855;
    assign _7844 = _7600[36:36];
    assign _7841 = _7836 - _7020;
    assign _7842 = _7838 ? _7841 : _7836;
    assign _7843 = _7842[62:0];
    assign _7845 = { _7843,
                     _7844 };
    assign _7846 = _7845 < _7020;
    assign _7847 = ~ _7846;
    assign _7835 = _7600[37:37];
    assign _7832 = _7827 - _7020;
    assign _7833 = _7829 ? _7832 : _7827;
    assign _7834 = _7833[62:0];
    assign _7836 = { _7834,
                     _7835 };
    assign _7837 = _7836 < _7020;
    assign _7838 = ~ _7837;
    assign _7826 = _7600[38:38];
    assign _7823 = _7818 - _7020;
    assign _7824 = _7820 ? _7823 : _7818;
    assign _7825 = _7824[62:0];
    assign _7827 = { _7825,
                     _7826 };
    assign _7828 = _7827 < _7020;
    assign _7829 = ~ _7828;
    assign _7817 = _7600[39:39];
    assign _7814 = _7809 - _7020;
    assign _7815 = _7811 ? _7814 : _7809;
    assign _7816 = _7815[62:0];
    assign _7818 = { _7816,
                     _7817 };
    assign _7819 = _7818 < _7020;
    assign _7820 = ~ _7819;
    assign _7808 = _7600[40:40];
    assign _7805 = _7800 - _7020;
    assign _7806 = _7802 ? _7805 : _7800;
    assign _7807 = _7806[62:0];
    assign _7809 = { _7807,
                     _7808 };
    assign _7810 = _7809 < _7020;
    assign _7811 = ~ _7810;
    assign _7799 = _7600[41:41];
    assign _7796 = _7791 - _7020;
    assign _7797 = _7793 ? _7796 : _7791;
    assign _7798 = _7797[62:0];
    assign _7800 = { _7798,
                     _7799 };
    assign _7801 = _7800 < _7020;
    assign _7802 = ~ _7801;
    assign _7790 = _7600[42:42];
    assign _7787 = _7782 - _7020;
    assign _7788 = _7784 ? _7787 : _7782;
    assign _7789 = _7788[62:0];
    assign _7791 = { _7789,
                     _7790 };
    assign _7792 = _7791 < _7020;
    assign _7793 = ~ _7792;
    assign _7781 = _7600[43:43];
    assign _7778 = _7773 - _7020;
    assign _7779 = _7775 ? _7778 : _7773;
    assign _7780 = _7779[62:0];
    assign _7782 = { _7780,
                     _7781 };
    assign _7783 = _7782 < _7020;
    assign _7784 = ~ _7783;
    assign _7772 = _7600[44:44];
    assign _7769 = _7764 - _7020;
    assign _7770 = _7766 ? _7769 : _7764;
    assign _7771 = _7770[62:0];
    assign _7773 = { _7771,
                     _7772 };
    assign _7774 = _7773 < _7020;
    assign _7775 = ~ _7774;
    assign _7763 = _7600[45:45];
    assign _7760 = _7755 - _7020;
    assign _7761 = _7757 ? _7760 : _7755;
    assign _7762 = _7761[62:0];
    assign _7764 = { _7762,
                     _7763 };
    assign _7765 = _7764 < _7020;
    assign _7766 = ~ _7765;
    assign _7754 = _7600[46:46];
    assign _7751 = _7746 - _7020;
    assign _7752 = _7748 ? _7751 : _7746;
    assign _7753 = _7752[62:0];
    assign _7755 = { _7753,
                     _7754 };
    assign _7756 = _7755 < _7020;
    assign _7757 = ~ _7756;
    assign _7745 = _7600[47:47];
    assign _7742 = _7737 - _7020;
    assign _7743 = _7739 ? _7742 : _7737;
    assign _7744 = _7743[62:0];
    assign _7746 = { _7744,
                     _7745 };
    assign _7747 = _7746 < _7020;
    assign _7748 = ~ _7747;
    assign _7736 = _7600[48:48];
    assign _7733 = _7728 - _7020;
    assign _7734 = _7730 ? _7733 : _7728;
    assign _7735 = _7734[62:0];
    assign _7737 = { _7735,
                     _7736 };
    assign _7738 = _7737 < _7020;
    assign _7739 = ~ _7738;
    assign _7727 = _7600[49:49];
    assign _7724 = _7719 - _7020;
    assign _7725 = _7721 ? _7724 : _7719;
    assign _7726 = _7725[62:0];
    assign _7728 = { _7726,
                     _7727 };
    assign _7729 = _7728 < _7020;
    assign _7730 = ~ _7729;
    assign _7718 = _7600[50:50];
    assign _7715 = _7710 - _7020;
    assign _7716 = _7712 ? _7715 : _7710;
    assign _7717 = _7716[62:0];
    assign _7719 = { _7717,
                     _7718 };
    assign _7720 = _7719 < _7020;
    assign _7721 = ~ _7720;
    assign _7709 = _7600[51:51];
    assign _7706 = _7701 - _7020;
    assign _7707 = _7703 ? _7706 : _7701;
    assign _7708 = _7707[62:0];
    assign _7710 = { _7708,
                     _7709 };
    assign _7711 = _7710 < _7020;
    assign _7712 = ~ _7711;
    assign _7700 = _7600[52:52];
    assign _7697 = _7692 - _7020;
    assign _7698 = _7694 ? _7697 : _7692;
    assign _7699 = _7698[62:0];
    assign _7701 = { _7699,
                     _7700 };
    assign _7702 = _7701 < _7020;
    assign _7703 = ~ _7702;
    assign _7691 = _7600[53:53];
    assign _7688 = _7683 - _7020;
    assign _7689 = _7685 ? _7688 : _7683;
    assign _7690 = _7689[62:0];
    assign _7692 = { _7690,
                     _7691 };
    assign _7693 = _7692 < _7020;
    assign _7694 = ~ _7693;
    assign _7682 = _7600[54:54];
    assign _7679 = _7674 - _7020;
    assign _7680 = _7676 ? _7679 : _7674;
    assign _7681 = _7680[62:0];
    assign _7683 = { _7681,
                     _7682 };
    assign _7684 = _7683 < _7020;
    assign _7685 = ~ _7684;
    assign _7673 = _7600[55:55];
    assign _7670 = _7665 - _7020;
    assign _7671 = _7667 ? _7670 : _7665;
    assign _7672 = _7671[62:0];
    assign _7674 = { _7672,
                     _7673 };
    assign _7675 = _7674 < _7020;
    assign _7676 = ~ _7675;
    assign _7664 = _7600[56:56];
    assign _7661 = _7656 - _7020;
    assign _7662 = _7658 ? _7661 : _7656;
    assign _7663 = _7662[62:0];
    assign _7665 = { _7663,
                     _7664 };
    assign _7666 = _7665 < _7020;
    assign _7667 = ~ _7666;
    assign _7655 = _7600[57:57];
    assign _7652 = _7647 - _7020;
    assign _7653 = _7649 ? _7652 : _7647;
    assign _7654 = _7653[62:0];
    assign _7656 = { _7654,
                     _7655 };
    assign _7657 = _7656 < _7020;
    assign _7658 = ~ _7657;
    assign _7646 = _7600[58:58];
    assign _7643 = _7638 - _7020;
    assign _7644 = _7640 ? _7643 : _7638;
    assign _7645 = _7644[62:0];
    assign _7647 = { _7645,
                     _7646 };
    assign _7648 = _7647 < _7020;
    assign _7649 = ~ _7648;
    assign _7637 = _7600[59:59];
    assign _7634 = _7629 - _7020;
    assign _7635 = _7631 ? _7634 : _7629;
    assign _7636 = _7635[62:0];
    assign _7638 = { _7636,
                     _7637 };
    assign _7639 = _7638 < _7020;
    assign _7640 = ~ _7639;
    assign _7628 = _7600[60:60];
    assign _7625 = _7620 - _7020;
    assign _7626 = _7622 ? _7625 : _7620;
    assign _7627 = _7626[62:0];
    assign _7629 = { _7627,
                     _7628 };
    assign _7630 = _7629 < _7020;
    assign _7631 = ~ _7630;
    assign _7619 = _7600[61:61];
    assign _7616 = _7611 - _7020;
    assign _7617 = _7613 ? _7616 : _7611;
    assign _7618 = _7617[62:0];
    assign _7620 = { _7618,
                     _7619 };
    assign _7621 = _7620 < _7020;
    assign _7622 = ~ _7621;
    assign _7610 = _7600[62:62];
    assign _7607 = _7602 - _7020;
    assign _7608 = _7604 ? _7607 : _7602;
    assign _7609 = _7608[62:0];
    assign _7611 = { _7609,
                     _7610 };
    assign _7612 = _7611 < _7020;
    assign _7613 = ~ _7612;
    assign _7600 = _7012 - _7594;
    assign _7601 = _7600[63:63];
    assign _7602 = { _22185,
                     _7601 };
    assign _7603 = _7602 < _7020;
    assign _7604 = ~ _7603;
    assign _7605 = { _22185,
                     _7604 };
    assign _7606 = _7605[62:0];
    assign _7614 = { _7606,
                     _7613 };
    assign _7615 = _7614[62:0];
    assign _7623 = { _7615,
                     _7622 };
    assign _7624 = _7623[62:0];
    assign _7632 = { _7624,
                     _7631 };
    assign _7633 = _7632[62:0];
    assign _7641 = { _7633,
                     _7640 };
    assign _7642 = _7641[62:0];
    assign _7650 = { _7642,
                     _7649 };
    assign _7651 = _7650[62:0];
    assign _7659 = { _7651,
                     _7658 };
    assign _7660 = _7659[62:0];
    assign _7668 = { _7660,
                     _7667 };
    assign _7669 = _7668[62:0];
    assign _7677 = { _7669,
                     _7676 };
    assign _7678 = _7677[62:0];
    assign _7686 = { _7678,
                     _7685 };
    assign _7687 = _7686[62:0];
    assign _7695 = { _7687,
                     _7694 };
    assign _7696 = _7695[62:0];
    assign _7704 = { _7696,
                     _7703 };
    assign _7705 = _7704[62:0];
    assign _7713 = { _7705,
                     _7712 };
    assign _7714 = _7713[62:0];
    assign _7722 = { _7714,
                     _7721 };
    assign _7723 = _7722[62:0];
    assign _7731 = { _7723,
                     _7730 };
    assign _7732 = _7731[62:0];
    assign _7740 = { _7732,
                     _7739 };
    assign _7741 = _7740[62:0];
    assign _7749 = { _7741,
                     _7748 };
    assign _7750 = _7749[62:0];
    assign _7758 = { _7750,
                     _7757 };
    assign _7759 = _7758[62:0];
    assign _7767 = { _7759,
                     _7766 };
    assign _7768 = _7767[62:0];
    assign _7776 = { _7768,
                     _7775 };
    assign _7777 = _7776[62:0];
    assign _7785 = { _7777,
                     _7784 };
    assign _7786 = _7785[62:0];
    assign _7794 = { _7786,
                     _7793 };
    assign _7795 = _7794[62:0];
    assign _7803 = { _7795,
                     _7802 };
    assign _7804 = _7803[62:0];
    assign _7812 = { _7804,
                     _7811 };
    assign _7813 = _7812[62:0];
    assign _7821 = { _7813,
                     _7820 };
    assign _7822 = _7821[62:0];
    assign _7830 = { _7822,
                     _7829 };
    assign _7831 = _7830[62:0];
    assign _7839 = { _7831,
                     _7838 };
    assign _7840 = _7839[62:0];
    assign _7848 = { _7840,
                     _7847 };
    assign _7849 = _7848[62:0];
    assign _7857 = { _7849,
                     _7856 };
    assign _7858 = _7857[62:0];
    assign _7866 = { _7858,
                     _7865 };
    assign _7867 = _7866[62:0];
    assign _7875 = { _7867,
                     _7874 };
    assign _7876 = _7875[62:0];
    assign _7884 = { _7876,
                     _7883 };
    assign _7885 = _7884[62:0];
    assign _7893 = { _7885,
                     _7892 };
    assign _7894 = _7893[62:0];
    assign _7902 = { _7894,
                     _7901 };
    assign _7903 = _7902[62:0];
    assign _7911 = { _7903,
                     _7910 };
    assign _7912 = _7911[62:0];
    assign _7920 = { _7912,
                     _7919 };
    assign _7921 = _7920[62:0];
    assign _7929 = { _7921,
                     _7928 };
    assign _7930 = _7929[62:0];
    assign _7938 = { _7930,
                     _7937 };
    assign _7939 = _7938[62:0];
    assign _7947 = { _7939,
                     _7946 };
    assign _7948 = _7947[62:0];
    assign _7956 = { _7948,
                     _7955 };
    assign _7957 = _7956[62:0];
    assign _7965 = { _7957,
                     _7964 };
    assign _7966 = _7965[62:0];
    assign _7974 = { _7966,
                     _7973 };
    assign _7975 = _7974[62:0];
    assign _7983 = { _7975,
                     _7982 };
    assign _7984 = _7983[62:0];
    assign _7992 = { _7984,
                     _7991 };
    assign _7993 = _7992[62:0];
    assign _8001 = { _7993,
                     _8000 };
    assign _8002 = _8001[62:0];
    assign _8010 = { _8002,
                     _8009 };
    assign _8011 = _8010[62:0];
    assign _8019 = { _8011,
                     _8018 };
    assign _8020 = _8019[62:0];
    assign _8028 = { _8020,
                     _8027 };
    assign _8029 = _8028[62:0];
    assign _8037 = { _8029,
                     _8036 };
    assign _8038 = _8037[62:0];
    assign _8046 = { _8038,
                     _8045 };
    assign _8047 = _8046[62:0];
    assign _8055 = { _8047,
                     _8054 };
    assign _8056 = _8055[62:0];
    assign _8064 = { _8056,
                     _8063 };
    assign _8065 = _8064[62:0];
    assign _8073 = { _8065,
                     _8072 };
    assign _8074 = _8073[62:0];
    assign _8082 = { _8074,
                     _8081 };
    assign _8083 = _8082[62:0];
    assign _8091 = { _8083,
                     _8090 };
    assign _8092 = _8091[62:0];
    assign _8100 = { _8092,
                     _8099 };
    assign _8101 = _8100[62:0];
    assign _8109 = { _8101,
                     _8108 };
    assign _8110 = _8109[62:0];
    assign _8118 = { _8110,
                     _8117 };
    assign _8119 = _8118[62:0];
    assign _8127 = { _8119,
                     _8126 };
    assign _8128 = _8127[62:0];
    assign _8136 = { _8128,
                     _8135 };
    assign _8137 = _8136[62:0];
    assign _8145 = { _8137,
                     _8144 };
    assign _8146 = _8145[62:0];
    assign _8154 = { _8146,
                     _8153 };
    assign _8155 = _8154[62:0];
    assign _8163 = { _8155,
                     _8162 };
    assign _8164 = _8163[62:0];
    assign _8172 = { _8164,
                     _8171 };
    assign _8174 = _8172 + _22186;
    assign _8175 = _8174 * _7594;
    assign _8176 = _8175[63:0];
    assign _8758 = _8176 + _8757;
    assign _7586 = _7017[0:0];
    assign _7583 = _7578 - _7020;
    assign _7584 = _7580 ? _7583 : _7578;
    assign _7585 = _7584[62:0];
    assign _7587 = { _7585,
                     _7586 };
    assign _7588 = _7587 < _7020;
    assign _7589 = ~ _7588;
    assign _7577 = _7017[1:1];
    assign _7574 = _7569 - _7020;
    assign _7575 = _7571 ? _7574 : _7569;
    assign _7576 = _7575[62:0];
    assign _7578 = { _7576,
                     _7577 };
    assign _7579 = _7578 < _7020;
    assign _7580 = ~ _7579;
    assign _7568 = _7017[2:2];
    assign _7565 = _7560 - _7020;
    assign _7566 = _7562 ? _7565 : _7560;
    assign _7567 = _7566[62:0];
    assign _7569 = { _7567,
                     _7568 };
    assign _7570 = _7569 < _7020;
    assign _7571 = ~ _7570;
    assign _7559 = _7017[3:3];
    assign _7556 = _7551 - _7020;
    assign _7557 = _7553 ? _7556 : _7551;
    assign _7558 = _7557[62:0];
    assign _7560 = { _7558,
                     _7559 };
    assign _7561 = _7560 < _7020;
    assign _7562 = ~ _7561;
    assign _7550 = _7017[4:4];
    assign _7547 = _7542 - _7020;
    assign _7548 = _7544 ? _7547 : _7542;
    assign _7549 = _7548[62:0];
    assign _7551 = { _7549,
                     _7550 };
    assign _7552 = _7551 < _7020;
    assign _7553 = ~ _7552;
    assign _7541 = _7017[5:5];
    assign _7538 = _7533 - _7020;
    assign _7539 = _7535 ? _7538 : _7533;
    assign _7540 = _7539[62:0];
    assign _7542 = { _7540,
                     _7541 };
    assign _7543 = _7542 < _7020;
    assign _7544 = ~ _7543;
    assign _7532 = _7017[6:6];
    assign _7529 = _7524 - _7020;
    assign _7530 = _7526 ? _7529 : _7524;
    assign _7531 = _7530[62:0];
    assign _7533 = { _7531,
                     _7532 };
    assign _7534 = _7533 < _7020;
    assign _7535 = ~ _7534;
    assign _7523 = _7017[7:7];
    assign _7520 = _7515 - _7020;
    assign _7521 = _7517 ? _7520 : _7515;
    assign _7522 = _7521[62:0];
    assign _7524 = { _7522,
                     _7523 };
    assign _7525 = _7524 < _7020;
    assign _7526 = ~ _7525;
    assign _7514 = _7017[8:8];
    assign _7511 = _7506 - _7020;
    assign _7512 = _7508 ? _7511 : _7506;
    assign _7513 = _7512[62:0];
    assign _7515 = { _7513,
                     _7514 };
    assign _7516 = _7515 < _7020;
    assign _7517 = ~ _7516;
    assign _7505 = _7017[9:9];
    assign _7502 = _7497 - _7020;
    assign _7503 = _7499 ? _7502 : _7497;
    assign _7504 = _7503[62:0];
    assign _7506 = { _7504,
                     _7505 };
    assign _7507 = _7506 < _7020;
    assign _7508 = ~ _7507;
    assign _7496 = _7017[10:10];
    assign _7493 = _7488 - _7020;
    assign _7494 = _7490 ? _7493 : _7488;
    assign _7495 = _7494[62:0];
    assign _7497 = { _7495,
                     _7496 };
    assign _7498 = _7497 < _7020;
    assign _7499 = ~ _7498;
    assign _7487 = _7017[11:11];
    assign _7484 = _7479 - _7020;
    assign _7485 = _7481 ? _7484 : _7479;
    assign _7486 = _7485[62:0];
    assign _7488 = { _7486,
                     _7487 };
    assign _7489 = _7488 < _7020;
    assign _7490 = ~ _7489;
    assign _7478 = _7017[12:12];
    assign _7475 = _7470 - _7020;
    assign _7476 = _7472 ? _7475 : _7470;
    assign _7477 = _7476[62:0];
    assign _7479 = { _7477,
                     _7478 };
    assign _7480 = _7479 < _7020;
    assign _7481 = ~ _7480;
    assign _7469 = _7017[13:13];
    assign _7466 = _7461 - _7020;
    assign _7467 = _7463 ? _7466 : _7461;
    assign _7468 = _7467[62:0];
    assign _7470 = { _7468,
                     _7469 };
    assign _7471 = _7470 < _7020;
    assign _7472 = ~ _7471;
    assign _7460 = _7017[14:14];
    assign _7457 = _7452 - _7020;
    assign _7458 = _7454 ? _7457 : _7452;
    assign _7459 = _7458[62:0];
    assign _7461 = { _7459,
                     _7460 };
    assign _7462 = _7461 < _7020;
    assign _7463 = ~ _7462;
    assign _7451 = _7017[15:15];
    assign _7448 = _7443 - _7020;
    assign _7449 = _7445 ? _7448 : _7443;
    assign _7450 = _7449[62:0];
    assign _7452 = { _7450,
                     _7451 };
    assign _7453 = _7452 < _7020;
    assign _7454 = ~ _7453;
    assign _7442 = _7017[16:16];
    assign _7439 = _7434 - _7020;
    assign _7440 = _7436 ? _7439 : _7434;
    assign _7441 = _7440[62:0];
    assign _7443 = { _7441,
                     _7442 };
    assign _7444 = _7443 < _7020;
    assign _7445 = ~ _7444;
    assign _7433 = _7017[17:17];
    assign _7430 = _7425 - _7020;
    assign _7431 = _7427 ? _7430 : _7425;
    assign _7432 = _7431[62:0];
    assign _7434 = { _7432,
                     _7433 };
    assign _7435 = _7434 < _7020;
    assign _7436 = ~ _7435;
    assign _7424 = _7017[18:18];
    assign _7421 = _7416 - _7020;
    assign _7422 = _7418 ? _7421 : _7416;
    assign _7423 = _7422[62:0];
    assign _7425 = { _7423,
                     _7424 };
    assign _7426 = _7425 < _7020;
    assign _7427 = ~ _7426;
    assign _7415 = _7017[19:19];
    assign _7412 = _7407 - _7020;
    assign _7413 = _7409 ? _7412 : _7407;
    assign _7414 = _7413[62:0];
    assign _7416 = { _7414,
                     _7415 };
    assign _7417 = _7416 < _7020;
    assign _7418 = ~ _7417;
    assign _7406 = _7017[20:20];
    assign _7403 = _7398 - _7020;
    assign _7404 = _7400 ? _7403 : _7398;
    assign _7405 = _7404[62:0];
    assign _7407 = { _7405,
                     _7406 };
    assign _7408 = _7407 < _7020;
    assign _7409 = ~ _7408;
    assign _7397 = _7017[21:21];
    assign _7394 = _7389 - _7020;
    assign _7395 = _7391 ? _7394 : _7389;
    assign _7396 = _7395[62:0];
    assign _7398 = { _7396,
                     _7397 };
    assign _7399 = _7398 < _7020;
    assign _7400 = ~ _7399;
    assign _7388 = _7017[22:22];
    assign _7385 = _7380 - _7020;
    assign _7386 = _7382 ? _7385 : _7380;
    assign _7387 = _7386[62:0];
    assign _7389 = { _7387,
                     _7388 };
    assign _7390 = _7389 < _7020;
    assign _7391 = ~ _7390;
    assign _7379 = _7017[23:23];
    assign _7376 = _7371 - _7020;
    assign _7377 = _7373 ? _7376 : _7371;
    assign _7378 = _7377[62:0];
    assign _7380 = { _7378,
                     _7379 };
    assign _7381 = _7380 < _7020;
    assign _7382 = ~ _7381;
    assign _7370 = _7017[24:24];
    assign _7367 = _7362 - _7020;
    assign _7368 = _7364 ? _7367 : _7362;
    assign _7369 = _7368[62:0];
    assign _7371 = { _7369,
                     _7370 };
    assign _7372 = _7371 < _7020;
    assign _7373 = ~ _7372;
    assign _7361 = _7017[25:25];
    assign _7358 = _7353 - _7020;
    assign _7359 = _7355 ? _7358 : _7353;
    assign _7360 = _7359[62:0];
    assign _7362 = { _7360,
                     _7361 };
    assign _7363 = _7362 < _7020;
    assign _7364 = ~ _7363;
    assign _7352 = _7017[26:26];
    assign _7349 = _7344 - _7020;
    assign _7350 = _7346 ? _7349 : _7344;
    assign _7351 = _7350[62:0];
    assign _7353 = { _7351,
                     _7352 };
    assign _7354 = _7353 < _7020;
    assign _7355 = ~ _7354;
    assign _7343 = _7017[27:27];
    assign _7340 = _7335 - _7020;
    assign _7341 = _7337 ? _7340 : _7335;
    assign _7342 = _7341[62:0];
    assign _7344 = { _7342,
                     _7343 };
    assign _7345 = _7344 < _7020;
    assign _7346 = ~ _7345;
    assign _7334 = _7017[28:28];
    assign _7331 = _7326 - _7020;
    assign _7332 = _7328 ? _7331 : _7326;
    assign _7333 = _7332[62:0];
    assign _7335 = { _7333,
                     _7334 };
    assign _7336 = _7335 < _7020;
    assign _7337 = ~ _7336;
    assign _7325 = _7017[29:29];
    assign _7322 = _7317 - _7020;
    assign _7323 = _7319 ? _7322 : _7317;
    assign _7324 = _7323[62:0];
    assign _7326 = { _7324,
                     _7325 };
    assign _7327 = _7326 < _7020;
    assign _7328 = ~ _7327;
    assign _7316 = _7017[30:30];
    assign _7313 = _7308 - _7020;
    assign _7314 = _7310 ? _7313 : _7308;
    assign _7315 = _7314[62:0];
    assign _7317 = { _7315,
                     _7316 };
    assign _7318 = _7317 < _7020;
    assign _7319 = ~ _7318;
    assign _7307 = _7017[31:31];
    assign _7304 = _7299 - _7020;
    assign _7305 = _7301 ? _7304 : _7299;
    assign _7306 = _7305[62:0];
    assign _7308 = { _7306,
                     _7307 };
    assign _7309 = _7308 < _7020;
    assign _7310 = ~ _7309;
    assign _7298 = _7017[32:32];
    assign _7295 = _7290 - _7020;
    assign _7296 = _7292 ? _7295 : _7290;
    assign _7297 = _7296[62:0];
    assign _7299 = { _7297,
                     _7298 };
    assign _7300 = _7299 < _7020;
    assign _7301 = ~ _7300;
    assign _7289 = _7017[33:33];
    assign _7286 = _7281 - _7020;
    assign _7287 = _7283 ? _7286 : _7281;
    assign _7288 = _7287[62:0];
    assign _7290 = { _7288,
                     _7289 };
    assign _7291 = _7290 < _7020;
    assign _7292 = ~ _7291;
    assign _7280 = _7017[34:34];
    assign _7277 = _7272 - _7020;
    assign _7278 = _7274 ? _7277 : _7272;
    assign _7279 = _7278[62:0];
    assign _7281 = { _7279,
                     _7280 };
    assign _7282 = _7281 < _7020;
    assign _7283 = ~ _7282;
    assign _7271 = _7017[35:35];
    assign _7268 = _7263 - _7020;
    assign _7269 = _7265 ? _7268 : _7263;
    assign _7270 = _7269[62:0];
    assign _7272 = { _7270,
                     _7271 };
    assign _7273 = _7272 < _7020;
    assign _7274 = ~ _7273;
    assign _7262 = _7017[36:36];
    assign _7259 = _7254 - _7020;
    assign _7260 = _7256 ? _7259 : _7254;
    assign _7261 = _7260[62:0];
    assign _7263 = { _7261,
                     _7262 };
    assign _7264 = _7263 < _7020;
    assign _7265 = ~ _7264;
    assign _7253 = _7017[37:37];
    assign _7250 = _7245 - _7020;
    assign _7251 = _7247 ? _7250 : _7245;
    assign _7252 = _7251[62:0];
    assign _7254 = { _7252,
                     _7253 };
    assign _7255 = _7254 < _7020;
    assign _7256 = ~ _7255;
    assign _7244 = _7017[38:38];
    assign _7241 = _7236 - _7020;
    assign _7242 = _7238 ? _7241 : _7236;
    assign _7243 = _7242[62:0];
    assign _7245 = { _7243,
                     _7244 };
    assign _7246 = _7245 < _7020;
    assign _7247 = ~ _7246;
    assign _7235 = _7017[39:39];
    assign _7232 = _7227 - _7020;
    assign _7233 = _7229 ? _7232 : _7227;
    assign _7234 = _7233[62:0];
    assign _7236 = { _7234,
                     _7235 };
    assign _7237 = _7236 < _7020;
    assign _7238 = ~ _7237;
    assign _7226 = _7017[40:40];
    assign _7223 = _7218 - _7020;
    assign _7224 = _7220 ? _7223 : _7218;
    assign _7225 = _7224[62:0];
    assign _7227 = { _7225,
                     _7226 };
    assign _7228 = _7227 < _7020;
    assign _7229 = ~ _7228;
    assign _7217 = _7017[41:41];
    assign _7214 = _7209 - _7020;
    assign _7215 = _7211 ? _7214 : _7209;
    assign _7216 = _7215[62:0];
    assign _7218 = { _7216,
                     _7217 };
    assign _7219 = _7218 < _7020;
    assign _7220 = ~ _7219;
    assign _7208 = _7017[42:42];
    assign _7205 = _7200 - _7020;
    assign _7206 = _7202 ? _7205 : _7200;
    assign _7207 = _7206[62:0];
    assign _7209 = { _7207,
                     _7208 };
    assign _7210 = _7209 < _7020;
    assign _7211 = ~ _7210;
    assign _7199 = _7017[43:43];
    assign _7196 = _7191 - _7020;
    assign _7197 = _7193 ? _7196 : _7191;
    assign _7198 = _7197[62:0];
    assign _7200 = { _7198,
                     _7199 };
    assign _7201 = _7200 < _7020;
    assign _7202 = ~ _7201;
    assign _7190 = _7017[44:44];
    assign _7187 = _7182 - _7020;
    assign _7188 = _7184 ? _7187 : _7182;
    assign _7189 = _7188[62:0];
    assign _7191 = { _7189,
                     _7190 };
    assign _7192 = _7191 < _7020;
    assign _7193 = ~ _7192;
    assign _7181 = _7017[45:45];
    assign _7178 = _7173 - _7020;
    assign _7179 = _7175 ? _7178 : _7173;
    assign _7180 = _7179[62:0];
    assign _7182 = { _7180,
                     _7181 };
    assign _7183 = _7182 < _7020;
    assign _7184 = ~ _7183;
    assign _7172 = _7017[46:46];
    assign _7169 = _7164 - _7020;
    assign _7170 = _7166 ? _7169 : _7164;
    assign _7171 = _7170[62:0];
    assign _7173 = { _7171,
                     _7172 };
    assign _7174 = _7173 < _7020;
    assign _7175 = ~ _7174;
    assign _7163 = _7017[47:47];
    assign _7160 = _7155 - _7020;
    assign _7161 = _7157 ? _7160 : _7155;
    assign _7162 = _7161[62:0];
    assign _7164 = { _7162,
                     _7163 };
    assign _7165 = _7164 < _7020;
    assign _7166 = ~ _7165;
    assign _7154 = _7017[48:48];
    assign _7151 = _7146 - _7020;
    assign _7152 = _7148 ? _7151 : _7146;
    assign _7153 = _7152[62:0];
    assign _7155 = { _7153,
                     _7154 };
    assign _7156 = _7155 < _7020;
    assign _7157 = ~ _7156;
    assign _7145 = _7017[49:49];
    assign _7142 = _7137 - _7020;
    assign _7143 = _7139 ? _7142 : _7137;
    assign _7144 = _7143[62:0];
    assign _7146 = { _7144,
                     _7145 };
    assign _7147 = _7146 < _7020;
    assign _7148 = ~ _7147;
    assign _7136 = _7017[50:50];
    assign _7133 = _7128 - _7020;
    assign _7134 = _7130 ? _7133 : _7128;
    assign _7135 = _7134[62:0];
    assign _7137 = { _7135,
                     _7136 };
    assign _7138 = _7137 < _7020;
    assign _7139 = ~ _7138;
    assign _7127 = _7017[51:51];
    assign _7124 = _7119 - _7020;
    assign _7125 = _7121 ? _7124 : _7119;
    assign _7126 = _7125[62:0];
    assign _7128 = { _7126,
                     _7127 };
    assign _7129 = _7128 < _7020;
    assign _7130 = ~ _7129;
    assign _7118 = _7017[52:52];
    assign _7115 = _7110 - _7020;
    assign _7116 = _7112 ? _7115 : _7110;
    assign _7117 = _7116[62:0];
    assign _7119 = { _7117,
                     _7118 };
    assign _7120 = _7119 < _7020;
    assign _7121 = ~ _7120;
    assign _7109 = _7017[53:53];
    assign _7106 = _7101 - _7020;
    assign _7107 = _7103 ? _7106 : _7101;
    assign _7108 = _7107[62:0];
    assign _7110 = { _7108,
                     _7109 };
    assign _7111 = _7110 < _7020;
    assign _7112 = ~ _7111;
    assign _7100 = _7017[54:54];
    assign _7097 = _7092 - _7020;
    assign _7098 = _7094 ? _7097 : _7092;
    assign _7099 = _7098[62:0];
    assign _7101 = { _7099,
                     _7100 };
    assign _7102 = _7101 < _7020;
    assign _7103 = ~ _7102;
    assign _7091 = _7017[55:55];
    assign _7088 = _7083 - _7020;
    assign _7089 = _7085 ? _7088 : _7083;
    assign _7090 = _7089[62:0];
    assign _7092 = { _7090,
                     _7091 };
    assign _7093 = _7092 < _7020;
    assign _7094 = ~ _7093;
    assign _7082 = _7017[56:56];
    assign _7079 = _7074 - _7020;
    assign _7080 = _7076 ? _7079 : _7074;
    assign _7081 = _7080[62:0];
    assign _7083 = { _7081,
                     _7082 };
    assign _7084 = _7083 < _7020;
    assign _7085 = ~ _7084;
    assign _7073 = _7017[57:57];
    assign _7070 = _7065 - _7020;
    assign _7071 = _7067 ? _7070 : _7065;
    assign _7072 = _7071[62:0];
    assign _7074 = { _7072,
                     _7073 };
    assign _7075 = _7074 < _7020;
    assign _7076 = ~ _7075;
    assign _7064 = _7017[58:58];
    assign _7061 = _7056 - _7020;
    assign _7062 = _7058 ? _7061 : _7056;
    assign _7063 = _7062[62:0];
    assign _7065 = { _7063,
                     _7064 };
    assign _7066 = _7065 < _7020;
    assign _7067 = ~ _7066;
    assign _7055 = _7017[59:59];
    assign _7052 = _7047 - _7020;
    assign _7053 = _7049 ? _7052 : _7047;
    assign _7054 = _7053[62:0];
    assign _7056 = { _7054,
                     _7055 };
    assign _7057 = _7056 < _7020;
    assign _7058 = ~ _7057;
    assign _7046 = _7017[60:60];
    assign _7043 = _7038 - _7020;
    assign _7044 = _7040 ? _7043 : _7038;
    assign _7045 = _7044[62:0];
    assign _7047 = { _7045,
                     _7046 };
    assign _7048 = _7047 < _7020;
    assign _7049 = ~ _7048;
    assign _7037 = _7017[61:61];
    assign _7034 = _7029 - _7020;
    assign _7035 = _7031 ? _7034 : _7029;
    assign _7036 = _7035[62:0];
    assign _7038 = { _7036,
                     _7037 };
    assign _7039 = _7038 < _7020;
    assign _7040 = ~ _7039;
    assign _7028 = _7017[62:62];
    assign _7025 = _7019 - _7020;
    assign _7026 = _7022 ? _7025 : _7019;
    assign _7027 = _7026[62:0];
    assign _7029 = { _7027,
                     _7028 };
    assign _7030 = _7029 < _7020;
    assign _7031 = ~ _7030;
    assign _7020 = 64'b0000000000000000000000000000000000000000000000011000011010100001;
    assign _7016 = 64'b0000000000000000000000000000000000000000000000011000011010100000;
    assign _7017 = _3 + _7016;
    assign _7018 = _7017[63:63];
    assign _7019 = { _22185,
                     _7018 };
    assign _7021 = _7019 < _7020;
    assign _7022 = ~ _7021;
    assign _7023 = { _22185,
                     _7022 };
    assign _7024 = _7023[62:0];
    assign _7032 = { _7024,
                     _7031 };
    assign _7033 = _7032[62:0];
    assign _7041 = { _7033,
                     _7040 };
    assign _7042 = _7041[62:0];
    assign _7050 = { _7042,
                     _7049 };
    assign _7051 = _7050[62:0];
    assign _7059 = { _7051,
                     _7058 };
    assign _7060 = _7059[62:0];
    assign _7068 = { _7060,
                     _7067 };
    assign _7069 = _7068[62:0];
    assign _7077 = { _7069,
                     _7076 };
    assign _7078 = _7077[62:0];
    assign _7086 = { _7078,
                     _7085 };
    assign _7087 = _7086[62:0];
    assign _7095 = { _7087,
                     _7094 };
    assign _7096 = _7095[62:0];
    assign _7104 = { _7096,
                     _7103 };
    assign _7105 = _7104[62:0];
    assign _7113 = { _7105,
                     _7112 };
    assign _7114 = _7113[62:0];
    assign _7122 = { _7114,
                     _7121 };
    assign _7123 = _7122[62:0];
    assign _7131 = { _7123,
                     _7130 };
    assign _7132 = _7131[62:0];
    assign _7140 = { _7132,
                     _7139 };
    assign _7141 = _7140[62:0];
    assign _7149 = { _7141,
                     _7148 };
    assign _7150 = _7149[62:0];
    assign _7158 = { _7150,
                     _7157 };
    assign _7159 = _7158[62:0];
    assign _7167 = { _7159,
                     _7166 };
    assign _7168 = _7167[62:0];
    assign _7176 = { _7168,
                     _7175 };
    assign _7177 = _7176[62:0];
    assign _7185 = { _7177,
                     _7184 };
    assign _7186 = _7185[62:0];
    assign _7194 = { _7186,
                     _7193 };
    assign _7195 = _7194[62:0];
    assign _7203 = { _7195,
                     _7202 };
    assign _7204 = _7203[62:0];
    assign _7212 = { _7204,
                     _7211 };
    assign _7213 = _7212[62:0];
    assign _7221 = { _7213,
                     _7220 };
    assign _7222 = _7221[62:0];
    assign _7230 = { _7222,
                     _7229 };
    assign _7231 = _7230[62:0];
    assign _7239 = { _7231,
                     _7238 };
    assign _7240 = _7239[62:0];
    assign _7248 = { _7240,
                     _7247 };
    assign _7249 = _7248[62:0];
    assign _7257 = { _7249,
                     _7256 };
    assign _7258 = _7257[62:0];
    assign _7266 = { _7258,
                     _7265 };
    assign _7267 = _7266[62:0];
    assign _7275 = { _7267,
                     _7274 };
    assign _7276 = _7275[62:0];
    assign _7284 = { _7276,
                     _7283 };
    assign _7285 = _7284[62:0];
    assign _7293 = { _7285,
                     _7292 };
    assign _7294 = _7293[62:0];
    assign _7302 = { _7294,
                     _7301 };
    assign _7303 = _7302[62:0];
    assign _7311 = { _7303,
                     _7310 };
    assign _7312 = _7311[62:0];
    assign _7320 = { _7312,
                     _7319 };
    assign _7321 = _7320[62:0];
    assign _7329 = { _7321,
                     _7328 };
    assign _7330 = _7329[62:0];
    assign _7338 = { _7330,
                     _7337 };
    assign _7339 = _7338[62:0];
    assign _7347 = { _7339,
                     _7346 };
    assign _7348 = _7347[62:0];
    assign _7356 = { _7348,
                     _7355 };
    assign _7357 = _7356[62:0];
    assign _7365 = { _7357,
                     _7364 };
    assign _7366 = _7365[62:0];
    assign _7374 = { _7366,
                     _7373 };
    assign _7375 = _7374[62:0];
    assign _7383 = { _7375,
                     _7382 };
    assign _7384 = _7383[62:0];
    assign _7392 = { _7384,
                     _7391 };
    assign _7393 = _7392[62:0];
    assign _7401 = { _7393,
                     _7400 };
    assign _7402 = _7401[62:0];
    assign _7410 = { _7402,
                     _7409 };
    assign _7411 = _7410[62:0];
    assign _7419 = { _7411,
                     _7418 };
    assign _7420 = _7419[62:0];
    assign _7428 = { _7420,
                     _7427 };
    assign _7429 = _7428[62:0];
    assign _7437 = { _7429,
                     _7436 };
    assign _7438 = _7437[62:0];
    assign _7446 = { _7438,
                     _7445 };
    assign _7447 = _7446[62:0];
    assign _7455 = { _7447,
                     _7454 };
    assign _7456 = _7455[62:0];
    assign _7464 = { _7456,
                     _7463 };
    assign _7465 = _7464[62:0];
    assign _7473 = { _7465,
                     _7472 };
    assign _7474 = _7473[62:0];
    assign _7482 = { _7474,
                     _7481 };
    assign _7483 = _7482[62:0];
    assign _7491 = { _7483,
                     _7490 };
    assign _7492 = _7491[62:0];
    assign _7500 = { _7492,
                     _7499 };
    assign _7501 = _7500[62:0];
    assign _7509 = { _7501,
                     _7508 };
    assign _7510 = _7509[62:0];
    assign _7518 = { _7510,
                     _7517 };
    assign _7519 = _7518[62:0];
    assign _7527 = { _7519,
                     _7526 };
    assign _7528 = _7527[62:0];
    assign _7536 = { _7528,
                     _7535 };
    assign _7537 = _7536[62:0];
    assign _7545 = { _7537,
                     _7544 };
    assign _7546 = _7545[62:0];
    assign _7554 = { _7546,
                     _7553 };
    assign _7555 = _7554[62:0];
    assign _7563 = { _7555,
                     _7562 };
    assign _7564 = _7563[62:0];
    assign _7572 = { _7564,
                     _7571 };
    assign _7573 = _7572[62:0];
    assign _7581 = { _7573,
                     _7580 };
    assign _7582 = _7581[62:0];
    assign _7590 = { _7582,
                     _7589 };
    assign _7591 = _7590 * _7020;
    assign _7592 = _7591[63:0];
    assign _7013 = 64'b0000000000000000000000000000000000111011100110101111000100010000;
    assign _7593 = _7013 < _7592;
    assign _7594 = _7593 ? _7592 : _7013;
    assign _7011 = _5 < _21017;
    assign _7012 = _7011 ? _5 : _21017;
    assign _7595 = _7012 < _7594;
    assign _7596 = ~ _7595;
    assign _8759 = _7596 ? _8758 : _21604;
    assign _7000 = _6431[0:0];
    assign _6997 = _6992 - _22192;
    assign _6998 = _6994 ? _6997 : _6992;
    assign _6999 = _6998[62:0];
    assign _7001 = { _6999,
                     _7000 };
    assign _7002 = _7001 < _22192;
    assign _7003 = ~ _7002;
    assign _6991 = _6431[1:1];
    assign _6988 = _6983 - _22192;
    assign _6989 = _6985 ? _6988 : _6983;
    assign _6990 = _6989[62:0];
    assign _6992 = { _6990,
                     _6991 };
    assign _6993 = _6992 < _22192;
    assign _6994 = ~ _6993;
    assign _6982 = _6431[2:2];
    assign _6979 = _6974 - _22192;
    assign _6980 = _6976 ? _6979 : _6974;
    assign _6981 = _6980[62:0];
    assign _6983 = { _6981,
                     _6982 };
    assign _6984 = _6983 < _22192;
    assign _6985 = ~ _6984;
    assign _6973 = _6431[3:3];
    assign _6970 = _6965 - _22192;
    assign _6971 = _6967 ? _6970 : _6965;
    assign _6972 = _6971[62:0];
    assign _6974 = { _6972,
                     _6973 };
    assign _6975 = _6974 < _22192;
    assign _6976 = ~ _6975;
    assign _6964 = _6431[4:4];
    assign _6961 = _6956 - _22192;
    assign _6962 = _6958 ? _6961 : _6956;
    assign _6963 = _6962[62:0];
    assign _6965 = { _6963,
                     _6964 };
    assign _6966 = _6965 < _22192;
    assign _6967 = ~ _6966;
    assign _6955 = _6431[5:5];
    assign _6952 = _6947 - _22192;
    assign _6953 = _6949 ? _6952 : _6947;
    assign _6954 = _6953[62:0];
    assign _6956 = { _6954,
                     _6955 };
    assign _6957 = _6956 < _22192;
    assign _6958 = ~ _6957;
    assign _6946 = _6431[6:6];
    assign _6943 = _6938 - _22192;
    assign _6944 = _6940 ? _6943 : _6938;
    assign _6945 = _6944[62:0];
    assign _6947 = { _6945,
                     _6946 };
    assign _6948 = _6947 < _22192;
    assign _6949 = ~ _6948;
    assign _6937 = _6431[7:7];
    assign _6934 = _6929 - _22192;
    assign _6935 = _6931 ? _6934 : _6929;
    assign _6936 = _6935[62:0];
    assign _6938 = { _6936,
                     _6937 };
    assign _6939 = _6938 < _22192;
    assign _6940 = ~ _6939;
    assign _6928 = _6431[8:8];
    assign _6925 = _6920 - _22192;
    assign _6926 = _6922 ? _6925 : _6920;
    assign _6927 = _6926[62:0];
    assign _6929 = { _6927,
                     _6928 };
    assign _6930 = _6929 < _22192;
    assign _6931 = ~ _6930;
    assign _6919 = _6431[9:9];
    assign _6916 = _6911 - _22192;
    assign _6917 = _6913 ? _6916 : _6911;
    assign _6918 = _6917[62:0];
    assign _6920 = { _6918,
                     _6919 };
    assign _6921 = _6920 < _22192;
    assign _6922 = ~ _6921;
    assign _6910 = _6431[10:10];
    assign _6907 = _6902 - _22192;
    assign _6908 = _6904 ? _6907 : _6902;
    assign _6909 = _6908[62:0];
    assign _6911 = { _6909,
                     _6910 };
    assign _6912 = _6911 < _22192;
    assign _6913 = ~ _6912;
    assign _6901 = _6431[11:11];
    assign _6898 = _6893 - _22192;
    assign _6899 = _6895 ? _6898 : _6893;
    assign _6900 = _6899[62:0];
    assign _6902 = { _6900,
                     _6901 };
    assign _6903 = _6902 < _22192;
    assign _6904 = ~ _6903;
    assign _6892 = _6431[12:12];
    assign _6889 = _6884 - _22192;
    assign _6890 = _6886 ? _6889 : _6884;
    assign _6891 = _6890[62:0];
    assign _6893 = { _6891,
                     _6892 };
    assign _6894 = _6893 < _22192;
    assign _6895 = ~ _6894;
    assign _6883 = _6431[13:13];
    assign _6880 = _6875 - _22192;
    assign _6881 = _6877 ? _6880 : _6875;
    assign _6882 = _6881[62:0];
    assign _6884 = { _6882,
                     _6883 };
    assign _6885 = _6884 < _22192;
    assign _6886 = ~ _6885;
    assign _6874 = _6431[14:14];
    assign _6871 = _6866 - _22192;
    assign _6872 = _6868 ? _6871 : _6866;
    assign _6873 = _6872[62:0];
    assign _6875 = { _6873,
                     _6874 };
    assign _6876 = _6875 < _22192;
    assign _6877 = ~ _6876;
    assign _6865 = _6431[15:15];
    assign _6862 = _6857 - _22192;
    assign _6863 = _6859 ? _6862 : _6857;
    assign _6864 = _6863[62:0];
    assign _6866 = { _6864,
                     _6865 };
    assign _6867 = _6866 < _22192;
    assign _6868 = ~ _6867;
    assign _6856 = _6431[16:16];
    assign _6853 = _6848 - _22192;
    assign _6854 = _6850 ? _6853 : _6848;
    assign _6855 = _6854[62:0];
    assign _6857 = { _6855,
                     _6856 };
    assign _6858 = _6857 < _22192;
    assign _6859 = ~ _6858;
    assign _6847 = _6431[17:17];
    assign _6844 = _6839 - _22192;
    assign _6845 = _6841 ? _6844 : _6839;
    assign _6846 = _6845[62:0];
    assign _6848 = { _6846,
                     _6847 };
    assign _6849 = _6848 < _22192;
    assign _6850 = ~ _6849;
    assign _6838 = _6431[18:18];
    assign _6835 = _6830 - _22192;
    assign _6836 = _6832 ? _6835 : _6830;
    assign _6837 = _6836[62:0];
    assign _6839 = { _6837,
                     _6838 };
    assign _6840 = _6839 < _22192;
    assign _6841 = ~ _6840;
    assign _6829 = _6431[19:19];
    assign _6826 = _6821 - _22192;
    assign _6827 = _6823 ? _6826 : _6821;
    assign _6828 = _6827[62:0];
    assign _6830 = { _6828,
                     _6829 };
    assign _6831 = _6830 < _22192;
    assign _6832 = ~ _6831;
    assign _6820 = _6431[20:20];
    assign _6817 = _6812 - _22192;
    assign _6818 = _6814 ? _6817 : _6812;
    assign _6819 = _6818[62:0];
    assign _6821 = { _6819,
                     _6820 };
    assign _6822 = _6821 < _22192;
    assign _6823 = ~ _6822;
    assign _6811 = _6431[21:21];
    assign _6808 = _6803 - _22192;
    assign _6809 = _6805 ? _6808 : _6803;
    assign _6810 = _6809[62:0];
    assign _6812 = { _6810,
                     _6811 };
    assign _6813 = _6812 < _22192;
    assign _6814 = ~ _6813;
    assign _6802 = _6431[22:22];
    assign _6799 = _6794 - _22192;
    assign _6800 = _6796 ? _6799 : _6794;
    assign _6801 = _6800[62:0];
    assign _6803 = { _6801,
                     _6802 };
    assign _6804 = _6803 < _22192;
    assign _6805 = ~ _6804;
    assign _6793 = _6431[23:23];
    assign _6790 = _6785 - _22192;
    assign _6791 = _6787 ? _6790 : _6785;
    assign _6792 = _6791[62:0];
    assign _6794 = { _6792,
                     _6793 };
    assign _6795 = _6794 < _22192;
    assign _6796 = ~ _6795;
    assign _6784 = _6431[24:24];
    assign _6781 = _6776 - _22192;
    assign _6782 = _6778 ? _6781 : _6776;
    assign _6783 = _6782[62:0];
    assign _6785 = { _6783,
                     _6784 };
    assign _6786 = _6785 < _22192;
    assign _6787 = ~ _6786;
    assign _6775 = _6431[25:25];
    assign _6772 = _6767 - _22192;
    assign _6773 = _6769 ? _6772 : _6767;
    assign _6774 = _6773[62:0];
    assign _6776 = { _6774,
                     _6775 };
    assign _6777 = _6776 < _22192;
    assign _6778 = ~ _6777;
    assign _6766 = _6431[26:26];
    assign _6763 = _6758 - _22192;
    assign _6764 = _6760 ? _6763 : _6758;
    assign _6765 = _6764[62:0];
    assign _6767 = { _6765,
                     _6766 };
    assign _6768 = _6767 < _22192;
    assign _6769 = ~ _6768;
    assign _6757 = _6431[27:27];
    assign _6754 = _6749 - _22192;
    assign _6755 = _6751 ? _6754 : _6749;
    assign _6756 = _6755[62:0];
    assign _6758 = { _6756,
                     _6757 };
    assign _6759 = _6758 < _22192;
    assign _6760 = ~ _6759;
    assign _6748 = _6431[28:28];
    assign _6745 = _6740 - _22192;
    assign _6746 = _6742 ? _6745 : _6740;
    assign _6747 = _6746[62:0];
    assign _6749 = { _6747,
                     _6748 };
    assign _6750 = _6749 < _22192;
    assign _6751 = ~ _6750;
    assign _6739 = _6431[29:29];
    assign _6736 = _6731 - _22192;
    assign _6737 = _6733 ? _6736 : _6731;
    assign _6738 = _6737[62:0];
    assign _6740 = { _6738,
                     _6739 };
    assign _6741 = _6740 < _22192;
    assign _6742 = ~ _6741;
    assign _6730 = _6431[30:30];
    assign _6727 = _6722 - _22192;
    assign _6728 = _6724 ? _6727 : _6722;
    assign _6729 = _6728[62:0];
    assign _6731 = { _6729,
                     _6730 };
    assign _6732 = _6731 < _22192;
    assign _6733 = ~ _6732;
    assign _6721 = _6431[31:31];
    assign _6718 = _6713 - _22192;
    assign _6719 = _6715 ? _6718 : _6713;
    assign _6720 = _6719[62:0];
    assign _6722 = { _6720,
                     _6721 };
    assign _6723 = _6722 < _22192;
    assign _6724 = ~ _6723;
    assign _6712 = _6431[32:32];
    assign _6709 = _6704 - _22192;
    assign _6710 = _6706 ? _6709 : _6704;
    assign _6711 = _6710[62:0];
    assign _6713 = { _6711,
                     _6712 };
    assign _6714 = _6713 < _22192;
    assign _6715 = ~ _6714;
    assign _6703 = _6431[33:33];
    assign _6700 = _6695 - _22192;
    assign _6701 = _6697 ? _6700 : _6695;
    assign _6702 = _6701[62:0];
    assign _6704 = { _6702,
                     _6703 };
    assign _6705 = _6704 < _22192;
    assign _6706 = ~ _6705;
    assign _6694 = _6431[34:34];
    assign _6691 = _6686 - _22192;
    assign _6692 = _6688 ? _6691 : _6686;
    assign _6693 = _6692[62:0];
    assign _6695 = { _6693,
                     _6694 };
    assign _6696 = _6695 < _22192;
    assign _6697 = ~ _6696;
    assign _6685 = _6431[35:35];
    assign _6682 = _6677 - _22192;
    assign _6683 = _6679 ? _6682 : _6677;
    assign _6684 = _6683[62:0];
    assign _6686 = { _6684,
                     _6685 };
    assign _6687 = _6686 < _22192;
    assign _6688 = ~ _6687;
    assign _6676 = _6431[36:36];
    assign _6673 = _6668 - _22192;
    assign _6674 = _6670 ? _6673 : _6668;
    assign _6675 = _6674[62:0];
    assign _6677 = { _6675,
                     _6676 };
    assign _6678 = _6677 < _22192;
    assign _6679 = ~ _6678;
    assign _6667 = _6431[37:37];
    assign _6664 = _6659 - _22192;
    assign _6665 = _6661 ? _6664 : _6659;
    assign _6666 = _6665[62:0];
    assign _6668 = { _6666,
                     _6667 };
    assign _6669 = _6668 < _22192;
    assign _6670 = ~ _6669;
    assign _6658 = _6431[38:38];
    assign _6655 = _6650 - _22192;
    assign _6656 = _6652 ? _6655 : _6650;
    assign _6657 = _6656[62:0];
    assign _6659 = { _6657,
                     _6658 };
    assign _6660 = _6659 < _22192;
    assign _6661 = ~ _6660;
    assign _6649 = _6431[39:39];
    assign _6646 = _6641 - _22192;
    assign _6647 = _6643 ? _6646 : _6641;
    assign _6648 = _6647[62:0];
    assign _6650 = { _6648,
                     _6649 };
    assign _6651 = _6650 < _22192;
    assign _6652 = ~ _6651;
    assign _6640 = _6431[40:40];
    assign _6637 = _6632 - _22192;
    assign _6638 = _6634 ? _6637 : _6632;
    assign _6639 = _6638[62:0];
    assign _6641 = { _6639,
                     _6640 };
    assign _6642 = _6641 < _22192;
    assign _6643 = ~ _6642;
    assign _6631 = _6431[41:41];
    assign _6628 = _6623 - _22192;
    assign _6629 = _6625 ? _6628 : _6623;
    assign _6630 = _6629[62:0];
    assign _6632 = { _6630,
                     _6631 };
    assign _6633 = _6632 < _22192;
    assign _6634 = ~ _6633;
    assign _6622 = _6431[42:42];
    assign _6619 = _6614 - _22192;
    assign _6620 = _6616 ? _6619 : _6614;
    assign _6621 = _6620[62:0];
    assign _6623 = { _6621,
                     _6622 };
    assign _6624 = _6623 < _22192;
    assign _6625 = ~ _6624;
    assign _6613 = _6431[43:43];
    assign _6610 = _6605 - _22192;
    assign _6611 = _6607 ? _6610 : _6605;
    assign _6612 = _6611[62:0];
    assign _6614 = { _6612,
                     _6613 };
    assign _6615 = _6614 < _22192;
    assign _6616 = ~ _6615;
    assign _6604 = _6431[44:44];
    assign _6601 = _6596 - _22192;
    assign _6602 = _6598 ? _6601 : _6596;
    assign _6603 = _6602[62:0];
    assign _6605 = { _6603,
                     _6604 };
    assign _6606 = _6605 < _22192;
    assign _6607 = ~ _6606;
    assign _6595 = _6431[45:45];
    assign _6592 = _6587 - _22192;
    assign _6593 = _6589 ? _6592 : _6587;
    assign _6594 = _6593[62:0];
    assign _6596 = { _6594,
                     _6595 };
    assign _6597 = _6596 < _22192;
    assign _6598 = ~ _6597;
    assign _6586 = _6431[46:46];
    assign _6583 = _6578 - _22192;
    assign _6584 = _6580 ? _6583 : _6578;
    assign _6585 = _6584[62:0];
    assign _6587 = { _6585,
                     _6586 };
    assign _6588 = _6587 < _22192;
    assign _6589 = ~ _6588;
    assign _6577 = _6431[47:47];
    assign _6574 = _6569 - _22192;
    assign _6575 = _6571 ? _6574 : _6569;
    assign _6576 = _6575[62:0];
    assign _6578 = { _6576,
                     _6577 };
    assign _6579 = _6578 < _22192;
    assign _6580 = ~ _6579;
    assign _6568 = _6431[48:48];
    assign _6565 = _6560 - _22192;
    assign _6566 = _6562 ? _6565 : _6560;
    assign _6567 = _6566[62:0];
    assign _6569 = { _6567,
                     _6568 };
    assign _6570 = _6569 < _22192;
    assign _6571 = ~ _6570;
    assign _6559 = _6431[49:49];
    assign _6556 = _6551 - _22192;
    assign _6557 = _6553 ? _6556 : _6551;
    assign _6558 = _6557[62:0];
    assign _6560 = { _6558,
                     _6559 };
    assign _6561 = _6560 < _22192;
    assign _6562 = ~ _6561;
    assign _6550 = _6431[50:50];
    assign _6547 = _6542 - _22192;
    assign _6548 = _6544 ? _6547 : _6542;
    assign _6549 = _6548[62:0];
    assign _6551 = { _6549,
                     _6550 };
    assign _6552 = _6551 < _22192;
    assign _6553 = ~ _6552;
    assign _6541 = _6431[51:51];
    assign _6538 = _6533 - _22192;
    assign _6539 = _6535 ? _6538 : _6533;
    assign _6540 = _6539[62:0];
    assign _6542 = { _6540,
                     _6541 };
    assign _6543 = _6542 < _22192;
    assign _6544 = ~ _6543;
    assign _6532 = _6431[52:52];
    assign _6529 = _6524 - _22192;
    assign _6530 = _6526 ? _6529 : _6524;
    assign _6531 = _6530[62:0];
    assign _6533 = { _6531,
                     _6532 };
    assign _6534 = _6533 < _22192;
    assign _6535 = ~ _6534;
    assign _6523 = _6431[53:53];
    assign _6520 = _6515 - _22192;
    assign _6521 = _6517 ? _6520 : _6515;
    assign _6522 = _6521[62:0];
    assign _6524 = { _6522,
                     _6523 };
    assign _6525 = _6524 < _22192;
    assign _6526 = ~ _6525;
    assign _6514 = _6431[54:54];
    assign _6511 = _6506 - _22192;
    assign _6512 = _6508 ? _6511 : _6506;
    assign _6513 = _6512[62:0];
    assign _6515 = { _6513,
                     _6514 };
    assign _6516 = _6515 < _22192;
    assign _6517 = ~ _6516;
    assign _6505 = _6431[55:55];
    assign _6502 = _6497 - _22192;
    assign _6503 = _6499 ? _6502 : _6497;
    assign _6504 = _6503[62:0];
    assign _6506 = { _6504,
                     _6505 };
    assign _6507 = _6506 < _22192;
    assign _6508 = ~ _6507;
    assign _6496 = _6431[56:56];
    assign _6493 = _6488 - _22192;
    assign _6494 = _6490 ? _6493 : _6488;
    assign _6495 = _6494[62:0];
    assign _6497 = { _6495,
                     _6496 };
    assign _6498 = _6497 < _22192;
    assign _6499 = ~ _6498;
    assign _6487 = _6431[57:57];
    assign _6484 = _6479 - _22192;
    assign _6485 = _6481 ? _6484 : _6479;
    assign _6486 = _6485[62:0];
    assign _6488 = { _6486,
                     _6487 };
    assign _6489 = _6488 < _22192;
    assign _6490 = ~ _6489;
    assign _6478 = _6431[58:58];
    assign _6475 = _6470 - _22192;
    assign _6476 = _6472 ? _6475 : _6470;
    assign _6477 = _6476[62:0];
    assign _6479 = { _6477,
                     _6478 };
    assign _6480 = _6479 < _22192;
    assign _6481 = ~ _6480;
    assign _6469 = _6431[59:59];
    assign _6466 = _6461 - _22192;
    assign _6467 = _6463 ? _6466 : _6461;
    assign _6468 = _6467[62:0];
    assign _6470 = { _6468,
                     _6469 };
    assign _6471 = _6470 < _22192;
    assign _6472 = ~ _6471;
    assign _6460 = _6431[60:60];
    assign _6457 = _6452 - _22192;
    assign _6458 = _6454 ? _6457 : _6452;
    assign _6459 = _6458[62:0];
    assign _6461 = { _6459,
                     _6460 };
    assign _6462 = _6461 < _22192;
    assign _6463 = ~ _6462;
    assign _6451 = _6431[61:61];
    assign _6448 = _6443 - _22192;
    assign _6449 = _6445 ? _6448 : _6443;
    assign _6450 = _6449[62:0];
    assign _6452 = { _6450,
                     _6451 };
    assign _6453 = _6452 < _22192;
    assign _6454 = ~ _6453;
    assign _6442 = _6431[62:62];
    assign _6439 = _6433 - _22192;
    assign _6440 = _6436 ? _6439 : _6433;
    assign _6441 = _6440[62:0];
    assign _6443 = { _6441,
                     _6442 };
    assign _6444 = _6443 < _22192;
    assign _6445 = ~ _6444;
    assign _6429 = _6421 + _22186;
    assign _6430 = _6421 * _6429;
    assign _6431 = _6430[63:0];
    assign _6432 = _6431[63:63];
    assign _6433 = { _22185,
                     _6432 };
    assign _6435 = _6433 < _22192;
    assign _6436 = ~ _6435;
    assign _6437 = { _22185,
                     _6436 };
    assign _6438 = _6437[62:0];
    assign _6446 = { _6438,
                     _6445 };
    assign _6447 = _6446[62:0];
    assign _6455 = { _6447,
                     _6454 };
    assign _6456 = _6455[62:0];
    assign _6464 = { _6456,
                     _6463 };
    assign _6465 = _6464[62:0];
    assign _6473 = { _6465,
                     _6472 };
    assign _6474 = _6473[62:0];
    assign _6482 = { _6474,
                     _6481 };
    assign _6483 = _6482[62:0];
    assign _6491 = { _6483,
                     _6490 };
    assign _6492 = _6491[62:0];
    assign _6500 = { _6492,
                     _6499 };
    assign _6501 = _6500[62:0];
    assign _6509 = { _6501,
                     _6508 };
    assign _6510 = _6509[62:0];
    assign _6518 = { _6510,
                     _6517 };
    assign _6519 = _6518[62:0];
    assign _6527 = { _6519,
                     _6526 };
    assign _6528 = _6527[62:0];
    assign _6536 = { _6528,
                     _6535 };
    assign _6537 = _6536[62:0];
    assign _6545 = { _6537,
                     _6544 };
    assign _6546 = _6545[62:0];
    assign _6554 = { _6546,
                     _6553 };
    assign _6555 = _6554[62:0];
    assign _6563 = { _6555,
                     _6562 };
    assign _6564 = _6563[62:0];
    assign _6572 = { _6564,
                     _6571 };
    assign _6573 = _6572[62:0];
    assign _6581 = { _6573,
                     _6580 };
    assign _6582 = _6581[62:0];
    assign _6590 = { _6582,
                     _6589 };
    assign _6591 = _6590[62:0];
    assign _6599 = { _6591,
                     _6598 };
    assign _6600 = _6599[62:0];
    assign _6608 = { _6600,
                     _6607 };
    assign _6609 = _6608[62:0];
    assign _6617 = { _6609,
                     _6616 };
    assign _6618 = _6617[62:0];
    assign _6626 = { _6618,
                     _6625 };
    assign _6627 = _6626[62:0];
    assign _6635 = { _6627,
                     _6634 };
    assign _6636 = _6635[62:0];
    assign _6644 = { _6636,
                     _6643 };
    assign _6645 = _6644[62:0];
    assign _6653 = { _6645,
                     _6652 };
    assign _6654 = _6653[62:0];
    assign _6662 = { _6654,
                     _6661 };
    assign _6663 = _6662[62:0];
    assign _6671 = { _6663,
                     _6670 };
    assign _6672 = _6671[62:0];
    assign _6680 = { _6672,
                     _6679 };
    assign _6681 = _6680[62:0];
    assign _6689 = { _6681,
                     _6688 };
    assign _6690 = _6689[62:0];
    assign _6698 = { _6690,
                     _6697 };
    assign _6699 = _6698[62:0];
    assign _6707 = { _6699,
                     _6706 };
    assign _6708 = _6707[62:0];
    assign _6716 = { _6708,
                     _6715 };
    assign _6717 = _6716[62:0];
    assign _6725 = { _6717,
                     _6724 };
    assign _6726 = _6725[62:0];
    assign _6734 = { _6726,
                     _6733 };
    assign _6735 = _6734[62:0];
    assign _6743 = { _6735,
                     _6742 };
    assign _6744 = _6743[62:0];
    assign _6752 = { _6744,
                     _6751 };
    assign _6753 = _6752[62:0];
    assign _6761 = { _6753,
                     _6760 };
    assign _6762 = _6761[62:0];
    assign _6770 = { _6762,
                     _6769 };
    assign _6771 = _6770[62:0];
    assign _6779 = { _6771,
                     _6778 };
    assign _6780 = _6779[62:0];
    assign _6788 = { _6780,
                     _6787 };
    assign _6789 = _6788[62:0];
    assign _6797 = { _6789,
                     _6796 };
    assign _6798 = _6797[62:0];
    assign _6806 = { _6798,
                     _6805 };
    assign _6807 = _6806[62:0];
    assign _6815 = { _6807,
                     _6814 };
    assign _6816 = _6815[62:0];
    assign _6824 = { _6816,
                     _6823 };
    assign _6825 = _6824[62:0];
    assign _6833 = { _6825,
                     _6832 };
    assign _6834 = _6833[62:0];
    assign _6842 = { _6834,
                     _6841 };
    assign _6843 = _6842[62:0];
    assign _6851 = { _6843,
                     _6850 };
    assign _6852 = _6851[62:0];
    assign _6860 = { _6852,
                     _6859 };
    assign _6861 = _6860[62:0];
    assign _6869 = { _6861,
                     _6868 };
    assign _6870 = _6869[62:0];
    assign _6878 = { _6870,
                     _6877 };
    assign _6879 = _6878[62:0];
    assign _6887 = { _6879,
                     _6886 };
    assign _6888 = _6887[62:0];
    assign _6896 = { _6888,
                     _6895 };
    assign _6897 = _6896[62:0];
    assign _6905 = { _6897,
                     _6904 };
    assign _6906 = _6905[62:0];
    assign _6914 = { _6906,
                     _6913 };
    assign _6915 = _6914[62:0];
    assign _6923 = { _6915,
                     _6922 };
    assign _6924 = _6923[62:0];
    assign _6932 = { _6924,
                     _6931 };
    assign _6933 = _6932[62:0];
    assign _6941 = { _6933,
                     _6940 };
    assign _6942 = _6941[62:0];
    assign _6950 = { _6942,
                     _6949 };
    assign _6951 = _6950[62:0];
    assign _6959 = { _6951,
                     _6958 };
    assign _6960 = _6959[62:0];
    assign _6968 = { _6960,
                     _6967 };
    assign _6969 = _6968[62:0];
    assign _6977 = { _6969,
                     _6976 };
    assign _6978 = _6977[62:0];
    assign _6986 = { _6978,
                     _6985 };
    assign _6987 = _6986[62:0];
    assign _6995 = { _6987,
                     _6994 };
    assign _6996 = _6995[62:0];
    assign _7004 = { _6996,
                     _7003 };
    assign _7005 = _5269 * _7004;
    assign _7006 = _7005[63:0];
    assign _6417 = _5849[0:0];
    assign _6414 = _6409 - _5269;
    assign _6415 = _6411 ? _6414 : _6409;
    assign _6416 = _6415[62:0];
    assign _6418 = { _6416,
                     _6417 };
    assign _6419 = _6418 < _5269;
    assign _6420 = ~ _6419;
    assign _6408 = _5849[1:1];
    assign _6405 = _6400 - _5269;
    assign _6406 = _6402 ? _6405 : _6400;
    assign _6407 = _6406[62:0];
    assign _6409 = { _6407,
                     _6408 };
    assign _6410 = _6409 < _5269;
    assign _6411 = ~ _6410;
    assign _6399 = _5849[2:2];
    assign _6396 = _6391 - _5269;
    assign _6397 = _6393 ? _6396 : _6391;
    assign _6398 = _6397[62:0];
    assign _6400 = { _6398,
                     _6399 };
    assign _6401 = _6400 < _5269;
    assign _6402 = ~ _6401;
    assign _6390 = _5849[3:3];
    assign _6387 = _6382 - _5269;
    assign _6388 = _6384 ? _6387 : _6382;
    assign _6389 = _6388[62:0];
    assign _6391 = { _6389,
                     _6390 };
    assign _6392 = _6391 < _5269;
    assign _6393 = ~ _6392;
    assign _6381 = _5849[4:4];
    assign _6378 = _6373 - _5269;
    assign _6379 = _6375 ? _6378 : _6373;
    assign _6380 = _6379[62:0];
    assign _6382 = { _6380,
                     _6381 };
    assign _6383 = _6382 < _5269;
    assign _6384 = ~ _6383;
    assign _6372 = _5849[5:5];
    assign _6369 = _6364 - _5269;
    assign _6370 = _6366 ? _6369 : _6364;
    assign _6371 = _6370[62:0];
    assign _6373 = { _6371,
                     _6372 };
    assign _6374 = _6373 < _5269;
    assign _6375 = ~ _6374;
    assign _6363 = _5849[6:6];
    assign _6360 = _6355 - _5269;
    assign _6361 = _6357 ? _6360 : _6355;
    assign _6362 = _6361[62:0];
    assign _6364 = { _6362,
                     _6363 };
    assign _6365 = _6364 < _5269;
    assign _6366 = ~ _6365;
    assign _6354 = _5849[7:7];
    assign _6351 = _6346 - _5269;
    assign _6352 = _6348 ? _6351 : _6346;
    assign _6353 = _6352[62:0];
    assign _6355 = { _6353,
                     _6354 };
    assign _6356 = _6355 < _5269;
    assign _6357 = ~ _6356;
    assign _6345 = _5849[8:8];
    assign _6342 = _6337 - _5269;
    assign _6343 = _6339 ? _6342 : _6337;
    assign _6344 = _6343[62:0];
    assign _6346 = { _6344,
                     _6345 };
    assign _6347 = _6346 < _5269;
    assign _6348 = ~ _6347;
    assign _6336 = _5849[9:9];
    assign _6333 = _6328 - _5269;
    assign _6334 = _6330 ? _6333 : _6328;
    assign _6335 = _6334[62:0];
    assign _6337 = { _6335,
                     _6336 };
    assign _6338 = _6337 < _5269;
    assign _6339 = ~ _6338;
    assign _6327 = _5849[10:10];
    assign _6324 = _6319 - _5269;
    assign _6325 = _6321 ? _6324 : _6319;
    assign _6326 = _6325[62:0];
    assign _6328 = { _6326,
                     _6327 };
    assign _6329 = _6328 < _5269;
    assign _6330 = ~ _6329;
    assign _6318 = _5849[11:11];
    assign _6315 = _6310 - _5269;
    assign _6316 = _6312 ? _6315 : _6310;
    assign _6317 = _6316[62:0];
    assign _6319 = { _6317,
                     _6318 };
    assign _6320 = _6319 < _5269;
    assign _6321 = ~ _6320;
    assign _6309 = _5849[12:12];
    assign _6306 = _6301 - _5269;
    assign _6307 = _6303 ? _6306 : _6301;
    assign _6308 = _6307[62:0];
    assign _6310 = { _6308,
                     _6309 };
    assign _6311 = _6310 < _5269;
    assign _6312 = ~ _6311;
    assign _6300 = _5849[13:13];
    assign _6297 = _6292 - _5269;
    assign _6298 = _6294 ? _6297 : _6292;
    assign _6299 = _6298[62:0];
    assign _6301 = { _6299,
                     _6300 };
    assign _6302 = _6301 < _5269;
    assign _6303 = ~ _6302;
    assign _6291 = _5849[14:14];
    assign _6288 = _6283 - _5269;
    assign _6289 = _6285 ? _6288 : _6283;
    assign _6290 = _6289[62:0];
    assign _6292 = { _6290,
                     _6291 };
    assign _6293 = _6292 < _5269;
    assign _6294 = ~ _6293;
    assign _6282 = _5849[15:15];
    assign _6279 = _6274 - _5269;
    assign _6280 = _6276 ? _6279 : _6274;
    assign _6281 = _6280[62:0];
    assign _6283 = { _6281,
                     _6282 };
    assign _6284 = _6283 < _5269;
    assign _6285 = ~ _6284;
    assign _6273 = _5849[16:16];
    assign _6270 = _6265 - _5269;
    assign _6271 = _6267 ? _6270 : _6265;
    assign _6272 = _6271[62:0];
    assign _6274 = { _6272,
                     _6273 };
    assign _6275 = _6274 < _5269;
    assign _6276 = ~ _6275;
    assign _6264 = _5849[17:17];
    assign _6261 = _6256 - _5269;
    assign _6262 = _6258 ? _6261 : _6256;
    assign _6263 = _6262[62:0];
    assign _6265 = { _6263,
                     _6264 };
    assign _6266 = _6265 < _5269;
    assign _6267 = ~ _6266;
    assign _6255 = _5849[18:18];
    assign _6252 = _6247 - _5269;
    assign _6253 = _6249 ? _6252 : _6247;
    assign _6254 = _6253[62:0];
    assign _6256 = { _6254,
                     _6255 };
    assign _6257 = _6256 < _5269;
    assign _6258 = ~ _6257;
    assign _6246 = _5849[19:19];
    assign _6243 = _6238 - _5269;
    assign _6244 = _6240 ? _6243 : _6238;
    assign _6245 = _6244[62:0];
    assign _6247 = { _6245,
                     _6246 };
    assign _6248 = _6247 < _5269;
    assign _6249 = ~ _6248;
    assign _6237 = _5849[20:20];
    assign _6234 = _6229 - _5269;
    assign _6235 = _6231 ? _6234 : _6229;
    assign _6236 = _6235[62:0];
    assign _6238 = { _6236,
                     _6237 };
    assign _6239 = _6238 < _5269;
    assign _6240 = ~ _6239;
    assign _6228 = _5849[21:21];
    assign _6225 = _6220 - _5269;
    assign _6226 = _6222 ? _6225 : _6220;
    assign _6227 = _6226[62:0];
    assign _6229 = { _6227,
                     _6228 };
    assign _6230 = _6229 < _5269;
    assign _6231 = ~ _6230;
    assign _6219 = _5849[22:22];
    assign _6216 = _6211 - _5269;
    assign _6217 = _6213 ? _6216 : _6211;
    assign _6218 = _6217[62:0];
    assign _6220 = { _6218,
                     _6219 };
    assign _6221 = _6220 < _5269;
    assign _6222 = ~ _6221;
    assign _6210 = _5849[23:23];
    assign _6207 = _6202 - _5269;
    assign _6208 = _6204 ? _6207 : _6202;
    assign _6209 = _6208[62:0];
    assign _6211 = { _6209,
                     _6210 };
    assign _6212 = _6211 < _5269;
    assign _6213 = ~ _6212;
    assign _6201 = _5849[24:24];
    assign _6198 = _6193 - _5269;
    assign _6199 = _6195 ? _6198 : _6193;
    assign _6200 = _6199[62:0];
    assign _6202 = { _6200,
                     _6201 };
    assign _6203 = _6202 < _5269;
    assign _6204 = ~ _6203;
    assign _6192 = _5849[25:25];
    assign _6189 = _6184 - _5269;
    assign _6190 = _6186 ? _6189 : _6184;
    assign _6191 = _6190[62:0];
    assign _6193 = { _6191,
                     _6192 };
    assign _6194 = _6193 < _5269;
    assign _6195 = ~ _6194;
    assign _6183 = _5849[26:26];
    assign _6180 = _6175 - _5269;
    assign _6181 = _6177 ? _6180 : _6175;
    assign _6182 = _6181[62:0];
    assign _6184 = { _6182,
                     _6183 };
    assign _6185 = _6184 < _5269;
    assign _6186 = ~ _6185;
    assign _6174 = _5849[27:27];
    assign _6171 = _6166 - _5269;
    assign _6172 = _6168 ? _6171 : _6166;
    assign _6173 = _6172[62:0];
    assign _6175 = { _6173,
                     _6174 };
    assign _6176 = _6175 < _5269;
    assign _6177 = ~ _6176;
    assign _6165 = _5849[28:28];
    assign _6162 = _6157 - _5269;
    assign _6163 = _6159 ? _6162 : _6157;
    assign _6164 = _6163[62:0];
    assign _6166 = { _6164,
                     _6165 };
    assign _6167 = _6166 < _5269;
    assign _6168 = ~ _6167;
    assign _6156 = _5849[29:29];
    assign _6153 = _6148 - _5269;
    assign _6154 = _6150 ? _6153 : _6148;
    assign _6155 = _6154[62:0];
    assign _6157 = { _6155,
                     _6156 };
    assign _6158 = _6157 < _5269;
    assign _6159 = ~ _6158;
    assign _6147 = _5849[30:30];
    assign _6144 = _6139 - _5269;
    assign _6145 = _6141 ? _6144 : _6139;
    assign _6146 = _6145[62:0];
    assign _6148 = { _6146,
                     _6147 };
    assign _6149 = _6148 < _5269;
    assign _6150 = ~ _6149;
    assign _6138 = _5849[31:31];
    assign _6135 = _6130 - _5269;
    assign _6136 = _6132 ? _6135 : _6130;
    assign _6137 = _6136[62:0];
    assign _6139 = { _6137,
                     _6138 };
    assign _6140 = _6139 < _5269;
    assign _6141 = ~ _6140;
    assign _6129 = _5849[32:32];
    assign _6126 = _6121 - _5269;
    assign _6127 = _6123 ? _6126 : _6121;
    assign _6128 = _6127[62:0];
    assign _6130 = { _6128,
                     _6129 };
    assign _6131 = _6130 < _5269;
    assign _6132 = ~ _6131;
    assign _6120 = _5849[33:33];
    assign _6117 = _6112 - _5269;
    assign _6118 = _6114 ? _6117 : _6112;
    assign _6119 = _6118[62:0];
    assign _6121 = { _6119,
                     _6120 };
    assign _6122 = _6121 < _5269;
    assign _6123 = ~ _6122;
    assign _6111 = _5849[34:34];
    assign _6108 = _6103 - _5269;
    assign _6109 = _6105 ? _6108 : _6103;
    assign _6110 = _6109[62:0];
    assign _6112 = { _6110,
                     _6111 };
    assign _6113 = _6112 < _5269;
    assign _6114 = ~ _6113;
    assign _6102 = _5849[35:35];
    assign _6099 = _6094 - _5269;
    assign _6100 = _6096 ? _6099 : _6094;
    assign _6101 = _6100[62:0];
    assign _6103 = { _6101,
                     _6102 };
    assign _6104 = _6103 < _5269;
    assign _6105 = ~ _6104;
    assign _6093 = _5849[36:36];
    assign _6090 = _6085 - _5269;
    assign _6091 = _6087 ? _6090 : _6085;
    assign _6092 = _6091[62:0];
    assign _6094 = { _6092,
                     _6093 };
    assign _6095 = _6094 < _5269;
    assign _6096 = ~ _6095;
    assign _6084 = _5849[37:37];
    assign _6081 = _6076 - _5269;
    assign _6082 = _6078 ? _6081 : _6076;
    assign _6083 = _6082[62:0];
    assign _6085 = { _6083,
                     _6084 };
    assign _6086 = _6085 < _5269;
    assign _6087 = ~ _6086;
    assign _6075 = _5849[38:38];
    assign _6072 = _6067 - _5269;
    assign _6073 = _6069 ? _6072 : _6067;
    assign _6074 = _6073[62:0];
    assign _6076 = { _6074,
                     _6075 };
    assign _6077 = _6076 < _5269;
    assign _6078 = ~ _6077;
    assign _6066 = _5849[39:39];
    assign _6063 = _6058 - _5269;
    assign _6064 = _6060 ? _6063 : _6058;
    assign _6065 = _6064[62:0];
    assign _6067 = { _6065,
                     _6066 };
    assign _6068 = _6067 < _5269;
    assign _6069 = ~ _6068;
    assign _6057 = _5849[40:40];
    assign _6054 = _6049 - _5269;
    assign _6055 = _6051 ? _6054 : _6049;
    assign _6056 = _6055[62:0];
    assign _6058 = { _6056,
                     _6057 };
    assign _6059 = _6058 < _5269;
    assign _6060 = ~ _6059;
    assign _6048 = _5849[41:41];
    assign _6045 = _6040 - _5269;
    assign _6046 = _6042 ? _6045 : _6040;
    assign _6047 = _6046[62:0];
    assign _6049 = { _6047,
                     _6048 };
    assign _6050 = _6049 < _5269;
    assign _6051 = ~ _6050;
    assign _6039 = _5849[42:42];
    assign _6036 = _6031 - _5269;
    assign _6037 = _6033 ? _6036 : _6031;
    assign _6038 = _6037[62:0];
    assign _6040 = { _6038,
                     _6039 };
    assign _6041 = _6040 < _5269;
    assign _6042 = ~ _6041;
    assign _6030 = _5849[43:43];
    assign _6027 = _6022 - _5269;
    assign _6028 = _6024 ? _6027 : _6022;
    assign _6029 = _6028[62:0];
    assign _6031 = { _6029,
                     _6030 };
    assign _6032 = _6031 < _5269;
    assign _6033 = ~ _6032;
    assign _6021 = _5849[44:44];
    assign _6018 = _6013 - _5269;
    assign _6019 = _6015 ? _6018 : _6013;
    assign _6020 = _6019[62:0];
    assign _6022 = { _6020,
                     _6021 };
    assign _6023 = _6022 < _5269;
    assign _6024 = ~ _6023;
    assign _6012 = _5849[45:45];
    assign _6009 = _6004 - _5269;
    assign _6010 = _6006 ? _6009 : _6004;
    assign _6011 = _6010[62:0];
    assign _6013 = { _6011,
                     _6012 };
    assign _6014 = _6013 < _5269;
    assign _6015 = ~ _6014;
    assign _6003 = _5849[46:46];
    assign _6000 = _5995 - _5269;
    assign _6001 = _5997 ? _6000 : _5995;
    assign _6002 = _6001[62:0];
    assign _6004 = { _6002,
                     _6003 };
    assign _6005 = _6004 < _5269;
    assign _6006 = ~ _6005;
    assign _5994 = _5849[47:47];
    assign _5991 = _5986 - _5269;
    assign _5992 = _5988 ? _5991 : _5986;
    assign _5993 = _5992[62:0];
    assign _5995 = { _5993,
                     _5994 };
    assign _5996 = _5995 < _5269;
    assign _5997 = ~ _5996;
    assign _5985 = _5849[48:48];
    assign _5982 = _5977 - _5269;
    assign _5983 = _5979 ? _5982 : _5977;
    assign _5984 = _5983[62:0];
    assign _5986 = { _5984,
                     _5985 };
    assign _5987 = _5986 < _5269;
    assign _5988 = ~ _5987;
    assign _5976 = _5849[49:49];
    assign _5973 = _5968 - _5269;
    assign _5974 = _5970 ? _5973 : _5968;
    assign _5975 = _5974[62:0];
    assign _5977 = { _5975,
                     _5976 };
    assign _5978 = _5977 < _5269;
    assign _5979 = ~ _5978;
    assign _5967 = _5849[50:50];
    assign _5964 = _5959 - _5269;
    assign _5965 = _5961 ? _5964 : _5959;
    assign _5966 = _5965[62:0];
    assign _5968 = { _5966,
                     _5967 };
    assign _5969 = _5968 < _5269;
    assign _5970 = ~ _5969;
    assign _5958 = _5849[51:51];
    assign _5955 = _5950 - _5269;
    assign _5956 = _5952 ? _5955 : _5950;
    assign _5957 = _5956[62:0];
    assign _5959 = { _5957,
                     _5958 };
    assign _5960 = _5959 < _5269;
    assign _5961 = ~ _5960;
    assign _5949 = _5849[52:52];
    assign _5946 = _5941 - _5269;
    assign _5947 = _5943 ? _5946 : _5941;
    assign _5948 = _5947[62:0];
    assign _5950 = { _5948,
                     _5949 };
    assign _5951 = _5950 < _5269;
    assign _5952 = ~ _5951;
    assign _5940 = _5849[53:53];
    assign _5937 = _5932 - _5269;
    assign _5938 = _5934 ? _5937 : _5932;
    assign _5939 = _5938[62:0];
    assign _5941 = { _5939,
                     _5940 };
    assign _5942 = _5941 < _5269;
    assign _5943 = ~ _5942;
    assign _5931 = _5849[54:54];
    assign _5928 = _5923 - _5269;
    assign _5929 = _5925 ? _5928 : _5923;
    assign _5930 = _5929[62:0];
    assign _5932 = { _5930,
                     _5931 };
    assign _5933 = _5932 < _5269;
    assign _5934 = ~ _5933;
    assign _5922 = _5849[55:55];
    assign _5919 = _5914 - _5269;
    assign _5920 = _5916 ? _5919 : _5914;
    assign _5921 = _5920[62:0];
    assign _5923 = { _5921,
                     _5922 };
    assign _5924 = _5923 < _5269;
    assign _5925 = ~ _5924;
    assign _5913 = _5849[56:56];
    assign _5910 = _5905 - _5269;
    assign _5911 = _5907 ? _5910 : _5905;
    assign _5912 = _5911[62:0];
    assign _5914 = { _5912,
                     _5913 };
    assign _5915 = _5914 < _5269;
    assign _5916 = ~ _5915;
    assign _5904 = _5849[57:57];
    assign _5901 = _5896 - _5269;
    assign _5902 = _5898 ? _5901 : _5896;
    assign _5903 = _5902[62:0];
    assign _5905 = { _5903,
                     _5904 };
    assign _5906 = _5905 < _5269;
    assign _5907 = ~ _5906;
    assign _5895 = _5849[58:58];
    assign _5892 = _5887 - _5269;
    assign _5893 = _5889 ? _5892 : _5887;
    assign _5894 = _5893[62:0];
    assign _5896 = { _5894,
                     _5895 };
    assign _5897 = _5896 < _5269;
    assign _5898 = ~ _5897;
    assign _5886 = _5849[59:59];
    assign _5883 = _5878 - _5269;
    assign _5884 = _5880 ? _5883 : _5878;
    assign _5885 = _5884[62:0];
    assign _5887 = { _5885,
                     _5886 };
    assign _5888 = _5887 < _5269;
    assign _5889 = ~ _5888;
    assign _5877 = _5849[60:60];
    assign _5874 = _5869 - _5269;
    assign _5875 = _5871 ? _5874 : _5869;
    assign _5876 = _5875[62:0];
    assign _5878 = { _5876,
                     _5877 };
    assign _5879 = _5878 < _5269;
    assign _5880 = ~ _5879;
    assign _5868 = _5849[61:61];
    assign _5865 = _5860 - _5269;
    assign _5866 = _5862 ? _5865 : _5860;
    assign _5867 = _5866[62:0];
    assign _5869 = { _5867,
                     _5868 };
    assign _5870 = _5869 < _5269;
    assign _5871 = ~ _5870;
    assign _5859 = _5849[62:62];
    assign _5856 = _5851 - _5269;
    assign _5857 = _5853 ? _5856 : _5851;
    assign _5858 = _5857[62:0];
    assign _5860 = { _5858,
                     _5859 };
    assign _5861 = _5860 < _5269;
    assign _5862 = ~ _5861;
    assign _5849 = _5261 - _5843;
    assign _5850 = _5849[63:63];
    assign _5851 = { _22185,
                     _5850 };
    assign _5852 = _5851 < _5269;
    assign _5853 = ~ _5852;
    assign _5854 = { _22185,
                     _5853 };
    assign _5855 = _5854[62:0];
    assign _5863 = { _5855,
                     _5862 };
    assign _5864 = _5863[62:0];
    assign _5872 = { _5864,
                     _5871 };
    assign _5873 = _5872[62:0];
    assign _5881 = { _5873,
                     _5880 };
    assign _5882 = _5881[62:0];
    assign _5890 = { _5882,
                     _5889 };
    assign _5891 = _5890[62:0];
    assign _5899 = { _5891,
                     _5898 };
    assign _5900 = _5899[62:0];
    assign _5908 = { _5900,
                     _5907 };
    assign _5909 = _5908[62:0];
    assign _5917 = { _5909,
                     _5916 };
    assign _5918 = _5917[62:0];
    assign _5926 = { _5918,
                     _5925 };
    assign _5927 = _5926[62:0];
    assign _5935 = { _5927,
                     _5934 };
    assign _5936 = _5935[62:0];
    assign _5944 = { _5936,
                     _5943 };
    assign _5945 = _5944[62:0];
    assign _5953 = { _5945,
                     _5952 };
    assign _5954 = _5953[62:0];
    assign _5962 = { _5954,
                     _5961 };
    assign _5963 = _5962[62:0];
    assign _5971 = { _5963,
                     _5970 };
    assign _5972 = _5971[62:0];
    assign _5980 = { _5972,
                     _5979 };
    assign _5981 = _5980[62:0];
    assign _5989 = { _5981,
                     _5988 };
    assign _5990 = _5989[62:0];
    assign _5998 = { _5990,
                     _5997 };
    assign _5999 = _5998[62:0];
    assign _6007 = { _5999,
                     _6006 };
    assign _6008 = _6007[62:0];
    assign _6016 = { _6008,
                     _6015 };
    assign _6017 = _6016[62:0];
    assign _6025 = { _6017,
                     _6024 };
    assign _6026 = _6025[62:0];
    assign _6034 = { _6026,
                     _6033 };
    assign _6035 = _6034[62:0];
    assign _6043 = { _6035,
                     _6042 };
    assign _6044 = _6043[62:0];
    assign _6052 = { _6044,
                     _6051 };
    assign _6053 = _6052[62:0];
    assign _6061 = { _6053,
                     _6060 };
    assign _6062 = _6061[62:0];
    assign _6070 = { _6062,
                     _6069 };
    assign _6071 = _6070[62:0];
    assign _6079 = { _6071,
                     _6078 };
    assign _6080 = _6079[62:0];
    assign _6088 = { _6080,
                     _6087 };
    assign _6089 = _6088[62:0];
    assign _6097 = { _6089,
                     _6096 };
    assign _6098 = _6097[62:0];
    assign _6106 = { _6098,
                     _6105 };
    assign _6107 = _6106[62:0];
    assign _6115 = { _6107,
                     _6114 };
    assign _6116 = _6115[62:0];
    assign _6124 = { _6116,
                     _6123 };
    assign _6125 = _6124[62:0];
    assign _6133 = { _6125,
                     _6132 };
    assign _6134 = _6133[62:0];
    assign _6142 = { _6134,
                     _6141 };
    assign _6143 = _6142[62:0];
    assign _6151 = { _6143,
                     _6150 };
    assign _6152 = _6151[62:0];
    assign _6160 = { _6152,
                     _6159 };
    assign _6161 = _6160[62:0];
    assign _6169 = { _6161,
                     _6168 };
    assign _6170 = _6169[62:0];
    assign _6178 = { _6170,
                     _6177 };
    assign _6179 = _6178[62:0];
    assign _6187 = { _6179,
                     _6186 };
    assign _6188 = _6187[62:0];
    assign _6196 = { _6188,
                     _6195 };
    assign _6197 = _6196[62:0];
    assign _6205 = { _6197,
                     _6204 };
    assign _6206 = _6205[62:0];
    assign _6214 = { _6206,
                     _6213 };
    assign _6215 = _6214[62:0];
    assign _6223 = { _6215,
                     _6222 };
    assign _6224 = _6223[62:0];
    assign _6232 = { _6224,
                     _6231 };
    assign _6233 = _6232[62:0];
    assign _6241 = { _6233,
                     _6240 };
    assign _6242 = _6241[62:0];
    assign _6250 = { _6242,
                     _6249 };
    assign _6251 = _6250[62:0];
    assign _6259 = { _6251,
                     _6258 };
    assign _6260 = _6259[62:0];
    assign _6268 = { _6260,
                     _6267 };
    assign _6269 = _6268[62:0];
    assign _6277 = { _6269,
                     _6276 };
    assign _6278 = _6277[62:0];
    assign _6286 = { _6278,
                     _6285 };
    assign _6287 = _6286[62:0];
    assign _6295 = { _6287,
                     _6294 };
    assign _6296 = _6295[62:0];
    assign _6304 = { _6296,
                     _6303 };
    assign _6305 = _6304[62:0];
    assign _6313 = { _6305,
                     _6312 };
    assign _6314 = _6313[62:0];
    assign _6322 = { _6314,
                     _6321 };
    assign _6323 = _6322[62:0];
    assign _6331 = { _6323,
                     _6330 };
    assign _6332 = _6331[62:0];
    assign _6340 = { _6332,
                     _6339 };
    assign _6341 = _6340[62:0];
    assign _6349 = { _6341,
                     _6348 };
    assign _6350 = _6349[62:0];
    assign _6358 = { _6350,
                     _6357 };
    assign _6359 = _6358[62:0];
    assign _6367 = { _6359,
                     _6366 };
    assign _6368 = _6367[62:0];
    assign _6376 = { _6368,
                     _6375 };
    assign _6377 = _6376[62:0];
    assign _6385 = { _6377,
                     _6384 };
    assign _6386 = _6385[62:0];
    assign _6394 = { _6386,
                     _6393 };
    assign _6395 = _6394[62:0];
    assign _6403 = { _6395,
                     _6402 };
    assign _6404 = _6403[62:0];
    assign _6412 = { _6404,
                     _6411 };
    assign _6413 = _6412[62:0];
    assign _6421 = { _6413,
                     _6420 };
    assign _6423 = _6421 + _22186;
    assign _6424 = _6423 * _5843;
    assign _6425 = _6424[63:0];
    assign _7007 = _6425 + _7006;
    assign _5835 = _5266[0:0];
    assign _5832 = _5827 - _5269;
    assign _5833 = _5829 ? _5832 : _5827;
    assign _5834 = _5833[62:0];
    assign _5836 = { _5834,
                     _5835 };
    assign _5837 = _5836 < _5269;
    assign _5838 = ~ _5837;
    assign _5826 = _5266[1:1];
    assign _5823 = _5818 - _5269;
    assign _5824 = _5820 ? _5823 : _5818;
    assign _5825 = _5824[62:0];
    assign _5827 = { _5825,
                     _5826 };
    assign _5828 = _5827 < _5269;
    assign _5829 = ~ _5828;
    assign _5817 = _5266[2:2];
    assign _5814 = _5809 - _5269;
    assign _5815 = _5811 ? _5814 : _5809;
    assign _5816 = _5815[62:0];
    assign _5818 = { _5816,
                     _5817 };
    assign _5819 = _5818 < _5269;
    assign _5820 = ~ _5819;
    assign _5808 = _5266[3:3];
    assign _5805 = _5800 - _5269;
    assign _5806 = _5802 ? _5805 : _5800;
    assign _5807 = _5806[62:0];
    assign _5809 = { _5807,
                     _5808 };
    assign _5810 = _5809 < _5269;
    assign _5811 = ~ _5810;
    assign _5799 = _5266[4:4];
    assign _5796 = _5791 - _5269;
    assign _5797 = _5793 ? _5796 : _5791;
    assign _5798 = _5797[62:0];
    assign _5800 = { _5798,
                     _5799 };
    assign _5801 = _5800 < _5269;
    assign _5802 = ~ _5801;
    assign _5790 = _5266[5:5];
    assign _5787 = _5782 - _5269;
    assign _5788 = _5784 ? _5787 : _5782;
    assign _5789 = _5788[62:0];
    assign _5791 = { _5789,
                     _5790 };
    assign _5792 = _5791 < _5269;
    assign _5793 = ~ _5792;
    assign _5781 = _5266[6:6];
    assign _5778 = _5773 - _5269;
    assign _5779 = _5775 ? _5778 : _5773;
    assign _5780 = _5779[62:0];
    assign _5782 = { _5780,
                     _5781 };
    assign _5783 = _5782 < _5269;
    assign _5784 = ~ _5783;
    assign _5772 = _5266[7:7];
    assign _5769 = _5764 - _5269;
    assign _5770 = _5766 ? _5769 : _5764;
    assign _5771 = _5770[62:0];
    assign _5773 = { _5771,
                     _5772 };
    assign _5774 = _5773 < _5269;
    assign _5775 = ~ _5774;
    assign _5763 = _5266[8:8];
    assign _5760 = _5755 - _5269;
    assign _5761 = _5757 ? _5760 : _5755;
    assign _5762 = _5761[62:0];
    assign _5764 = { _5762,
                     _5763 };
    assign _5765 = _5764 < _5269;
    assign _5766 = ~ _5765;
    assign _5754 = _5266[9:9];
    assign _5751 = _5746 - _5269;
    assign _5752 = _5748 ? _5751 : _5746;
    assign _5753 = _5752[62:0];
    assign _5755 = { _5753,
                     _5754 };
    assign _5756 = _5755 < _5269;
    assign _5757 = ~ _5756;
    assign _5745 = _5266[10:10];
    assign _5742 = _5737 - _5269;
    assign _5743 = _5739 ? _5742 : _5737;
    assign _5744 = _5743[62:0];
    assign _5746 = { _5744,
                     _5745 };
    assign _5747 = _5746 < _5269;
    assign _5748 = ~ _5747;
    assign _5736 = _5266[11:11];
    assign _5733 = _5728 - _5269;
    assign _5734 = _5730 ? _5733 : _5728;
    assign _5735 = _5734[62:0];
    assign _5737 = { _5735,
                     _5736 };
    assign _5738 = _5737 < _5269;
    assign _5739 = ~ _5738;
    assign _5727 = _5266[12:12];
    assign _5724 = _5719 - _5269;
    assign _5725 = _5721 ? _5724 : _5719;
    assign _5726 = _5725[62:0];
    assign _5728 = { _5726,
                     _5727 };
    assign _5729 = _5728 < _5269;
    assign _5730 = ~ _5729;
    assign _5718 = _5266[13:13];
    assign _5715 = _5710 - _5269;
    assign _5716 = _5712 ? _5715 : _5710;
    assign _5717 = _5716[62:0];
    assign _5719 = { _5717,
                     _5718 };
    assign _5720 = _5719 < _5269;
    assign _5721 = ~ _5720;
    assign _5709 = _5266[14:14];
    assign _5706 = _5701 - _5269;
    assign _5707 = _5703 ? _5706 : _5701;
    assign _5708 = _5707[62:0];
    assign _5710 = { _5708,
                     _5709 };
    assign _5711 = _5710 < _5269;
    assign _5712 = ~ _5711;
    assign _5700 = _5266[15:15];
    assign _5697 = _5692 - _5269;
    assign _5698 = _5694 ? _5697 : _5692;
    assign _5699 = _5698[62:0];
    assign _5701 = { _5699,
                     _5700 };
    assign _5702 = _5701 < _5269;
    assign _5703 = ~ _5702;
    assign _5691 = _5266[16:16];
    assign _5688 = _5683 - _5269;
    assign _5689 = _5685 ? _5688 : _5683;
    assign _5690 = _5689[62:0];
    assign _5692 = { _5690,
                     _5691 };
    assign _5693 = _5692 < _5269;
    assign _5694 = ~ _5693;
    assign _5682 = _5266[17:17];
    assign _5679 = _5674 - _5269;
    assign _5680 = _5676 ? _5679 : _5674;
    assign _5681 = _5680[62:0];
    assign _5683 = { _5681,
                     _5682 };
    assign _5684 = _5683 < _5269;
    assign _5685 = ~ _5684;
    assign _5673 = _5266[18:18];
    assign _5670 = _5665 - _5269;
    assign _5671 = _5667 ? _5670 : _5665;
    assign _5672 = _5671[62:0];
    assign _5674 = { _5672,
                     _5673 };
    assign _5675 = _5674 < _5269;
    assign _5676 = ~ _5675;
    assign _5664 = _5266[19:19];
    assign _5661 = _5656 - _5269;
    assign _5662 = _5658 ? _5661 : _5656;
    assign _5663 = _5662[62:0];
    assign _5665 = { _5663,
                     _5664 };
    assign _5666 = _5665 < _5269;
    assign _5667 = ~ _5666;
    assign _5655 = _5266[20:20];
    assign _5652 = _5647 - _5269;
    assign _5653 = _5649 ? _5652 : _5647;
    assign _5654 = _5653[62:0];
    assign _5656 = { _5654,
                     _5655 };
    assign _5657 = _5656 < _5269;
    assign _5658 = ~ _5657;
    assign _5646 = _5266[21:21];
    assign _5643 = _5638 - _5269;
    assign _5644 = _5640 ? _5643 : _5638;
    assign _5645 = _5644[62:0];
    assign _5647 = { _5645,
                     _5646 };
    assign _5648 = _5647 < _5269;
    assign _5649 = ~ _5648;
    assign _5637 = _5266[22:22];
    assign _5634 = _5629 - _5269;
    assign _5635 = _5631 ? _5634 : _5629;
    assign _5636 = _5635[62:0];
    assign _5638 = { _5636,
                     _5637 };
    assign _5639 = _5638 < _5269;
    assign _5640 = ~ _5639;
    assign _5628 = _5266[23:23];
    assign _5625 = _5620 - _5269;
    assign _5626 = _5622 ? _5625 : _5620;
    assign _5627 = _5626[62:0];
    assign _5629 = { _5627,
                     _5628 };
    assign _5630 = _5629 < _5269;
    assign _5631 = ~ _5630;
    assign _5619 = _5266[24:24];
    assign _5616 = _5611 - _5269;
    assign _5617 = _5613 ? _5616 : _5611;
    assign _5618 = _5617[62:0];
    assign _5620 = { _5618,
                     _5619 };
    assign _5621 = _5620 < _5269;
    assign _5622 = ~ _5621;
    assign _5610 = _5266[25:25];
    assign _5607 = _5602 - _5269;
    assign _5608 = _5604 ? _5607 : _5602;
    assign _5609 = _5608[62:0];
    assign _5611 = { _5609,
                     _5610 };
    assign _5612 = _5611 < _5269;
    assign _5613 = ~ _5612;
    assign _5601 = _5266[26:26];
    assign _5598 = _5593 - _5269;
    assign _5599 = _5595 ? _5598 : _5593;
    assign _5600 = _5599[62:0];
    assign _5602 = { _5600,
                     _5601 };
    assign _5603 = _5602 < _5269;
    assign _5604 = ~ _5603;
    assign _5592 = _5266[27:27];
    assign _5589 = _5584 - _5269;
    assign _5590 = _5586 ? _5589 : _5584;
    assign _5591 = _5590[62:0];
    assign _5593 = { _5591,
                     _5592 };
    assign _5594 = _5593 < _5269;
    assign _5595 = ~ _5594;
    assign _5583 = _5266[28:28];
    assign _5580 = _5575 - _5269;
    assign _5581 = _5577 ? _5580 : _5575;
    assign _5582 = _5581[62:0];
    assign _5584 = { _5582,
                     _5583 };
    assign _5585 = _5584 < _5269;
    assign _5586 = ~ _5585;
    assign _5574 = _5266[29:29];
    assign _5571 = _5566 - _5269;
    assign _5572 = _5568 ? _5571 : _5566;
    assign _5573 = _5572[62:0];
    assign _5575 = { _5573,
                     _5574 };
    assign _5576 = _5575 < _5269;
    assign _5577 = ~ _5576;
    assign _5565 = _5266[30:30];
    assign _5562 = _5557 - _5269;
    assign _5563 = _5559 ? _5562 : _5557;
    assign _5564 = _5563[62:0];
    assign _5566 = { _5564,
                     _5565 };
    assign _5567 = _5566 < _5269;
    assign _5568 = ~ _5567;
    assign _5556 = _5266[31:31];
    assign _5553 = _5548 - _5269;
    assign _5554 = _5550 ? _5553 : _5548;
    assign _5555 = _5554[62:0];
    assign _5557 = { _5555,
                     _5556 };
    assign _5558 = _5557 < _5269;
    assign _5559 = ~ _5558;
    assign _5547 = _5266[32:32];
    assign _5544 = _5539 - _5269;
    assign _5545 = _5541 ? _5544 : _5539;
    assign _5546 = _5545[62:0];
    assign _5548 = { _5546,
                     _5547 };
    assign _5549 = _5548 < _5269;
    assign _5550 = ~ _5549;
    assign _5538 = _5266[33:33];
    assign _5535 = _5530 - _5269;
    assign _5536 = _5532 ? _5535 : _5530;
    assign _5537 = _5536[62:0];
    assign _5539 = { _5537,
                     _5538 };
    assign _5540 = _5539 < _5269;
    assign _5541 = ~ _5540;
    assign _5529 = _5266[34:34];
    assign _5526 = _5521 - _5269;
    assign _5527 = _5523 ? _5526 : _5521;
    assign _5528 = _5527[62:0];
    assign _5530 = { _5528,
                     _5529 };
    assign _5531 = _5530 < _5269;
    assign _5532 = ~ _5531;
    assign _5520 = _5266[35:35];
    assign _5517 = _5512 - _5269;
    assign _5518 = _5514 ? _5517 : _5512;
    assign _5519 = _5518[62:0];
    assign _5521 = { _5519,
                     _5520 };
    assign _5522 = _5521 < _5269;
    assign _5523 = ~ _5522;
    assign _5511 = _5266[36:36];
    assign _5508 = _5503 - _5269;
    assign _5509 = _5505 ? _5508 : _5503;
    assign _5510 = _5509[62:0];
    assign _5512 = { _5510,
                     _5511 };
    assign _5513 = _5512 < _5269;
    assign _5514 = ~ _5513;
    assign _5502 = _5266[37:37];
    assign _5499 = _5494 - _5269;
    assign _5500 = _5496 ? _5499 : _5494;
    assign _5501 = _5500[62:0];
    assign _5503 = { _5501,
                     _5502 };
    assign _5504 = _5503 < _5269;
    assign _5505 = ~ _5504;
    assign _5493 = _5266[38:38];
    assign _5490 = _5485 - _5269;
    assign _5491 = _5487 ? _5490 : _5485;
    assign _5492 = _5491[62:0];
    assign _5494 = { _5492,
                     _5493 };
    assign _5495 = _5494 < _5269;
    assign _5496 = ~ _5495;
    assign _5484 = _5266[39:39];
    assign _5481 = _5476 - _5269;
    assign _5482 = _5478 ? _5481 : _5476;
    assign _5483 = _5482[62:0];
    assign _5485 = { _5483,
                     _5484 };
    assign _5486 = _5485 < _5269;
    assign _5487 = ~ _5486;
    assign _5475 = _5266[40:40];
    assign _5472 = _5467 - _5269;
    assign _5473 = _5469 ? _5472 : _5467;
    assign _5474 = _5473[62:0];
    assign _5476 = { _5474,
                     _5475 };
    assign _5477 = _5476 < _5269;
    assign _5478 = ~ _5477;
    assign _5466 = _5266[41:41];
    assign _5463 = _5458 - _5269;
    assign _5464 = _5460 ? _5463 : _5458;
    assign _5465 = _5464[62:0];
    assign _5467 = { _5465,
                     _5466 };
    assign _5468 = _5467 < _5269;
    assign _5469 = ~ _5468;
    assign _5457 = _5266[42:42];
    assign _5454 = _5449 - _5269;
    assign _5455 = _5451 ? _5454 : _5449;
    assign _5456 = _5455[62:0];
    assign _5458 = { _5456,
                     _5457 };
    assign _5459 = _5458 < _5269;
    assign _5460 = ~ _5459;
    assign _5448 = _5266[43:43];
    assign _5445 = _5440 - _5269;
    assign _5446 = _5442 ? _5445 : _5440;
    assign _5447 = _5446[62:0];
    assign _5449 = { _5447,
                     _5448 };
    assign _5450 = _5449 < _5269;
    assign _5451 = ~ _5450;
    assign _5439 = _5266[44:44];
    assign _5436 = _5431 - _5269;
    assign _5437 = _5433 ? _5436 : _5431;
    assign _5438 = _5437[62:0];
    assign _5440 = { _5438,
                     _5439 };
    assign _5441 = _5440 < _5269;
    assign _5442 = ~ _5441;
    assign _5430 = _5266[45:45];
    assign _5427 = _5422 - _5269;
    assign _5428 = _5424 ? _5427 : _5422;
    assign _5429 = _5428[62:0];
    assign _5431 = { _5429,
                     _5430 };
    assign _5432 = _5431 < _5269;
    assign _5433 = ~ _5432;
    assign _5421 = _5266[46:46];
    assign _5418 = _5413 - _5269;
    assign _5419 = _5415 ? _5418 : _5413;
    assign _5420 = _5419[62:0];
    assign _5422 = { _5420,
                     _5421 };
    assign _5423 = _5422 < _5269;
    assign _5424 = ~ _5423;
    assign _5412 = _5266[47:47];
    assign _5409 = _5404 - _5269;
    assign _5410 = _5406 ? _5409 : _5404;
    assign _5411 = _5410[62:0];
    assign _5413 = { _5411,
                     _5412 };
    assign _5414 = _5413 < _5269;
    assign _5415 = ~ _5414;
    assign _5403 = _5266[48:48];
    assign _5400 = _5395 - _5269;
    assign _5401 = _5397 ? _5400 : _5395;
    assign _5402 = _5401[62:0];
    assign _5404 = { _5402,
                     _5403 };
    assign _5405 = _5404 < _5269;
    assign _5406 = ~ _5405;
    assign _5394 = _5266[49:49];
    assign _5391 = _5386 - _5269;
    assign _5392 = _5388 ? _5391 : _5386;
    assign _5393 = _5392[62:0];
    assign _5395 = { _5393,
                     _5394 };
    assign _5396 = _5395 < _5269;
    assign _5397 = ~ _5396;
    assign _5385 = _5266[50:50];
    assign _5382 = _5377 - _5269;
    assign _5383 = _5379 ? _5382 : _5377;
    assign _5384 = _5383[62:0];
    assign _5386 = { _5384,
                     _5385 };
    assign _5387 = _5386 < _5269;
    assign _5388 = ~ _5387;
    assign _5376 = _5266[51:51];
    assign _5373 = _5368 - _5269;
    assign _5374 = _5370 ? _5373 : _5368;
    assign _5375 = _5374[62:0];
    assign _5377 = { _5375,
                     _5376 };
    assign _5378 = _5377 < _5269;
    assign _5379 = ~ _5378;
    assign _5367 = _5266[52:52];
    assign _5364 = _5359 - _5269;
    assign _5365 = _5361 ? _5364 : _5359;
    assign _5366 = _5365[62:0];
    assign _5368 = { _5366,
                     _5367 };
    assign _5369 = _5368 < _5269;
    assign _5370 = ~ _5369;
    assign _5358 = _5266[53:53];
    assign _5355 = _5350 - _5269;
    assign _5356 = _5352 ? _5355 : _5350;
    assign _5357 = _5356[62:0];
    assign _5359 = { _5357,
                     _5358 };
    assign _5360 = _5359 < _5269;
    assign _5361 = ~ _5360;
    assign _5349 = _5266[54:54];
    assign _5346 = _5341 - _5269;
    assign _5347 = _5343 ? _5346 : _5341;
    assign _5348 = _5347[62:0];
    assign _5350 = { _5348,
                     _5349 };
    assign _5351 = _5350 < _5269;
    assign _5352 = ~ _5351;
    assign _5340 = _5266[55:55];
    assign _5337 = _5332 - _5269;
    assign _5338 = _5334 ? _5337 : _5332;
    assign _5339 = _5338[62:0];
    assign _5341 = { _5339,
                     _5340 };
    assign _5342 = _5341 < _5269;
    assign _5343 = ~ _5342;
    assign _5331 = _5266[56:56];
    assign _5328 = _5323 - _5269;
    assign _5329 = _5325 ? _5328 : _5323;
    assign _5330 = _5329[62:0];
    assign _5332 = { _5330,
                     _5331 };
    assign _5333 = _5332 < _5269;
    assign _5334 = ~ _5333;
    assign _5322 = _5266[57:57];
    assign _5319 = _5314 - _5269;
    assign _5320 = _5316 ? _5319 : _5314;
    assign _5321 = _5320[62:0];
    assign _5323 = { _5321,
                     _5322 };
    assign _5324 = _5323 < _5269;
    assign _5325 = ~ _5324;
    assign _5313 = _5266[58:58];
    assign _5310 = _5305 - _5269;
    assign _5311 = _5307 ? _5310 : _5305;
    assign _5312 = _5311[62:0];
    assign _5314 = { _5312,
                     _5313 };
    assign _5315 = _5314 < _5269;
    assign _5316 = ~ _5315;
    assign _5304 = _5266[59:59];
    assign _5301 = _5296 - _5269;
    assign _5302 = _5298 ? _5301 : _5296;
    assign _5303 = _5302[62:0];
    assign _5305 = { _5303,
                     _5304 };
    assign _5306 = _5305 < _5269;
    assign _5307 = ~ _5306;
    assign _5295 = _5266[60:60];
    assign _5292 = _5287 - _5269;
    assign _5293 = _5289 ? _5292 : _5287;
    assign _5294 = _5293[62:0];
    assign _5296 = { _5294,
                     _5295 };
    assign _5297 = _5296 < _5269;
    assign _5298 = ~ _5297;
    assign _5286 = _5266[61:61];
    assign _5283 = _5278 - _5269;
    assign _5284 = _5280 ? _5283 : _5278;
    assign _5285 = _5284[62:0];
    assign _5287 = { _5285,
                     _5286 };
    assign _5288 = _5287 < _5269;
    assign _5289 = ~ _5288;
    assign _5277 = _5266[62:62];
    assign _5274 = _5268 - _5269;
    assign _5275 = _5271 ? _5274 : _5268;
    assign _5276 = _5275[62:0];
    assign _5278 = { _5276,
                     _5277 };
    assign _5279 = _5278 < _5269;
    assign _5280 = ~ _5279;
    assign _5269 = 64'b0000000000000000000000000000000000000000000000000010011100010001;
    assign _5265 = 64'b0000000000000000000000000000000000000000000000000010011100010000;
    assign _5266 = _3 + _5265;
    assign _5267 = _5266[63:63];
    assign _5268 = { _22185,
                     _5267 };
    assign _5270 = _5268 < _5269;
    assign _5271 = ~ _5270;
    assign _5272 = { _22185,
                     _5271 };
    assign _5273 = _5272[62:0];
    assign _5281 = { _5273,
                     _5280 };
    assign _5282 = _5281[62:0];
    assign _5290 = { _5282,
                     _5289 };
    assign _5291 = _5290[62:0];
    assign _5299 = { _5291,
                     _5298 };
    assign _5300 = _5299[62:0];
    assign _5308 = { _5300,
                     _5307 };
    assign _5309 = _5308[62:0];
    assign _5317 = { _5309,
                     _5316 };
    assign _5318 = _5317[62:0];
    assign _5326 = { _5318,
                     _5325 };
    assign _5327 = _5326[62:0];
    assign _5335 = { _5327,
                     _5334 };
    assign _5336 = _5335[62:0];
    assign _5344 = { _5336,
                     _5343 };
    assign _5345 = _5344[62:0];
    assign _5353 = { _5345,
                     _5352 };
    assign _5354 = _5353[62:0];
    assign _5362 = { _5354,
                     _5361 };
    assign _5363 = _5362[62:0];
    assign _5371 = { _5363,
                     _5370 };
    assign _5372 = _5371[62:0];
    assign _5380 = { _5372,
                     _5379 };
    assign _5381 = _5380[62:0];
    assign _5389 = { _5381,
                     _5388 };
    assign _5390 = _5389[62:0];
    assign _5398 = { _5390,
                     _5397 };
    assign _5399 = _5398[62:0];
    assign _5407 = { _5399,
                     _5406 };
    assign _5408 = _5407[62:0];
    assign _5416 = { _5408,
                     _5415 };
    assign _5417 = _5416[62:0];
    assign _5425 = { _5417,
                     _5424 };
    assign _5426 = _5425[62:0];
    assign _5434 = { _5426,
                     _5433 };
    assign _5435 = _5434[62:0];
    assign _5443 = { _5435,
                     _5442 };
    assign _5444 = _5443[62:0];
    assign _5452 = { _5444,
                     _5451 };
    assign _5453 = _5452[62:0];
    assign _5461 = { _5453,
                     _5460 };
    assign _5462 = _5461[62:0];
    assign _5470 = { _5462,
                     _5469 };
    assign _5471 = _5470[62:0];
    assign _5479 = { _5471,
                     _5478 };
    assign _5480 = _5479[62:0];
    assign _5488 = { _5480,
                     _5487 };
    assign _5489 = _5488[62:0];
    assign _5497 = { _5489,
                     _5496 };
    assign _5498 = _5497[62:0];
    assign _5506 = { _5498,
                     _5505 };
    assign _5507 = _5506[62:0];
    assign _5515 = { _5507,
                     _5514 };
    assign _5516 = _5515[62:0];
    assign _5524 = { _5516,
                     _5523 };
    assign _5525 = _5524[62:0];
    assign _5533 = { _5525,
                     _5532 };
    assign _5534 = _5533[62:0];
    assign _5542 = { _5534,
                     _5541 };
    assign _5543 = _5542[62:0];
    assign _5551 = { _5543,
                     _5550 };
    assign _5552 = _5551[62:0];
    assign _5560 = { _5552,
                     _5559 };
    assign _5561 = _5560[62:0];
    assign _5569 = { _5561,
                     _5568 };
    assign _5570 = _5569[62:0];
    assign _5578 = { _5570,
                     _5577 };
    assign _5579 = _5578[62:0];
    assign _5587 = { _5579,
                     _5586 };
    assign _5588 = _5587[62:0];
    assign _5596 = { _5588,
                     _5595 };
    assign _5597 = _5596[62:0];
    assign _5605 = { _5597,
                     _5604 };
    assign _5606 = _5605[62:0];
    assign _5614 = { _5606,
                     _5613 };
    assign _5615 = _5614[62:0];
    assign _5623 = { _5615,
                     _5622 };
    assign _5624 = _5623[62:0];
    assign _5632 = { _5624,
                     _5631 };
    assign _5633 = _5632[62:0];
    assign _5641 = { _5633,
                     _5640 };
    assign _5642 = _5641[62:0];
    assign _5650 = { _5642,
                     _5649 };
    assign _5651 = _5650[62:0];
    assign _5659 = { _5651,
                     _5658 };
    assign _5660 = _5659[62:0];
    assign _5668 = { _5660,
                     _5667 };
    assign _5669 = _5668[62:0];
    assign _5677 = { _5669,
                     _5676 };
    assign _5678 = _5677[62:0];
    assign _5686 = { _5678,
                     _5685 };
    assign _5687 = _5686[62:0];
    assign _5695 = { _5687,
                     _5694 };
    assign _5696 = _5695[62:0];
    assign _5704 = { _5696,
                     _5703 };
    assign _5705 = _5704[62:0];
    assign _5713 = { _5705,
                     _5712 };
    assign _5714 = _5713[62:0];
    assign _5722 = { _5714,
                     _5721 };
    assign _5723 = _5722[62:0];
    assign _5731 = { _5723,
                     _5730 };
    assign _5732 = _5731[62:0];
    assign _5740 = { _5732,
                     _5739 };
    assign _5741 = _5740[62:0];
    assign _5749 = { _5741,
                     _5748 };
    assign _5750 = _5749[62:0];
    assign _5758 = { _5750,
                     _5757 };
    assign _5759 = _5758[62:0];
    assign _5767 = { _5759,
                     _5766 };
    assign _5768 = _5767[62:0];
    assign _5776 = { _5768,
                     _5775 };
    assign _5777 = _5776[62:0];
    assign _5785 = { _5777,
                     _5784 };
    assign _5786 = _5785[62:0];
    assign _5794 = { _5786,
                     _5793 };
    assign _5795 = _5794[62:0];
    assign _5803 = { _5795,
                     _5802 };
    assign _5804 = _5803[62:0];
    assign _5812 = { _5804,
                     _5811 };
    assign _5813 = _5812[62:0];
    assign _5821 = { _5813,
                     _5820 };
    assign _5822 = _5821[62:0];
    assign _5830 = { _5822,
                     _5829 };
    assign _5831 = _5830[62:0];
    assign _5839 = { _5831,
                     _5838 };
    assign _5840 = _5839 * _5269;
    assign _5841 = _5840[63:0];
    assign _5262 = 64'b0000000000000000000000000000000000000000100110001001101001101000;
    assign _5842 = _5262 < _5841;
    assign _5843 = _5842 ? _5841 : _5262;
    assign _5259 = 64'b0000000000000000000000000000000000000101111101011110000011111111;
    assign _5260 = _5 < _5259;
    assign _5261 = _5260 ? _5 : _5259;
    assign _5844 = _5261 < _5843;
    assign _5845 = ~ _5844;
    assign _7008 = _5845 ? _7007 : _21604;
    assign _5249 = _4680[0:0];
    assign _5246 = _5241 - _22192;
    assign _5247 = _5243 ? _5246 : _5241;
    assign _5248 = _5247[62:0];
    assign _5250 = { _5248,
                     _5249 };
    assign _5251 = _5250 < _22192;
    assign _5252 = ~ _5251;
    assign _5240 = _4680[1:1];
    assign _5237 = _5232 - _22192;
    assign _5238 = _5234 ? _5237 : _5232;
    assign _5239 = _5238[62:0];
    assign _5241 = { _5239,
                     _5240 };
    assign _5242 = _5241 < _22192;
    assign _5243 = ~ _5242;
    assign _5231 = _4680[2:2];
    assign _5228 = _5223 - _22192;
    assign _5229 = _5225 ? _5228 : _5223;
    assign _5230 = _5229[62:0];
    assign _5232 = { _5230,
                     _5231 };
    assign _5233 = _5232 < _22192;
    assign _5234 = ~ _5233;
    assign _5222 = _4680[3:3];
    assign _5219 = _5214 - _22192;
    assign _5220 = _5216 ? _5219 : _5214;
    assign _5221 = _5220[62:0];
    assign _5223 = { _5221,
                     _5222 };
    assign _5224 = _5223 < _22192;
    assign _5225 = ~ _5224;
    assign _5213 = _4680[4:4];
    assign _5210 = _5205 - _22192;
    assign _5211 = _5207 ? _5210 : _5205;
    assign _5212 = _5211[62:0];
    assign _5214 = { _5212,
                     _5213 };
    assign _5215 = _5214 < _22192;
    assign _5216 = ~ _5215;
    assign _5204 = _4680[5:5];
    assign _5201 = _5196 - _22192;
    assign _5202 = _5198 ? _5201 : _5196;
    assign _5203 = _5202[62:0];
    assign _5205 = { _5203,
                     _5204 };
    assign _5206 = _5205 < _22192;
    assign _5207 = ~ _5206;
    assign _5195 = _4680[6:6];
    assign _5192 = _5187 - _22192;
    assign _5193 = _5189 ? _5192 : _5187;
    assign _5194 = _5193[62:0];
    assign _5196 = { _5194,
                     _5195 };
    assign _5197 = _5196 < _22192;
    assign _5198 = ~ _5197;
    assign _5186 = _4680[7:7];
    assign _5183 = _5178 - _22192;
    assign _5184 = _5180 ? _5183 : _5178;
    assign _5185 = _5184[62:0];
    assign _5187 = { _5185,
                     _5186 };
    assign _5188 = _5187 < _22192;
    assign _5189 = ~ _5188;
    assign _5177 = _4680[8:8];
    assign _5174 = _5169 - _22192;
    assign _5175 = _5171 ? _5174 : _5169;
    assign _5176 = _5175[62:0];
    assign _5178 = { _5176,
                     _5177 };
    assign _5179 = _5178 < _22192;
    assign _5180 = ~ _5179;
    assign _5168 = _4680[9:9];
    assign _5165 = _5160 - _22192;
    assign _5166 = _5162 ? _5165 : _5160;
    assign _5167 = _5166[62:0];
    assign _5169 = { _5167,
                     _5168 };
    assign _5170 = _5169 < _22192;
    assign _5171 = ~ _5170;
    assign _5159 = _4680[10:10];
    assign _5156 = _5151 - _22192;
    assign _5157 = _5153 ? _5156 : _5151;
    assign _5158 = _5157[62:0];
    assign _5160 = { _5158,
                     _5159 };
    assign _5161 = _5160 < _22192;
    assign _5162 = ~ _5161;
    assign _5150 = _4680[11:11];
    assign _5147 = _5142 - _22192;
    assign _5148 = _5144 ? _5147 : _5142;
    assign _5149 = _5148[62:0];
    assign _5151 = { _5149,
                     _5150 };
    assign _5152 = _5151 < _22192;
    assign _5153 = ~ _5152;
    assign _5141 = _4680[12:12];
    assign _5138 = _5133 - _22192;
    assign _5139 = _5135 ? _5138 : _5133;
    assign _5140 = _5139[62:0];
    assign _5142 = { _5140,
                     _5141 };
    assign _5143 = _5142 < _22192;
    assign _5144 = ~ _5143;
    assign _5132 = _4680[13:13];
    assign _5129 = _5124 - _22192;
    assign _5130 = _5126 ? _5129 : _5124;
    assign _5131 = _5130[62:0];
    assign _5133 = { _5131,
                     _5132 };
    assign _5134 = _5133 < _22192;
    assign _5135 = ~ _5134;
    assign _5123 = _4680[14:14];
    assign _5120 = _5115 - _22192;
    assign _5121 = _5117 ? _5120 : _5115;
    assign _5122 = _5121[62:0];
    assign _5124 = { _5122,
                     _5123 };
    assign _5125 = _5124 < _22192;
    assign _5126 = ~ _5125;
    assign _5114 = _4680[15:15];
    assign _5111 = _5106 - _22192;
    assign _5112 = _5108 ? _5111 : _5106;
    assign _5113 = _5112[62:0];
    assign _5115 = { _5113,
                     _5114 };
    assign _5116 = _5115 < _22192;
    assign _5117 = ~ _5116;
    assign _5105 = _4680[16:16];
    assign _5102 = _5097 - _22192;
    assign _5103 = _5099 ? _5102 : _5097;
    assign _5104 = _5103[62:0];
    assign _5106 = { _5104,
                     _5105 };
    assign _5107 = _5106 < _22192;
    assign _5108 = ~ _5107;
    assign _5096 = _4680[17:17];
    assign _5093 = _5088 - _22192;
    assign _5094 = _5090 ? _5093 : _5088;
    assign _5095 = _5094[62:0];
    assign _5097 = { _5095,
                     _5096 };
    assign _5098 = _5097 < _22192;
    assign _5099 = ~ _5098;
    assign _5087 = _4680[18:18];
    assign _5084 = _5079 - _22192;
    assign _5085 = _5081 ? _5084 : _5079;
    assign _5086 = _5085[62:0];
    assign _5088 = { _5086,
                     _5087 };
    assign _5089 = _5088 < _22192;
    assign _5090 = ~ _5089;
    assign _5078 = _4680[19:19];
    assign _5075 = _5070 - _22192;
    assign _5076 = _5072 ? _5075 : _5070;
    assign _5077 = _5076[62:0];
    assign _5079 = { _5077,
                     _5078 };
    assign _5080 = _5079 < _22192;
    assign _5081 = ~ _5080;
    assign _5069 = _4680[20:20];
    assign _5066 = _5061 - _22192;
    assign _5067 = _5063 ? _5066 : _5061;
    assign _5068 = _5067[62:0];
    assign _5070 = { _5068,
                     _5069 };
    assign _5071 = _5070 < _22192;
    assign _5072 = ~ _5071;
    assign _5060 = _4680[21:21];
    assign _5057 = _5052 - _22192;
    assign _5058 = _5054 ? _5057 : _5052;
    assign _5059 = _5058[62:0];
    assign _5061 = { _5059,
                     _5060 };
    assign _5062 = _5061 < _22192;
    assign _5063 = ~ _5062;
    assign _5051 = _4680[22:22];
    assign _5048 = _5043 - _22192;
    assign _5049 = _5045 ? _5048 : _5043;
    assign _5050 = _5049[62:0];
    assign _5052 = { _5050,
                     _5051 };
    assign _5053 = _5052 < _22192;
    assign _5054 = ~ _5053;
    assign _5042 = _4680[23:23];
    assign _5039 = _5034 - _22192;
    assign _5040 = _5036 ? _5039 : _5034;
    assign _5041 = _5040[62:0];
    assign _5043 = { _5041,
                     _5042 };
    assign _5044 = _5043 < _22192;
    assign _5045 = ~ _5044;
    assign _5033 = _4680[24:24];
    assign _5030 = _5025 - _22192;
    assign _5031 = _5027 ? _5030 : _5025;
    assign _5032 = _5031[62:0];
    assign _5034 = { _5032,
                     _5033 };
    assign _5035 = _5034 < _22192;
    assign _5036 = ~ _5035;
    assign _5024 = _4680[25:25];
    assign _5021 = _5016 - _22192;
    assign _5022 = _5018 ? _5021 : _5016;
    assign _5023 = _5022[62:0];
    assign _5025 = { _5023,
                     _5024 };
    assign _5026 = _5025 < _22192;
    assign _5027 = ~ _5026;
    assign _5015 = _4680[26:26];
    assign _5012 = _5007 - _22192;
    assign _5013 = _5009 ? _5012 : _5007;
    assign _5014 = _5013[62:0];
    assign _5016 = { _5014,
                     _5015 };
    assign _5017 = _5016 < _22192;
    assign _5018 = ~ _5017;
    assign _5006 = _4680[27:27];
    assign _5003 = _4998 - _22192;
    assign _5004 = _5000 ? _5003 : _4998;
    assign _5005 = _5004[62:0];
    assign _5007 = { _5005,
                     _5006 };
    assign _5008 = _5007 < _22192;
    assign _5009 = ~ _5008;
    assign _4997 = _4680[28:28];
    assign _4994 = _4989 - _22192;
    assign _4995 = _4991 ? _4994 : _4989;
    assign _4996 = _4995[62:0];
    assign _4998 = { _4996,
                     _4997 };
    assign _4999 = _4998 < _22192;
    assign _5000 = ~ _4999;
    assign _4988 = _4680[29:29];
    assign _4985 = _4980 - _22192;
    assign _4986 = _4982 ? _4985 : _4980;
    assign _4987 = _4986[62:0];
    assign _4989 = { _4987,
                     _4988 };
    assign _4990 = _4989 < _22192;
    assign _4991 = ~ _4990;
    assign _4979 = _4680[30:30];
    assign _4976 = _4971 - _22192;
    assign _4977 = _4973 ? _4976 : _4971;
    assign _4978 = _4977[62:0];
    assign _4980 = { _4978,
                     _4979 };
    assign _4981 = _4980 < _22192;
    assign _4982 = ~ _4981;
    assign _4970 = _4680[31:31];
    assign _4967 = _4962 - _22192;
    assign _4968 = _4964 ? _4967 : _4962;
    assign _4969 = _4968[62:0];
    assign _4971 = { _4969,
                     _4970 };
    assign _4972 = _4971 < _22192;
    assign _4973 = ~ _4972;
    assign _4961 = _4680[32:32];
    assign _4958 = _4953 - _22192;
    assign _4959 = _4955 ? _4958 : _4953;
    assign _4960 = _4959[62:0];
    assign _4962 = { _4960,
                     _4961 };
    assign _4963 = _4962 < _22192;
    assign _4964 = ~ _4963;
    assign _4952 = _4680[33:33];
    assign _4949 = _4944 - _22192;
    assign _4950 = _4946 ? _4949 : _4944;
    assign _4951 = _4950[62:0];
    assign _4953 = { _4951,
                     _4952 };
    assign _4954 = _4953 < _22192;
    assign _4955 = ~ _4954;
    assign _4943 = _4680[34:34];
    assign _4940 = _4935 - _22192;
    assign _4941 = _4937 ? _4940 : _4935;
    assign _4942 = _4941[62:0];
    assign _4944 = { _4942,
                     _4943 };
    assign _4945 = _4944 < _22192;
    assign _4946 = ~ _4945;
    assign _4934 = _4680[35:35];
    assign _4931 = _4926 - _22192;
    assign _4932 = _4928 ? _4931 : _4926;
    assign _4933 = _4932[62:0];
    assign _4935 = { _4933,
                     _4934 };
    assign _4936 = _4935 < _22192;
    assign _4937 = ~ _4936;
    assign _4925 = _4680[36:36];
    assign _4922 = _4917 - _22192;
    assign _4923 = _4919 ? _4922 : _4917;
    assign _4924 = _4923[62:0];
    assign _4926 = { _4924,
                     _4925 };
    assign _4927 = _4926 < _22192;
    assign _4928 = ~ _4927;
    assign _4916 = _4680[37:37];
    assign _4913 = _4908 - _22192;
    assign _4914 = _4910 ? _4913 : _4908;
    assign _4915 = _4914[62:0];
    assign _4917 = { _4915,
                     _4916 };
    assign _4918 = _4917 < _22192;
    assign _4919 = ~ _4918;
    assign _4907 = _4680[38:38];
    assign _4904 = _4899 - _22192;
    assign _4905 = _4901 ? _4904 : _4899;
    assign _4906 = _4905[62:0];
    assign _4908 = { _4906,
                     _4907 };
    assign _4909 = _4908 < _22192;
    assign _4910 = ~ _4909;
    assign _4898 = _4680[39:39];
    assign _4895 = _4890 - _22192;
    assign _4896 = _4892 ? _4895 : _4890;
    assign _4897 = _4896[62:0];
    assign _4899 = { _4897,
                     _4898 };
    assign _4900 = _4899 < _22192;
    assign _4901 = ~ _4900;
    assign _4889 = _4680[40:40];
    assign _4886 = _4881 - _22192;
    assign _4887 = _4883 ? _4886 : _4881;
    assign _4888 = _4887[62:0];
    assign _4890 = { _4888,
                     _4889 };
    assign _4891 = _4890 < _22192;
    assign _4892 = ~ _4891;
    assign _4880 = _4680[41:41];
    assign _4877 = _4872 - _22192;
    assign _4878 = _4874 ? _4877 : _4872;
    assign _4879 = _4878[62:0];
    assign _4881 = { _4879,
                     _4880 };
    assign _4882 = _4881 < _22192;
    assign _4883 = ~ _4882;
    assign _4871 = _4680[42:42];
    assign _4868 = _4863 - _22192;
    assign _4869 = _4865 ? _4868 : _4863;
    assign _4870 = _4869[62:0];
    assign _4872 = { _4870,
                     _4871 };
    assign _4873 = _4872 < _22192;
    assign _4874 = ~ _4873;
    assign _4862 = _4680[43:43];
    assign _4859 = _4854 - _22192;
    assign _4860 = _4856 ? _4859 : _4854;
    assign _4861 = _4860[62:0];
    assign _4863 = { _4861,
                     _4862 };
    assign _4864 = _4863 < _22192;
    assign _4865 = ~ _4864;
    assign _4853 = _4680[44:44];
    assign _4850 = _4845 - _22192;
    assign _4851 = _4847 ? _4850 : _4845;
    assign _4852 = _4851[62:0];
    assign _4854 = { _4852,
                     _4853 };
    assign _4855 = _4854 < _22192;
    assign _4856 = ~ _4855;
    assign _4844 = _4680[45:45];
    assign _4841 = _4836 - _22192;
    assign _4842 = _4838 ? _4841 : _4836;
    assign _4843 = _4842[62:0];
    assign _4845 = { _4843,
                     _4844 };
    assign _4846 = _4845 < _22192;
    assign _4847 = ~ _4846;
    assign _4835 = _4680[46:46];
    assign _4832 = _4827 - _22192;
    assign _4833 = _4829 ? _4832 : _4827;
    assign _4834 = _4833[62:0];
    assign _4836 = { _4834,
                     _4835 };
    assign _4837 = _4836 < _22192;
    assign _4838 = ~ _4837;
    assign _4826 = _4680[47:47];
    assign _4823 = _4818 - _22192;
    assign _4824 = _4820 ? _4823 : _4818;
    assign _4825 = _4824[62:0];
    assign _4827 = { _4825,
                     _4826 };
    assign _4828 = _4827 < _22192;
    assign _4829 = ~ _4828;
    assign _4817 = _4680[48:48];
    assign _4814 = _4809 - _22192;
    assign _4815 = _4811 ? _4814 : _4809;
    assign _4816 = _4815[62:0];
    assign _4818 = { _4816,
                     _4817 };
    assign _4819 = _4818 < _22192;
    assign _4820 = ~ _4819;
    assign _4808 = _4680[49:49];
    assign _4805 = _4800 - _22192;
    assign _4806 = _4802 ? _4805 : _4800;
    assign _4807 = _4806[62:0];
    assign _4809 = { _4807,
                     _4808 };
    assign _4810 = _4809 < _22192;
    assign _4811 = ~ _4810;
    assign _4799 = _4680[50:50];
    assign _4796 = _4791 - _22192;
    assign _4797 = _4793 ? _4796 : _4791;
    assign _4798 = _4797[62:0];
    assign _4800 = { _4798,
                     _4799 };
    assign _4801 = _4800 < _22192;
    assign _4802 = ~ _4801;
    assign _4790 = _4680[51:51];
    assign _4787 = _4782 - _22192;
    assign _4788 = _4784 ? _4787 : _4782;
    assign _4789 = _4788[62:0];
    assign _4791 = { _4789,
                     _4790 };
    assign _4792 = _4791 < _22192;
    assign _4793 = ~ _4792;
    assign _4781 = _4680[52:52];
    assign _4778 = _4773 - _22192;
    assign _4779 = _4775 ? _4778 : _4773;
    assign _4780 = _4779[62:0];
    assign _4782 = { _4780,
                     _4781 };
    assign _4783 = _4782 < _22192;
    assign _4784 = ~ _4783;
    assign _4772 = _4680[53:53];
    assign _4769 = _4764 - _22192;
    assign _4770 = _4766 ? _4769 : _4764;
    assign _4771 = _4770[62:0];
    assign _4773 = { _4771,
                     _4772 };
    assign _4774 = _4773 < _22192;
    assign _4775 = ~ _4774;
    assign _4763 = _4680[54:54];
    assign _4760 = _4755 - _22192;
    assign _4761 = _4757 ? _4760 : _4755;
    assign _4762 = _4761[62:0];
    assign _4764 = { _4762,
                     _4763 };
    assign _4765 = _4764 < _22192;
    assign _4766 = ~ _4765;
    assign _4754 = _4680[55:55];
    assign _4751 = _4746 - _22192;
    assign _4752 = _4748 ? _4751 : _4746;
    assign _4753 = _4752[62:0];
    assign _4755 = { _4753,
                     _4754 };
    assign _4756 = _4755 < _22192;
    assign _4757 = ~ _4756;
    assign _4745 = _4680[56:56];
    assign _4742 = _4737 - _22192;
    assign _4743 = _4739 ? _4742 : _4737;
    assign _4744 = _4743[62:0];
    assign _4746 = { _4744,
                     _4745 };
    assign _4747 = _4746 < _22192;
    assign _4748 = ~ _4747;
    assign _4736 = _4680[57:57];
    assign _4733 = _4728 - _22192;
    assign _4734 = _4730 ? _4733 : _4728;
    assign _4735 = _4734[62:0];
    assign _4737 = { _4735,
                     _4736 };
    assign _4738 = _4737 < _22192;
    assign _4739 = ~ _4738;
    assign _4727 = _4680[58:58];
    assign _4724 = _4719 - _22192;
    assign _4725 = _4721 ? _4724 : _4719;
    assign _4726 = _4725[62:0];
    assign _4728 = { _4726,
                     _4727 };
    assign _4729 = _4728 < _22192;
    assign _4730 = ~ _4729;
    assign _4718 = _4680[59:59];
    assign _4715 = _4710 - _22192;
    assign _4716 = _4712 ? _4715 : _4710;
    assign _4717 = _4716[62:0];
    assign _4719 = { _4717,
                     _4718 };
    assign _4720 = _4719 < _22192;
    assign _4721 = ~ _4720;
    assign _4709 = _4680[60:60];
    assign _4706 = _4701 - _22192;
    assign _4707 = _4703 ? _4706 : _4701;
    assign _4708 = _4707[62:0];
    assign _4710 = { _4708,
                     _4709 };
    assign _4711 = _4710 < _22192;
    assign _4712 = ~ _4711;
    assign _4700 = _4680[61:61];
    assign _4697 = _4692 - _22192;
    assign _4698 = _4694 ? _4697 : _4692;
    assign _4699 = _4698[62:0];
    assign _4701 = { _4699,
                     _4700 };
    assign _4702 = _4701 < _22192;
    assign _4703 = ~ _4702;
    assign _4691 = _4680[62:62];
    assign _4688 = _4682 - _22192;
    assign _4689 = _4685 ? _4688 : _4682;
    assign _4690 = _4689[62:0];
    assign _4692 = { _4690,
                     _4691 };
    assign _4693 = _4692 < _22192;
    assign _4694 = ~ _4693;
    assign _4678 = _4670 + _22186;
    assign _4679 = _4670 * _4678;
    assign _4680 = _4679[63:0];
    assign _4681 = _4680[63:63];
    assign _4682 = { _22185,
                     _4681 };
    assign _4684 = _4682 < _22192;
    assign _4685 = ~ _4684;
    assign _4686 = { _22185,
                     _4685 };
    assign _4687 = _4686[62:0];
    assign _4695 = { _4687,
                     _4694 };
    assign _4696 = _4695[62:0];
    assign _4704 = { _4696,
                     _4703 };
    assign _4705 = _4704[62:0];
    assign _4713 = { _4705,
                     _4712 };
    assign _4714 = _4713[62:0];
    assign _4722 = { _4714,
                     _4721 };
    assign _4723 = _4722[62:0];
    assign _4731 = { _4723,
                     _4730 };
    assign _4732 = _4731[62:0];
    assign _4740 = { _4732,
                     _4739 };
    assign _4741 = _4740[62:0];
    assign _4749 = { _4741,
                     _4748 };
    assign _4750 = _4749[62:0];
    assign _4758 = { _4750,
                     _4757 };
    assign _4759 = _4758[62:0];
    assign _4767 = { _4759,
                     _4766 };
    assign _4768 = _4767[62:0];
    assign _4776 = { _4768,
                     _4775 };
    assign _4777 = _4776[62:0];
    assign _4785 = { _4777,
                     _4784 };
    assign _4786 = _4785[62:0];
    assign _4794 = { _4786,
                     _4793 };
    assign _4795 = _4794[62:0];
    assign _4803 = { _4795,
                     _4802 };
    assign _4804 = _4803[62:0];
    assign _4812 = { _4804,
                     _4811 };
    assign _4813 = _4812[62:0];
    assign _4821 = { _4813,
                     _4820 };
    assign _4822 = _4821[62:0];
    assign _4830 = { _4822,
                     _4829 };
    assign _4831 = _4830[62:0];
    assign _4839 = { _4831,
                     _4838 };
    assign _4840 = _4839[62:0];
    assign _4848 = { _4840,
                     _4847 };
    assign _4849 = _4848[62:0];
    assign _4857 = { _4849,
                     _4856 };
    assign _4858 = _4857[62:0];
    assign _4866 = { _4858,
                     _4865 };
    assign _4867 = _4866[62:0];
    assign _4875 = { _4867,
                     _4874 };
    assign _4876 = _4875[62:0];
    assign _4884 = { _4876,
                     _4883 };
    assign _4885 = _4884[62:0];
    assign _4893 = { _4885,
                     _4892 };
    assign _4894 = _4893[62:0];
    assign _4902 = { _4894,
                     _4901 };
    assign _4903 = _4902[62:0];
    assign _4911 = { _4903,
                     _4910 };
    assign _4912 = _4911[62:0];
    assign _4920 = { _4912,
                     _4919 };
    assign _4921 = _4920[62:0];
    assign _4929 = { _4921,
                     _4928 };
    assign _4930 = _4929[62:0];
    assign _4938 = { _4930,
                     _4937 };
    assign _4939 = _4938[62:0];
    assign _4947 = { _4939,
                     _4946 };
    assign _4948 = _4947[62:0];
    assign _4956 = { _4948,
                     _4955 };
    assign _4957 = _4956[62:0];
    assign _4965 = { _4957,
                     _4964 };
    assign _4966 = _4965[62:0];
    assign _4974 = { _4966,
                     _4973 };
    assign _4975 = _4974[62:0];
    assign _4983 = { _4975,
                     _4982 };
    assign _4984 = _4983[62:0];
    assign _4992 = { _4984,
                     _4991 };
    assign _4993 = _4992[62:0];
    assign _5001 = { _4993,
                     _5000 };
    assign _5002 = _5001[62:0];
    assign _5010 = { _5002,
                     _5009 };
    assign _5011 = _5010[62:0];
    assign _5019 = { _5011,
                     _5018 };
    assign _5020 = _5019[62:0];
    assign _5028 = { _5020,
                     _5027 };
    assign _5029 = _5028[62:0];
    assign _5037 = { _5029,
                     _5036 };
    assign _5038 = _5037[62:0];
    assign _5046 = { _5038,
                     _5045 };
    assign _5047 = _5046[62:0];
    assign _5055 = { _5047,
                     _5054 };
    assign _5056 = _5055[62:0];
    assign _5064 = { _5056,
                     _5063 };
    assign _5065 = _5064[62:0];
    assign _5073 = { _5065,
                     _5072 };
    assign _5074 = _5073[62:0];
    assign _5082 = { _5074,
                     _5081 };
    assign _5083 = _5082[62:0];
    assign _5091 = { _5083,
                     _5090 };
    assign _5092 = _5091[62:0];
    assign _5100 = { _5092,
                     _5099 };
    assign _5101 = _5100[62:0];
    assign _5109 = { _5101,
                     _5108 };
    assign _5110 = _5109[62:0];
    assign _5118 = { _5110,
                     _5117 };
    assign _5119 = _5118[62:0];
    assign _5127 = { _5119,
                     _5126 };
    assign _5128 = _5127[62:0];
    assign _5136 = { _5128,
                     _5135 };
    assign _5137 = _5136[62:0];
    assign _5145 = { _5137,
                     _5144 };
    assign _5146 = _5145[62:0];
    assign _5154 = { _5146,
                     _5153 };
    assign _5155 = _5154[62:0];
    assign _5163 = { _5155,
                     _5162 };
    assign _5164 = _5163[62:0];
    assign _5172 = { _5164,
                     _5171 };
    assign _5173 = _5172[62:0];
    assign _5181 = { _5173,
                     _5180 };
    assign _5182 = _5181[62:0];
    assign _5190 = { _5182,
                     _5189 };
    assign _5191 = _5190[62:0];
    assign _5199 = { _5191,
                     _5198 };
    assign _5200 = _5199[62:0];
    assign _5208 = { _5200,
                     _5207 };
    assign _5209 = _5208[62:0];
    assign _5217 = { _5209,
                     _5216 };
    assign _5218 = _5217[62:0];
    assign _5226 = { _5218,
                     _5225 };
    assign _5227 = _5226[62:0];
    assign _5235 = { _5227,
                     _5234 };
    assign _5236 = _5235[62:0];
    assign _5244 = { _5236,
                     _5243 };
    assign _5245 = _5244[62:0];
    assign _5253 = { _5245,
                     _5252 };
    assign _5254 = _3518 * _5253;
    assign _5255 = _5254[63:0];
    assign _4666 = _4098[0:0];
    assign _4663 = _4658 - _3518;
    assign _4664 = _4660 ? _4663 : _4658;
    assign _4665 = _4664[62:0];
    assign _4667 = { _4665,
                     _4666 };
    assign _4668 = _4667 < _3518;
    assign _4669 = ~ _4668;
    assign _4657 = _4098[1:1];
    assign _4654 = _4649 - _3518;
    assign _4655 = _4651 ? _4654 : _4649;
    assign _4656 = _4655[62:0];
    assign _4658 = { _4656,
                     _4657 };
    assign _4659 = _4658 < _3518;
    assign _4660 = ~ _4659;
    assign _4648 = _4098[2:2];
    assign _4645 = _4640 - _3518;
    assign _4646 = _4642 ? _4645 : _4640;
    assign _4647 = _4646[62:0];
    assign _4649 = { _4647,
                     _4648 };
    assign _4650 = _4649 < _3518;
    assign _4651 = ~ _4650;
    assign _4639 = _4098[3:3];
    assign _4636 = _4631 - _3518;
    assign _4637 = _4633 ? _4636 : _4631;
    assign _4638 = _4637[62:0];
    assign _4640 = { _4638,
                     _4639 };
    assign _4641 = _4640 < _3518;
    assign _4642 = ~ _4641;
    assign _4630 = _4098[4:4];
    assign _4627 = _4622 - _3518;
    assign _4628 = _4624 ? _4627 : _4622;
    assign _4629 = _4628[62:0];
    assign _4631 = { _4629,
                     _4630 };
    assign _4632 = _4631 < _3518;
    assign _4633 = ~ _4632;
    assign _4621 = _4098[5:5];
    assign _4618 = _4613 - _3518;
    assign _4619 = _4615 ? _4618 : _4613;
    assign _4620 = _4619[62:0];
    assign _4622 = { _4620,
                     _4621 };
    assign _4623 = _4622 < _3518;
    assign _4624 = ~ _4623;
    assign _4612 = _4098[6:6];
    assign _4609 = _4604 - _3518;
    assign _4610 = _4606 ? _4609 : _4604;
    assign _4611 = _4610[62:0];
    assign _4613 = { _4611,
                     _4612 };
    assign _4614 = _4613 < _3518;
    assign _4615 = ~ _4614;
    assign _4603 = _4098[7:7];
    assign _4600 = _4595 - _3518;
    assign _4601 = _4597 ? _4600 : _4595;
    assign _4602 = _4601[62:0];
    assign _4604 = { _4602,
                     _4603 };
    assign _4605 = _4604 < _3518;
    assign _4606 = ~ _4605;
    assign _4594 = _4098[8:8];
    assign _4591 = _4586 - _3518;
    assign _4592 = _4588 ? _4591 : _4586;
    assign _4593 = _4592[62:0];
    assign _4595 = { _4593,
                     _4594 };
    assign _4596 = _4595 < _3518;
    assign _4597 = ~ _4596;
    assign _4585 = _4098[9:9];
    assign _4582 = _4577 - _3518;
    assign _4583 = _4579 ? _4582 : _4577;
    assign _4584 = _4583[62:0];
    assign _4586 = { _4584,
                     _4585 };
    assign _4587 = _4586 < _3518;
    assign _4588 = ~ _4587;
    assign _4576 = _4098[10:10];
    assign _4573 = _4568 - _3518;
    assign _4574 = _4570 ? _4573 : _4568;
    assign _4575 = _4574[62:0];
    assign _4577 = { _4575,
                     _4576 };
    assign _4578 = _4577 < _3518;
    assign _4579 = ~ _4578;
    assign _4567 = _4098[11:11];
    assign _4564 = _4559 - _3518;
    assign _4565 = _4561 ? _4564 : _4559;
    assign _4566 = _4565[62:0];
    assign _4568 = { _4566,
                     _4567 };
    assign _4569 = _4568 < _3518;
    assign _4570 = ~ _4569;
    assign _4558 = _4098[12:12];
    assign _4555 = _4550 - _3518;
    assign _4556 = _4552 ? _4555 : _4550;
    assign _4557 = _4556[62:0];
    assign _4559 = { _4557,
                     _4558 };
    assign _4560 = _4559 < _3518;
    assign _4561 = ~ _4560;
    assign _4549 = _4098[13:13];
    assign _4546 = _4541 - _3518;
    assign _4547 = _4543 ? _4546 : _4541;
    assign _4548 = _4547[62:0];
    assign _4550 = { _4548,
                     _4549 };
    assign _4551 = _4550 < _3518;
    assign _4552 = ~ _4551;
    assign _4540 = _4098[14:14];
    assign _4537 = _4532 - _3518;
    assign _4538 = _4534 ? _4537 : _4532;
    assign _4539 = _4538[62:0];
    assign _4541 = { _4539,
                     _4540 };
    assign _4542 = _4541 < _3518;
    assign _4543 = ~ _4542;
    assign _4531 = _4098[15:15];
    assign _4528 = _4523 - _3518;
    assign _4529 = _4525 ? _4528 : _4523;
    assign _4530 = _4529[62:0];
    assign _4532 = { _4530,
                     _4531 };
    assign _4533 = _4532 < _3518;
    assign _4534 = ~ _4533;
    assign _4522 = _4098[16:16];
    assign _4519 = _4514 - _3518;
    assign _4520 = _4516 ? _4519 : _4514;
    assign _4521 = _4520[62:0];
    assign _4523 = { _4521,
                     _4522 };
    assign _4524 = _4523 < _3518;
    assign _4525 = ~ _4524;
    assign _4513 = _4098[17:17];
    assign _4510 = _4505 - _3518;
    assign _4511 = _4507 ? _4510 : _4505;
    assign _4512 = _4511[62:0];
    assign _4514 = { _4512,
                     _4513 };
    assign _4515 = _4514 < _3518;
    assign _4516 = ~ _4515;
    assign _4504 = _4098[18:18];
    assign _4501 = _4496 - _3518;
    assign _4502 = _4498 ? _4501 : _4496;
    assign _4503 = _4502[62:0];
    assign _4505 = { _4503,
                     _4504 };
    assign _4506 = _4505 < _3518;
    assign _4507 = ~ _4506;
    assign _4495 = _4098[19:19];
    assign _4492 = _4487 - _3518;
    assign _4493 = _4489 ? _4492 : _4487;
    assign _4494 = _4493[62:0];
    assign _4496 = { _4494,
                     _4495 };
    assign _4497 = _4496 < _3518;
    assign _4498 = ~ _4497;
    assign _4486 = _4098[20:20];
    assign _4483 = _4478 - _3518;
    assign _4484 = _4480 ? _4483 : _4478;
    assign _4485 = _4484[62:0];
    assign _4487 = { _4485,
                     _4486 };
    assign _4488 = _4487 < _3518;
    assign _4489 = ~ _4488;
    assign _4477 = _4098[21:21];
    assign _4474 = _4469 - _3518;
    assign _4475 = _4471 ? _4474 : _4469;
    assign _4476 = _4475[62:0];
    assign _4478 = { _4476,
                     _4477 };
    assign _4479 = _4478 < _3518;
    assign _4480 = ~ _4479;
    assign _4468 = _4098[22:22];
    assign _4465 = _4460 - _3518;
    assign _4466 = _4462 ? _4465 : _4460;
    assign _4467 = _4466[62:0];
    assign _4469 = { _4467,
                     _4468 };
    assign _4470 = _4469 < _3518;
    assign _4471 = ~ _4470;
    assign _4459 = _4098[23:23];
    assign _4456 = _4451 - _3518;
    assign _4457 = _4453 ? _4456 : _4451;
    assign _4458 = _4457[62:0];
    assign _4460 = { _4458,
                     _4459 };
    assign _4461 = _4460 < _3518;
    assign _4462 = ~ _4461;
    assign _4450 = _4098[24:24];
    assign _4447 = _4442 - _3518;
    assign _4448 = _4444 ? _4447 : _4442;
    assign _4449 = _4448[62:0];
    assign _4451 = { _4449,
                     _4450 };
    assign _4452 = _4451 < _3518;
    assign _4453 = ~ _4452;
    assign _4441 = _4098[25:25];
    assign _4438 = _4433 - _3518;
    assign _4439 = _4435 ? _4438 : _4433;
    assign _4440 = _4439[62:0];
    assign _4442 = { _4440,
                     _4441 };
    assign _4443 = _4442 < _3518;
    assign _4444 = ~ _4443;
    assign _4432 = _4098[26:26];
    assign _4429 = _4424 - _3518;
    assign _4430 = _4426 ? _4429 : _4424;
    assign _4431 = _4430[62:0];
    assign _4433 = { _4431,
                     _4432 };
    assign _4434 = _4433 < _3518;
    assign _4435 = ~ _4434;
    assign _4423 = _4098[27:27];
    assign _4420 = _4415 - _3518;
    assign _4421 = _4417 ? _4420 : _4415;
    assign _4422 = _4421[62:0];
    assign _4424 = { _4422,
                     _4423 };
    assign _4425 = _4424 < _3518;
    assign _4426 = ~ _4425;
    assign _4414 = _4098[28:28];
    assign _4411 = _4406 - _3518;
    assign _4412 = _4408 ? _4411 : _4406;
    assign _4413 = _4412[62:0];
    assign _4415 = { _4413,
                     _4414 };
    assign _4416 = _4415 < _3518;
    assign _4417 = ~ _4416;
    assign _4405 = _4098[29:29];
    assign _4402 = _4397 - _3518;
    assign _4403 = _4399 ? _4402 : _4397;
    assign _4404 = _4403[62:0];
    assign _4406 = { _4404,
                     _4405 };
    assign _4407 = _4406 < _3518;
    assign _4408 = ~ _4407;
    assign _4396 = _4098[30:30];
    assign _4393 = _4388 - _3518;
    assign _4394 = _4390 ? _4393 : _4388;
    assign _4395 = _4394[62:0];
    assign _4397 = { _4395,
                     _4396 };
    assign _4398 = _4397 < _3518;
    assign _4399 = ~ _4398;
    assign _4387 = _4098[31:31];
    assign _4384 = _4379 - _3518;
    assign _4385 = _4381 ? _4384 : _4379;
    assign _4386 = _4385[62:0];
    assign _4388 = { _4386,
                     _4387 };
    assign _4389 = _4388 < _3518;
    assign _4390 = ~ _4389;
    assign _4378 = _4098[32:32];
    assign _4375 = _4370 - _3518;
    assign _4376 = _4372 ? _4375 : _4370;
    assign _4377 = _4376[62:0];
    assign _4379 = { _4377,
                     _4378 };
    assign _4380 = _4379 < _3518;
    assign _4381 = ~ _4380;
    assign _4369 = _4098[33:33];
    assign _4366 = _4361 - _3518;
    assign _4367 = _4363 ? _4366 : _4361;
    assign _4368 = _4367[62:0];
    assign _4370 = { _4368,
                     _4369 };
    assign _4371 = _4370 < _3518;
    assign _4372 = ~ _4371;
    assign _4360 = _4098[34:34];
    assign _4357 = _4352 - _3518;
    assign _4358 = _4354 ? _4357 : _4352;
    assign _4359 = _4358[62:0];
    assign _4361 = { _4359,
                     _4360 };
    assign _4362 = _4361 < _3518;
    assign _4363 = ~ _4362;
    assign _4351 = _4098[35:35];
    assign _4348 = _4343 - _3518;
    assign _4349 = _4345 ? _4348 : _4343;
    assign _4350 = _4349[62:0];
    assign _4352 = { _4350,
                     _4351 };
    assign _4353 = _4352 < _3518;
    assign _4354 = ~ _4353;
    assign _4342 = _4098[36:36];
    assign _4339 = _4334 - _3518;
    assign _4340 = _4336 ? _4339 : _4334;
    assign _4341 = _4340[62:0];
    assign _4343 = { _4341,
                     _4342 };
    assign _4344 = _4343 < _3518;
    assign _4345 = ~ _4344;
    assign _4333 = _4098[37:37];
    assign _4330 = _4325 - _3518;
    assign _4331 = _4327 ? _4330 : _4325;
    assign _4332 = _4331[62:0];
    assign _4334 = { _4332,
                     _4333 };
    assign _4335 = _4334 < _3518;
    assign _4336 = ~ _4335;
    assign _4324 = _4098[38:38];
    assign _4321 = _4316 - _3518;
    assign _4322 = _4318 ? _4321 : _4316;
    assign _4323 = _4322[62:0];
    assign _4325 = { _4323,
                     _4324 };
    assign _4326 = _4325 < _3518;
    assign _4327 = ~ _4326;
    assign _4315 = _4098[39:39];
    assign _4312 = _4307 - _3518;
    assign _4313 = _4309 ? _4312 : _4307;
    assign _4314 = _4313[62:0];
    assign _4316 = { _4314,
                     _4315 };
    assign _4317 = _4316 < _3518;
    assign _4318 = ~ _4317;
    assign _4306 = _4098[40:40];
    assign _4303 = _4298 - _3518;
    assign _4304 = _4300 ? _4303 : _4298;
    assign _4305 = _4304[62:0];
    assign _4307 = { _4305,
                     _4306 };
    assign _4308 = _4307 < _3518;
    assign _4309 = ~ _4308;
    assign _4297 = _4098[41:41];
    assign _4294 = _4289 - _3518;
    assign _4295 = _4291 ? _4294 : _4289;
    assign _4296 = _4295[62:0];
    assign _4298 = { _4296,
                     _4297 };
    assign _4299 = _4298 < _3518;
    assign _4300 = ~ _4299;
    assign _4288 = _4098[42:42];
    assign _4285 = _4280 - _3518;
    assign _4286 = _4282 ? _4285 : _4280;
    assign _4287 = _4286[62:0];
    assign _4289 = { _4287,
                     _4288 };
    assign _4290 = _4289 < _3518;
    assign _4291 = ~ _4290;
    assign _4279 = _4098[43:43];
    assign _4276 = _4271 - _3518;
    assign _4277 = _4273 ? _4276 : _4271;
    assign _4278 = _4277[62:0];
    assign _4280 = { _4278,
                     _4279 };
    assign _4281 = _4280 < _3518;
    assign _4282 = ~ _4281;
    assign _4270 = _4098[44:44];
    assign _4267 = _4262 - _3518;
    assign _4268 = _4264 ? _4267 : _4262;
    assign _4269 = _4268[62:0];
    assign _4271 = { _4269,
                     _4270 };
    assign _4272 = _4271 < _3518;
    assign _4273 = ~ _4272;
    assign _4261 = _4098[45:45];
    assign _4258 = _4253 - _3518;
    assign _4259 = _4255 ? _4258 : _4253;
    assign _4260 = _4259[62:0];
    assign _4262 = { _4260,
                     _4261 };
    assign _4263 = _4262 < _3518;
    assign _4264 = ~ _4263;
    assign _4252 = _4098[46:46];
    assign _4249 = _4244 - _3518;
    assign _4250 = _4246 ? _4249 : _4244;
    assign _4251 = _4250[62:0];
    assign _4253 = { _4251,
                     _4252 };
    assign _4254 = _4253 < _3518;
    assign _4255 = ~ _4254;
    assign _4243 = _4098[47:47];
    assign _4240 = _4235 - _3518;
    assign _4241 = _4237 ? _4240 : _4235;
    assign _4242 = _4241[62:0];
    assign _4244 = { _4242,
                     _4243 };
    assign _4245 = _4244 < _3518;
    assign _4246 = ~ _4245;
    assign _4234 = _4098[48:48];
    assign _4231 = _4226 - _3518;
    assign _4232 = _4228 ? _4231 : _4226;
    assign _4233 = _4232[62:0];
    assign _4235 = { _4233,
                     _4234 };
    assign _4236 = _4235 < _3518;
    assign _4237 = ~ _4236;
    assign _4225 = _4098[49:49];
    assign _4222 = _4217 - _3518;
    assign _4223 = _4219 ? _4222 : _4217;
    assign _4224 = _4223[62:0];
    assign _4226 = { _4224,
                     _4225 };
    assign _4227 = _4226 < _3518;
    assign _4228 = ~ _4227;
    assign _4216 = _4098[50:50];
    assign _4213 = _4208 - _3518;
    assign _4214 = _4210 ? _4213 : _4208;
    assign _4215 = _4214[62:0];
    assign _4217 = { _4215,
                     _4216 };
    assign _4218 = _4217 < _3518;
    assign _4219 = ~ _4218;
    assign _4207 = _4098[51:51];
    assign _4204 = _4199 - _3518;
    assign _4205 = _4201 ? _4204 : _4199;
    assign _4206 = _4205[62:0];
    assign _4208 = { _4206,
                     _4207 };
    assign _4209 = _4208 < _3518;
    assign _4210 = ~ _4209;
    assign _4198 = _4098[52:52];
    assign _4195 = _4190 - _3518;
    assign _4196 = _4192 ? _4195 : _4190;
    assign _4197 = _4196[62:0];
    assign _4199 = { _4197,
                     _4198 };
    assign _4200 = _4199 < _3518;
    assign _4201 = ~ _4200;
    assign _4189 = _4098[53:53];
    assign _4186 = _4181 - _3518;
    assign _4187 = _4183 ? _4186 : _4181;
    assign _4188 = _4187[62:0];
    assign _4190 = { _4188,
                     _4189 };
    assign _4191 = _4190 < _3518;
    assign _4192 = ~ _4191;
    assign _4180 = _4098[54:54];
    assign _4177 = _4172 - _3518;
    assign _4178 = _4174 ? _4177 : _4172;
    assign _4179 = _4178[62:0];
    assign _4181 = { _4179,
                     _4180 };
    assign _4182 = _4181 < _3518;
    assign _4183 = ~ _4182;
    assign _4171 = _4098[55:55];
    assign _4168 = _4163 - _3518;
    assign _4169 = _4165 ? _4168 : _4163;
    assign _4170 = _4169[62:0];
    assign _4172 = { _4170,
                     _4171 };
    assign _4173 = _4172 < _3518;
    assign _4174 = ~ _4173;
    assign _4162 = _4098[56:56];
    assign _4159 = _4154 - _3518;
    assign _4160 = _4156 ? _4159 : _4154;
    assign _4161 = _4160[62:0];
    assign _4163 = { _4161,
                     _4162 };
    assign _4164 = _4163 < _3518;
    assign _4165 = ~ _4164;
    assign _4153 = _4098[57:57];
    assign _4150 = _4145 - _3518;
    assign _4151 = _4147 ? _4150 : _4145;
    assign _4152 = _4151[62:0];
    assign _4154 = { _4152,
                     _4153 };
    assign _4155 = _4154 < _3518;
    assign _4156 = ~ _4155;
    assign _4144 = _4098[58:58];
    assign _4141 = _4136 - _3518;
    assign _4142 = _4138 ? _4141 : _4136;
    assign _4143 = _4142[62:0];
    assign _4145 = { _4143,
                     _4144 };
    assign _4146 = _4145 < _3518;
    assign _4147 = ~ _4146;
    assign _4135 = _4098[59:59];
    assign _4132 = _4127 - _3518;
    assign _4133 = _4129 ? _4132 : _4127;
    assign _4134 = _4133[62:0];
    assign _4136 = { _4134,
                     _4135 };
    assign _4137 = _4136 < _3518;
    assign _4138 = ~ _4137;
    assign _4126 = _4098[60:60];
    assign _4123 = _4118 - _3518;
    assign _4124 = _4120 ? _4123 : _4118;
    assign _4125 = _4124[62:0];
    assign _4127 = { _4125,
                     _4126 };
    assign _4128 = _4127 < _3518;
    assign _4129 = ~ _4128;
    assign _4117 = _4098[61:61];
    assign _4114 = _4109 - _3518;
    assign _4115 = _4111 ? _4114 : _4109;
    assign _4116 = _4115[62:0];
    assign _4118 = { _4116,
                     _4117 };
    assign _4119 = _4118 < _3518;
    assign _4120 = ~ _4119;
    assign _4108 = _4098[62:62];
    assign _4105 = _4100 - _3518;
    assign _4106 = _4102 ? _4105 : _4100;
    assign _4107 = _4106[62:0];
    assign _4109 = { _4107,
                     _4108 };
    assign _4110 = _4109 < _3518;
    assign _4111 = ~ _4110;
    assign _4098 = _3510 - _4092;
    assign _4099 = _4098[63:63];
    assign _4100 = { _22185,
                     _4099 };
    assign _4101 = _4100 < _3518;
    assign _4102 = ~ _4101;
    assign _4103 = { _22185,
                     _4102 };
    assign _4104 = _4103[62:0];
    assign _4112 = { _4104,
                     _4111 };
    assign _4113 = _4112[62:0];
    assign _4121 = { _4113,
                     _4120 };
    assign _4122 = _4121[62:0];
    assign _4130 = { _4122,
                     _4129 };
    assign _4131 = _4130[62:0];
    assign _4139 = { _4131,
                     _4138 };
    assign _4140 = _4139[62:0];
    assign _4148 = { _4140,
                     _4147 };
    assign _4149 = _4148[62:0];
    assign _4157 = { _4149,
                     _4156 };
    assign _4158 = _4157[62:0];
    assign _4166 = { _4158,
                     _4165 };
    assign _4167 = _4166[62:0];
    assign _4175 = { _4167,
                     _4174 };
    assign _4176 = _4175[62:0];
    assign _4184 = { _4176,
                     _4183 };
    assign _4185 = _4184[62:0];
    assign _4193 = { _4185,
                     _4192 };
    assign _4194 = _4193[62:0];
    assign _4202 = { _4194,
                     _4201 };
    assign _4203 = _4202[62:0];
    assign _4211 = { _4203,
                     _4210 };
    assign _4212 = _4211[62:0];
    assign _4220 = { _4212,
                     _4219 };
    assign _4221 = _4220[62:0];
    assign _4229 = { _4221,
                     _4228 };
    assign _4230 = _4229[62:0];
    assign _4238 = { _4230,
                     _4237 };
    assign _4239 = _4238[62:0];
    assign _4247 = { _4239,
                     _4246 };
    assign _4248 = _4247[62:0];
    assign _4256 = { _4248,
                     _4255 };
    assign _4257 = _4256[62:0];
    assign _4265 = { _4257,
                     _4264 };
    assign _4266 = _4265[62:0];
    assign _4274 = { _4266,
                     _4273 };
    assign _4275 = _4274[62:0];
    assign _4283 = { _4275,
                     _4282 };
    assign _4284 = _4283[62:0];
    assign _4292 = { _4284,
                     _4291 };
    assign _4293 = _4292[62:0];
    assign _4301 = { _4293,
                     _4300 };
    assign _4302 = _4301[62:0];
    assign _4310 = { _4302,
                     _4309 };
    assign _4311 = _4310[62:0];
    assign _4319 = { _4311,
                     _4318 };
    assign _4320 = _4319[62:0];
    assign _4328 = { _4320,
                     _4327 };
    assign _4329 = _4328[62:0];
    assign _4337 = { _4329,
                     _4336 };
    assign _4338 = _4337[62:0];
    assign _4346 = { _4338,
                     _4345 };
    assign _4347 = _4346[62:0];
    assign _4355 = { _4347,
                     _4354 };
    assign _4356 = _4355[62:0];
    assign _4364 = { _4356,
                     _4363 };
    assign _4365 = _4364[62:0];
    assign _4373 = { _4365,
                     _4372 };
    assign _4374 = _4373[62:0];
    assign _4382 = { _4374,
                     _4381 };
    assign _4383 = _4382[62:0];
    assign _4391 = { _4383,
                     _4390 };
    assign _4392 = _4391[62:0];
    assign _4400 = { _4392,
                     _4399 };
    assign _4401 = _4400[62:0];
    assign _4409 = { _4401,
                     _4408 };
    assign _4410 = _4409[62:0];
    assign _4418 = { _4410,
                     _4417 };
    assign _4419 = _4418[62:0];
    assign _4427 = { _4419,
                     _4426 };
    assign _4428 = _4427[62:0];
    assign _4436 = { _4428,
                     _4435 };
    assign _4437 = _4436[62:0];
    assign _4445 = { _4437,
                     _4444 };
    assign _4446 = _4445[62:0];
    assign _4454 = { _4446,
                     _4453 };
    assign _4455 = _4454[62:0];
    assign _4463 = { _4455,
                     _4462 };
    assign _4464 = _4463[62:0];
    assign _4472 = { _4464,
                     _4471 };
    assign _4473 = _4472[62:0];
    assign _4481 = { _4473,
                     _4480 };
    assign _4482 = _4481[62:0];
    assign _4490 = { _4482,
                     _4489 };
    assign _4491 = _4490[62:0];
    assign _4499 = { _4491,
                     _4498 };
    assign _4500 = _4499[62:0];
    assign _4508 = { _4500,
                     _4507 };
    assign _4509 = _4508[62:0];
    assign _4517 = { _4509,
                     _4516 };
    assign _4518 = _4517[62:0];
    assign _4526 = { _4518,
                     _4525 };
    assign _4527 = _4526[62:0];
    assign _4535 = { _4527,
                     _4534 };
    assign _4536 = _4535[62:0];
    assign _4544 = { _4536,
                     _4543 };
    assign _4545 = _4544[62:0];
    assign _4553 = { _4545,
                     _4552 };
    assign _4554 = _4553[62:0];
    assign _4562 = { _4554,
                     _4561 };
    assign _4563 = _4562[62:0];
    assign _4571 = { _4563,
                     _4570 };
    assign _4572 = _4571[62:0];
    assign _4580 = { _4572,
                     _4579 };
    assign _4581 = _4580[62:0];
    assign _4589 = { _4581,
                     _4588 };
    assign _4590 = _4589[62:0];
    assign _4598 = { _4590,
                     _4597 };
    assign _4599 = _4598[62:0];
    assign _4607 = { _4599,
                     _4606 };
    assign _4608 = _4607[62:0];
    assign _4616 = { _4608,
                     _4615 };
    assign _4617 = _4616[62:0];
    assign _4625 = { _4617,
                     _4624 };
    assign _4626 = _4625[62:0];
    assign _4634 = { _4626,
                     _4633 };
    assign _4635 = _4634[62:0];
    assign _4643 = { _4635,
                     _4642 };
    assign _4644 = _4643[62:0];
    assign _4652 = { _4644,
                     _4651 };
    assign _4653 = _4652[62:0];
    assign _4661 = { _4653,
                     _4660 };
    assign _4662 = _4661[62:0];
    assign _4670 = { _4662,
                     _4669 };
    assign _4672 = _4670 + _22186;
    assign _4673 = _4672 * _4092;
    assign _4674 = _4673[63:0];
    assign _5256 = _4674 + _5255;
    assign _4084 = _3515[0:0];
    assign _4081 = _4076 - _3518;
    assign _4082 = _4078 ? _4081 : _4076;
    assign _4083 = _4082[62:0];
    assign _4085 = { _4083,
                     _4084 };
    assign _4086 = _4085 < _3518;
    assign _4087 = ~ _4086;
    assign _4075 = _3515[1:1];
    assign _4072 = _4067 - _3518;
    assign _4073 = _4069 ? _4072 : _4067;
    assign _4074 = _4073[62:0];
    assign _4076 = { _4074,
                     _4075 };
    assign _4077 = _4076 < _3518;
    assign _4078 = ~ _4077;
    assign _4066 = _3515[2:2];
    assign _4063 = _4058 - _3518;
    assign _4064 = _4060 ? _4063 : _4058;
    assign _4065 = _4064[62:0];
    assign _4067 = { _4065,
                     _4066 };
    assign _4068 = _4067 < _3518;
    assign _4069 = ~ _4068;
    assign _4057 = _3515[3:3];
    assign _4054 = _4049 - _3518;
    assign _4055 = _4051 ? _4054 : _4049;
    assign _4056 = _4055[62:0];
    assign _4058 = { _4056,
                     _4057 };
    assign _4059 = _4058 < _3518;
    assign _4060 = ~ _4059;
    assign _4048 = _3515[4:4];
    assign _4045 = _4040 - _3518;
    assign _4046 = _4042 ? _4045 : _4040;
    assign _4047 = _4046[62:0];
    assign _4049 = { _4047,
                     _4048 };
    assign _4050 = _4049 < _3518;
    assign _4051 = ~ _4050;
    assign _4039 = _3515[5:5];
    assign _4036 = _4031 - _3518;
    assign _4037 = _4033 ? _4036 : _4031;
    assign _4038 = _4037[62:0];
    assign _4040 = { _4038,
                     _4039 };
    assign _4041 = _4040 < _3518;
    assign _4042 = ~ _4041;
    assign _4030 = _3515[6:6];
    assign _4027 = _4022 - _3518;
    assign _4028 = _4024 ? _4027 : _4022;
    assign _4029 = _4028[62:0];
    assign _4031 = { _4029,
                     _4030 };
    assign _4032 = _4031 < _3518;
    assign _4033 = ~ _4032;
    assign _4021 = _3515[7:7];
    assign _4018 = _4013 - _3518;
    assign _4019 = _4015 ? _4018 : _4013;
    assign _4020 = _4019[62:0];
    assign _4022 = { _4020,
                     _4021 };
    assign _4023 = _4022 < _3518;
    assign _4024 = ~ _4023;
    assign _4012 = _3515[8:8];
    assign _4009 = _4004 - _3518;
    assign _4010 = _4006 ? _4009 : _4004;
    assign _4011 = _4010[62:0];
    assign _4013 = { _4011,
                     _4012 };
    assign _4014 = _4013 < _3518;
    assign _4015 = ~ _4014;
    assign _4003 = _3515[9:9];
    assign _4000 = _3995 - _3518;
    assign _4001 = _3997 ? _4000 : _3995;
    assign _4002 = _4001[62:0];
    assign _4004 = { _4002,
                     _4003 };
    assign _4005 = _4004 < _3518;
    assign _4006 = ~ _4005;
    assign _3994 = _3515[10:10];
    assign _3991 = _3986 - _3518;
    assign _3992 = _3988 ? _3991 : _3986;
    assign _3993 = _3992[62:0];
    assign _3995 = { _3993,
                     _3994 };
    assign _3996 = _3995 < _3518;
    assign _3997 = ~ _3996;
    assign _3985 = _3515[11:11];
    assign _3982 = _3977 - _3518;
    assign _3983 = _3979 ? _3982 : _3977;
    assign _3984 = _3983[62:0];
    assign _3986 = { _3984,
                     _3985 };
    assign _3987 = _3986 < _3518;
    assign _3988 = ~ _3987;
    assign _3976 = _3515[12:12];
    assign _3973 = _3968 - _3518;
    assign _3974 = _3970 ? _3973 : _3968;
    assign _3975 = _3974[62:0];
    assign _3977 = { _3975,
                     _3976 };
    assign _3978 = _3977 < _3518;
    assign _3979 = ~ _3978;
    assign _3967 = _3515[13:13];
    assign _3964 = _3959 - _3518;
    assign _3965 = _3961 ? _3964 : _3959;
    assign _3966 = _3965[62:0];
    assign _3968 = { _3966,
                     _3967 };
    assign _3969 = _3968 < _3518;
    assign _3970 = ~ _3969;
    assign _3958 = _3515[14:14];
    assign _3955 = _3950 - _3518;
    assign _3956 = _3952 ? _3955 : _3950;
    assign _3957 = _3956[62:0];
    assign _3959 = { _3957,
                     _3958 };
    assign _3960 = _3959 < _3518;
    assign _3961 = ~ _3960;
    assign _3949 = _3515[15:15];
    assign _3946 = _3941 - _3518;
    assign _3947 = _3943 ? _3946 : _3941;
    assign _3948 = _3947[62:0];
    assign _3950 = { _3948,
                     _3949 };
    assign _3951 = _3950 < _3518;
    assign _3952 = ~ _3951;
    assign _3940 = _3515[16:16];
    assign _3937 = _3932 - _3518;
    assign _3938 = _3934 ? _3937 : _3932;
    assign _3939 = _3938[62:0];
    assign _3941 = { _3939,
                     _3940 };
    assign _3942 = _3941 < _3518;
    assign _3943 = ~ _3942;
    assign _3931 = _3515[17:17];
    assign _3928 = _3923 - _3518;
    assign _3929 = _3925 ? _3928 : _3923;
    assign _3930 = _3929[62:0];
    assign _3932 = { _3930,
                     _3931 };
    assign _3933 = _3932 < _3518;
    assign _3934 = ~ _3933;
    assign _3922 = _3515[18:18];
    assign _3919 = _3914 - _3518;
    assign _3920 = _3916 ? _3919 : _3914;
    assign _3921 = _3920[62:0];
    assign _3923 = { _3921,
                     _3922 };
    assign _3924 = _3923 < _3518;
    assign _3925 = ~ _3924;
    assign _3913 = _3515[19:19];
    assign _3910 = _3905 - _3518;
    assign _3911 = _3907 ? _3910 : _3905;
    assign _3912 = _3911[62:0];
    assign _3914 = { _3912,
                     _3913 };
    assign _3915 = _3914 < _3518;
    assign _3916 = ~ _3915;
    assign _3904 = _3515[20:20];
    assign _3901 = _3896 - _3518;
    assign _3902 = _3898 ? _3901 : _3896;
    assign _3903 = _3902[62:0];
    assign _3905 = { _3903,
                     _3904 };
    assign _3906 = _3905 < _3518;
    assign _3907 = ~ _3906;
    assign _3895 = _3515[21:21];
    assign _3892 = _3887 - _3518;
    assign _3893 = _3889 ? _3892 : _3887;
    assign _3894 = _3893[62:0];
    assign _3896 = { _3894,
                     _3895 };
    assign _3897 = _3896 < _3518;
    assign _3898 = ~ _3897;
    assign _3886 = _3515[22:22];
    assign _3883 = _3878 - _3518;
    assign _3884 = _3880 ? _3883 : _3878;
    assign _3885 = _3884[62:0];
    assign _3887 = { _3885,
                     _3886 };
    assign _3888 = _3887 < _3518;
    assign _3889 = ~ _3888;
    assign _3877 = _3515[23:23];
    assign _3874 = _3869 - _3518;
    assign _3875 = _3871 ? _3874 : _3869;
    assign _3876 = _3875[62:0];
    assign _3878 = { _3876,
                     _3877 };
    assign _3879 = _3878 < _3518;
    assign _3880 = ~ _3879;
    assign _3868 = _3515[24:24];
    assign _3865 = _3860 - _3518;
    assign _3866 = _3862 ? _3865 : _3860;
    assign _3867 = _3866[62:0];
    assign _3869 = { _3867,
                     _3868 };
    assign _3870 = _3869 < _3518;
    assign _3871 = ~ _3870;
    assign _3859 = _3515[25:25];
    assign _3856 = _3851 - _3518;
    assign _3857 = _3853 ? _3856 : _3851;
    assign _3858 = _3857[62:0];
    assign _3860 = { _3858,
                     _3859 };
    assign _3861 = _3860 < _3518;
    assign _3862 = ~ _3861;
    assign _3850 = _3515[26:26];
    assign _3847 = _3842 - _3518;
    assign _3848 = _3844 ? _3847 : _3842;
    assign _3849 = _3848[62:0];
    assign _3851 = { _3849,
                     _3850 };
    assign _3852 = _3851 < _3518;
    assign _3853 = ~ _3852;
    assign _3841 = _3515[27:27];
    assign _3838 = _3833 - _3518;
    assign _3839 = _3835 ? _3838 : _3833;
    assign _3840 = _3839[62:0];
    assign _3842 = { _3840,
                     _3841 };
    assign _3843 = _3842 < _3518;
    assign _3844 = ~ _3843;
    assign _3832 = _3515[28:28];
    assign _3829 = _3824 - _3518;
    assign _3830 = _3826 ? _3829 : _3824;
    assign _3831 = _3830[62:0];
    assign _3833 = { _3831,
                     _3832 };
    assign _3834 = _3833 < _3518;
    assign _3835 = ~ _3834;
    assign _3823 = _3515[29:29];
    assign _3820 = _3815 - _3518;
    assign _3821 = _3817 ? _3820 : _3815;
    assign _3822 = _3821[62:0];
    assign _3824 = { _3822,
                     _3823 };
    assign _3825 = _3824 < _3518;
    assign _3826 = ~ _3825;
    assign _3814 = _3515[30:30];
    assign _3811 = _3806 - _3518;
    assign _3812 = _3808 ? _3811 : _3806;
    assign _3813 = _3812[62:0];
    assign _3815 = { _3813,
                     _3814 };
    assign _3816 = _3815 < _3518;
    assign _3817 = ~ _3816;
    assign _3805 = _3515[31:31];
    assign _3802 = _3797 - _3518;
    assign _3803 = _3799 ? _3802 : _3797;
    assign _3804 = _3803[62:0];
    assign _3806 = { _3804,
                     _3805 };
    assign _3807 = _3806 < _3518;
    assign _3808 = ~ _3807;
    assign _3796 = _3515[32:32];
    assign _3793 = _3788 - _3518;
    assign _3794 = _3790 ? _3793 : _3788;
    assign _3795 = _3794[62:0];
    assign _3797 = { _3795,
                     _3796 };
    assign _3798 = _3797 < _3518;
    assign _3799 = ~ _3798;
    assign _3787 = _3515[33:33];
    assign _3784 = _3779 - _3518;
    assign _3785 = _3781 ? _3784 : _3779;
    assign _3786 = _3785[62:0];
    assign _3788 = { _3786,
                     _3787 };
    assign _3789 = _3788 < _3518;
    assign _3790 = ~ _3789;
    assign _3778 = _3515[34:34];
    assign _3775 = _3770 - _3518;
    assign _3776 = _3772 ? _3775 : _3770;
    assign _3777 = _3776[62:0];
    assign _3779 = { _3777,
                     _3778 };
    assign _3780 = _3779 < _3518;
    assign _3781 = ~ _3780;
    assign _3769 = _3515[35:35];
    assign _3766 = _3761 - _3518;
    assign _3767 = _3763 ? _3766 : _3761;
    assign _3768 = _3767[62:0];
    assign _3770 = { _3768,
                     _3769 };
    assign _3771 = _3770 < _3518;
    assign _3772 = ~ _3771;
    assign _3760 = _3515[36:36];
    assign _3757 = _3752 - _3518;
    assign _3758 = _3754 ? _3757 : _3752;
    assign _3759 = _3758[62:0];
    assign _3761 = { _3759,
                     _3760 };
    assign _3762 = _3761 < _3518;
    assign _3763 = ~ _3762;
    assign _3751 = _3515[37:37];
    assign _3748 = _3743 - _3518;
    assign _3749 = _3745 ? _3748 : _3743;
    assign _3750 = _3749[62:0];
    assign _3752 = { _3750,
                     _3751 };
    assign _3753 = _3752 < _3518;
    assign _3754 = ~ _3753;
    assign _3742 = _3515[38:38];
    assign _3739 = _3734 - _3518;
    assign _3740 = _3736 ? _3739 : _3734;
    assign _3741 = _3740[62:0];
    assign _3743 = { _3741,
                     _3742 };
    assign _3744 = _3743 < _3518;
    assign _3745 = ~ _3744;
    assign _3733 = _3515[39:39];
    assign _3730 = _3725 - _3518;
    assign _3731 = _3727 ? _3730 : _3725;
    assign _3732 = _3731[62:0];
    assign _3734 = { _3732,
                     _3733 };
    assign _3735 = _3734 < _3518;
    assign _3736 = ~ _3735;
    assign _3724 = _3515[40:40];
    assign _3721 = _3716 - _3518;
    assign _3722 = _3718 ? _3721 : _3716;
    assign _3723 = _3722[62:0];
    assign _3725 = { _3723,
                     _3724 };
    assign _3726 = _3725 < _3518;
    assign _3727 = ~ _3726;
    assign _3715 = _3515[41:41];
    assign _3712 = _3707 - _3518;
    assign _3713 = _3709 ? _3712 : _3707;
    assign _3714 = _3713[62:0];
    assign _3716 = { _3714,
                     _3715 };
    assign _3717 = _3716 < _3518;
    assign _3718 = ~ _3717;
    assign _3706 = _3515[42:42];
    assign _3703 = _3698 - _3518;
    assign _3704 = _3700 ? _3703 : _3698;
    assign _3705 = _3704[62:0];
    assign _3707 = { _3705,
                     _3706 };
    assign _3708 = _3707 < _3518;
    assign _3709 = ~ _3708;
    assign _3697 = _3515[43:43];
    assign _3694 = _3689 - _3518;
    assign _3695 = _3691 ? _3694 : _3689;
    assign _3696 = _3695[62:0];
    assign _3698 = { _3696,
                     _3697 };
    assign _3699 = _3698 < _3518;
    assign _3700 = ~ _3699;
    assign _3688 = _3515[44:44];
    assign _3685 = _3680 - _3518;
    assign _3686 = _3682 ? _3685 : _3680;
    assign _3687 = _3686[62:0];
    assign _3689 = { _3687,
                     _3688 };
    assign _3690 = _3689 < _3518;
    assign _3691 = ~ _3690;
    assign _3679 = _3515[45:45];
    assign _3676 = _3671 - _3518;
    assign _3677 = _3673 ? _3676 : _3671;
    assign _3678 = _3677[62:0];
    assign _3680 = { _3678,
                     _3679 };
    assign _3681 = _3680 < _3518;
    assign _3682 = ~ _3681;
    assign _3670 = _3515[46:46];
    assign _3667 = _3662 - _3518;
    assign _3668 = _3664 ? _3667 : _3662;
    assign _3669 = _3668[62:0];
    assign _3671 = { _3669,
                     _3670 };
    assign _3672 = _3671 < _3518;
    assign _3673 = ~ _3672;
    assign _3661 = _3515[47:47];
    assign _3658 = _3653 - _3518;
    assign _3659 = _3655 ? _3658 : _3653;
    assign _3660 = _3659[62:0];
    assign _3662 = { _3660,
                     _3661 };
    assign _3663 = _3662 < _3518;
    assign _3664 = ~ _3663;
    assign _3652 = _3515[48:48];
    assign _3649 = _3644 - _3518;
    assign _3650 = _3646 ? _3649 : _3644;
    assign _3651 = _3650[62:0];
    assign _3653 = { _3651,
                     _3652 };
    assign _3654 = _3653 < _3518;
    assign _3655 = ~ _3654;
    assign _3643 = _3515[49:49];
    assign _3640 = _3635 - _3518;
    assign _3641 = _3637 ? _3640 : _3635;
    assign _3642 = _3641[62:0];
    assign _3644 = { _3642,
                     _3643 };
    assign _3645 = _3644 < _3518;
    assign _3646 = ~ _3645;
    assign _3634 = _3515[50:50];
    assign _3631 = _3626 - _3518;
    assign _3632 = _3628 ? _3631 : _3626;
    assign _3633 = _3632[62:0];
    assign _3635 = { _3633,
                     _3634 };
    assign _3636 = _3635 < _3518;
    assign _3637 = ~ _3636;
    assign _3625 = _3515[51:51];
    assign _3622 = _3617 - _3518;
    assign _3623 = _3619 ? _3622 : _3617;
    assign _3624 = _3623[62:0];
    assign _3626 = { _3624,
                     _3625 };
    assign _3627 = _3626 < _3518;
    assign _3628 = ~ _3627;
    assign _3616 = _3515[52:52];
    assign _3613 = _3608 - _3518;
    assign _3614 = _3610 ? _3613 : _3608;
    assign _3615 = _3614[62:0];
    assign _3617 = { _3615,
                     _3616 };
    assign _3618 = _3617 < _3518;
    assign _3619 = ~ _3618;
    assign _3607 = _3515[53:53];
    assign _3604 = _3599 - _3518;
    assign _3605 = _3601 ? _3604 : _3599;
    assign _3606 = _3605[62:0];
    assign _3608 = { _3606,
                     _3607 };
    assign _3609 = _3608 < _3518;
    assign _3610 = ~ _3609;
    assign _3598 = _3515[54:54];
    assign _3595 = _3590 - _3518;
    assign _3596 = _3592 ? _3595 : _3590;
    assign _3597 = _3596[62:0];
    assign _3599 = { _3597,
                     _3598 };
    assign _3600 = _3599 < _3518;
    assign _3601 = ~ _3600;
    assign _3589 = _3515[55:55];
    assign _3586 = _3581 - _3518;
    assign _3587 = _3583 ? _3586 : _3581;
    assign _3588 = _3587[62:0];
    assign _3590 = { _3588,
                     _3589 };
    assign _3591 = _3590 < _3518;
    assign _3592 = ~ _3591;
    assign _3580 = _3515[56:56];
    assign _3577 = _3572 - _3518;
    assign _3578 = _3574 ? _3577 : _3572;
    assign _3579 = _3578[62:0];
    assign _3581 = { _3579,
                     _3580 };
    assign _3582 = _3581 < _3518;
    assign _3583 = ~ _3582;
    assign _3571 = _3515[57:57];
    assign _3568 = _3563 - _3518;
    assign _3569 = _3565 ? _3568 : _3563;
    assign _3570 = _3569[62:0];
    assign _3572 = { _3570,
                     _3571 };
    assign _3573 = _3572 < _3518;
    assign _3574 = ~ _3573;
    assign _3562 = _3515[58:58];
    assign _3559 = _3554 - _3518;
    assign _3560 = _3556 ? _3559 : _3554;
    assign _3561 = _3560[62:0];
    assign _3563 = { _3561,
                     _3562 };
    assign _3564 = _3563 < _3518;
    assign _3565 = ~ _3564;
    assign _3553 = _3515[59:59];
    assign _3550 = _3545 - _3518;
    assign _3551 = _3547 ? _3550 : _3545;
    assign _3552 = _3551[62:0];
    assign _3554 = { _3552,
                     _3553 };
    assign _3555 = _3554 < _3518;
    assign _3556 = ~ _3555;
    assign _3544 = _3515[60:60];
    assign _3541 = _3536 - _3518;
    assign _3542 = _3538 ? _3541 : _3536;
    assign _3543 = _3542[62:0];
    assign _3545 = { _3543,
                     _3544 };
    assign _3546 = _3545 < _3518;
    assign _3547 = ~ _3546;
    assign _3535 = _3515[61:61];
    assign _3532 = _3527 - _3518;
    assign _3533 = _3529 ? _3532 : _3527;
    assign _3534 = _3533[62:0];
    assign _3536 = { _3534,
                     _3535 };
    assign _3537 = _3536 < _3518;
    assign _3538 = ~ _3537;
    assign _3526 = _3515[62:62];
    assign _3523 = _3517 - _3518;
    assign _3524 = _3520 ? _3523 : _3517;
    assign _3525 = _3524[62:0];
    assign _3527 = { _3525,
                     _3526 };
    assign _3528 = _3527 < _3518;
    assign _3529 = ~ _3528;
    assign _3518 = 64'b0000000000000000000000000000000000000000000000000000001111101001;
    assign _3514 = 64'b0000000000000000000000000000000000000000000000000000001111101000;
    assign _3515 = _3 + _3514;
    assign _3516 = _3515[63:63];
    assign _3517 = { _22185,
                     _3516 };
    assign _3519 = _3517 < _3518;
    assign _3520 = ~ _3519;
    assign _3521 = { _22185,
                     _3520 };
    assign _3522 = _3521[62:0];
    assign _3530 = { _3522,
                     _3529 };
    assign _3531 = _3530[62:0];
    assign _3539 = { _3531,
                     _3538 };
    assign _3540 = _3539[62:0];
    assign _3548 = { _3540,
                     _3547 };
    assign _3549 = _3548[62:0];
    assign _3557 = { _3549,
                     _3556 };
    assign _3558 = _3557[62:0];
    assign _3566 = { _3558,
                     _3565 };
    assign _3567 = _3566[62:0];
    assign _3575 = { _3567,
                     _3574 };
    assign _3576 = _3575[62:0];
    assign _3584 = { _3576,
                     _3583 };
    assign _3585 = _3584[62:0];
    assign _3593 = { _3585,
                     _3592 };
    assign _3594 = _3593[62:0];
    assign _3602 = { _3594,
                     _3601 };
    assign _3603 = _3602[62:0];
    assign _3611 = { _3603,
                     _3610 };
    assign _3612 = _3611[62:0];
    assign _3620 = { _3612,
                     _3619 };
    assign _3621 = _3620[62:0];
    assign _3629 = { _3621,
                     _3628 };
    assign _3630 = _3629[62:0];
    assign _3638 = { _3630,
                     _3637 };
    assign _3639 = _3638[62:0];
    assign _3647 = { _3639,
                     _3646 };
    assign _3648 = _3647[62:0];
    assign _3656 = { _3648,
                     _3655 };
    assign _3657 = _3656[62:0];
    assign _3665 = { _3657,
                     _3664 };
    assign _3666 = _3665[62:0];
    assign _3674 = { _3666,
                     _3673 };
    assign _3675 = _3674[62:0];
    assign _3683 = { _3675,
                     _3682 };
    assign _3684 = _3683[62:0];
    assign _3692 = { _3684,
                     _3691 };
    assign _3693 = _3692[62:0];
    assign _3701 = { _3693,
                     _3700 };
    assign _3702 = _3701[62:0];
    assign _3710 = { _3702,
                     _3709 };
    assign _3711 = _3710[62:0];
    assign _3719 = { _3711,
                     _3718 };
    assign _3720 = _3719[62:0];
    assign _3728 = { _3720,
                     _3727 };
    assign _3729 = _3728[62:0];
    assign _3737 = { _3729,
                     _3736 };
    assign _3738 = _3737[62:0];
    assign _3746 = { _3738,
                     _3745 };
    assign _3747 = _3746[62:0];
    assign _3755 = { _3747,
                     _3754 };
    assign _3756 = _3755[62:0];
    assign _3764 = { _3756,
                     _3763 };
    assign _3765 = _3764[62:0];
    assign _3773 = { _3765,
                     _3772 };
    assign _3774 = _3773[62:0];
    assign _3782 = { _3774,
                     _3781 };
    assign _3783 = _3782[62:0];
    assign _3791 = { _3783,
                     _3790 };
    assign _3792 = _3791[62:0];
    assign _3800 = { _3792,
                     _3799 };
    assign _3801 = _3800[62:0];
    assign _3809 = { _3801,
                     _3808 };
    assign _3810 = _3809[62:0];
    assign _3818 = { _3810,
                     _3817 };
    assign _3819 = _3818[62:0];
    assign _3827 = { _3819,
                     _3826 };
    assign _3828 = _3827[62:0];
    assign _3836 = { _3828,
                     _3835 };
    assign _3837 = _3836[62:0];
    assign _3845 = { _3837,
                     _3844 };
    assign _3846 = _3845[62:0];
    assign _3854 = { _3846,
                     _3853 };
    assign _3855 = _3854[62:0];
    assign _3863 = { _3855,
                     _3862 };
    assign _3864 = _3863[62:0];
    assign _3872 = { _3864,
                     _3871 };
    assign _3873 = _3872[62:0];
    assign _3881 = { _3873,
                     _3880 };
    assign _3882 = _3881[62:0];
    assign _3890 = { _3882,
                     _3889 };
    assign _3891 = _3890[62:0];
    assign _3899 = { _3891,
                     _3898 };
    assign _3900 = _3899[62:0];
    assign _3908 = { _3900,
                     _3907 };
    assign _3909 = _3908[62:0];
    assign _3917 = { _3909,
                     _3916 };
    assign _3918 = _3917[62:0];
    assign _3926 = { _3918,
                     _3925 };
    assign _3927 = _3926[62:0];
    assign _3935 = { _3927,
                     _3934 };
    assign _3936 = _3935[62:0];
    assign _3944 = { _3936,
                     _3943 };
    assign _3945 = _3944[62:0];
    assign _3953 = { _3945,
                     _3952 };
    assign _3954 = _3953[62:0];
    assign _3962 = { _3954,
                     _3961 };
    assign _3963 = _3962[62:0];
    assign _3971 = { _3963,
                     _3970 };
    assign _3972 = _3971[62:0];
    assign _3980 = { _3972,
                     _3979 };
    assign _3981 = _3980[62:0];
    assign _3989 = { _3981,
                     _3988 };
    assign _3990 = _3989[62:0];
    assign _3998 = { _3990,
                     _3997 };
    assign _3999 = _3998[62:0];
    assign _4007 = { _3999,
                     _4006 };
    assign _4008 = _4007[62:0];
    assign _4016 = { _4008,
                     _4015 };
    assign _4017 = _4016[62:0];
    assign _4025 = { _4017,
                     _4024 };
    assign _4026 = _4025[62:0];
    assign _4034 = { _4026,
                     _4033 };
    assign _4035 = _4034[62:0];
    assign _4043 = { _4035,
                     _4042 };
    assign _4044 = _4043[62:0];
    assign _4052 = { _4044,
                     _4051 };
    assign _4053 = _4052[62:0];
    assign _4061 = { _4053,
                     _4060 };
    assign _4062 = _4061[62:0];
    assign _4070 = { _4062,
                     _4069 };
    assign _4071 = _4070[62:0];
    assign _4079 = { _4071,
                     _4078 };
    assign _4080 = _4079[62:0];
    assign _4088 = { _4080,
                     _4087 };
    assign _4089 = _4088 * _3518;
    assign _4090 = _4089[63:0];
    assign _3511 = 64'b0000000000000000000000000000000000000000000000011000011100000100;
    assign _4091 = _3511 < _4090;
    assign _4092 = _4091 ? _4090 : _3511;
    assign _3509 = _5 < _19267;
    assign _3510 = _3509 ? _5 : _19267;
    assign _4093 = _3510 < _4092;
    assign _4094 = ~ _4093;
    assign _5257 = _4094 ? _5256 : _21604;
    assign _3498 = _2929[0:0];
    assign _3495 = _3490 - _22192;
    assign _3496 = _3492 ? _3495 : _3490;
    assign _3497 = _3496[62:0];
    assign _3499 = { _3497,
                     _3498 };
    assign _3500 = _3499 < _22192;
    assign _3501 = ~ _3500;
    assign _3489 = _2929[1:1];
    assign _3486 = _3481 - _22192;
    assign _3487 = _3483 ? _3486 : _3481;
    assign _3488 = _3487[62:0];
    assign _3490 = { _3488,
                     _3489 };
    assign _3491 = _3490 < _22192;
    assign _3492 = ~ _3491;
    assign _3480 = _2929[2:2];
    assign _3477 = _3472 - _22192;
    assign _3478 = _3474 ? _3477 : _3472;
    assign _3479 = _3478[62:0];
    assign _3481 = { _3479,
                     _3480 };
    assign _3482 = _3481 < _22192;
    assign _3483 = ~ _3482;
    assign _3471 = _2929[3:3];
    assign _3468 = _3463 - _22192;
    assign _3469 = _3465 ? _3468 : _3463;
    assign _3470 = _3469[62:0];
    assign _3472 = { _3470,
                     _3471 };
    assign _3473 = _3472 < _22192;
    assign _3474 = ~ _3473;
    assign _3462 = _2929[4:4];
    assign _3459 = _3454 - _22192;
    assign _3460 = _3456 ? _3459 : _3454;
    assign _3461 = _3460[62:0];
    assign _3463 = { _3461,
                     _3462 };
    assign _3464 = _3463 < _22192;
    assign _3465 = ~ _3464;
    assign _3453 = _2929[5:5];
    assign _3450 = _3445 - _22192;
    assign _3451 = _3447 ? _3450 : _3445;
    assign _3452 = _3451[62:0];
    assign _3454 = { _3452,
                     _3453 };
    assign _3455 = _3454 < _22192;
    assign _3456 = ~ _3455;
    assign _3444 = _2929[6:6];
    assign _3441 = _3436 - _22192;
    assign _3442 = _3438 ? _3441 : _3436;
    assign _3443 = _3442[62:0];
    assign _3445 = { _3443,
                     _3444 };
    assign _3446 = _3445 < _22192;
    assign _3447 = ~ _3446;
    assign _3435 = _2929[7:7];
    assign _3432 = _3427 - _22192;
    assign _3433 = _3429 ? _3432 : _3427;
    assign _3434 = _3433[62:0];
    assign _3436 = { _3434,
                     _3435 };
    assign _3437 = _3436 < _22192;
    assign _3438 = ~ _3437;
    assign _3426 = _2929[8:8];
    assign _3423 = _3418 - _22192;
    assign _3424 = _3420 ? _3423 : _3418;
    assign _3425 = _3424[62:0];
    assign _3427 = { _3425,
                     _3426 };
    assign _3428 = _3427 < _22192;
    assign _3429 = ~ _3428;
    assign _3417 = _2929[9:9];
    assign _3414 = _3409 - _22192;
    assign _3415 = _3411 ? _3414 : _3409;
    assign _3416 = _3415[62:0];
    assign _3418 = { _3416,
                     _3417 };
    assign _3419 = _3418 < _22192;
    assign _3420 = ~ _3419;
    assign _3408 = _2929[10:10];
    assign _3405 = _3400 - _22192;
    assign _3406 = _3402 ? _3405 : _3400;
    assign _3407 = _3406[62:0];
    assign _3409 = { _3407,
                     _3408 };
    assign _3410 = _3409 < _22192;
    assign _3411 = ~ _3410;
    assign _3399 = _2929[11:11];
    assign _3396 = _3391 - _22192;
    assign _3397 = _3393 ? _3396 : _3391;
    assign _3398 = _3397[62:0];
    assign _3400 = { _3398,
                     _3399 };
    assign _3401 = _3400 < _22192;
    assign _3402 = ~ _3401;
    assign _3390 = _2929[12:12];
    assign _3387 = _3382 - _22192;
    assign _3388 = _3384 ? _3387 : _3382;
    assign _3389 = _3388[62:0];
    assign _3391 = { _3389,
                     _3390 };
    assign _3392 = _3391 < _22192;
    assign _3393 = ~ _3392;
    assign _3381 = _2929[13:13];
    assign _3378 = _3373 - _22192;
    assign _3379 = _3375 ? _3378 : _3373;
    assign _3380 = _3379[62:0];
    assign _3382 = { _3380,
                     _3381 };
    assign _3383 = _3382 < _22192;
    assign _3384 = ~ _3383;
    assign _3372 = _2929[14:14];
    assign _3369 = _3364 - _22192;
    assign _3370 = _3366 ? _3369 : _3364;
    assign _3371 = _3370[62:0];
    assign _3373 = { _3371,
                     _3372 };
    assign _3374 = _3373 < _22192;
    assign _3375 = ~ _3374;
    assign _3363 = _2929[15:15];
    assign _3360 = _3355 - _22192;
    assign _3361 = _3357 ? _3360 : _3355;
    assign _3362 = _3361[62:0];
    assign _3364 = { _3362,
                     _3363 };
    assign _3365 = _3364 < _22192;
    assign _3366 = ~ _3365;
    assign _3354 = _2929[16:16];
    assign _3351 = _3346 - _22192;
    assign _3352 = _3348 ? _3351 : _3346;
    assign _3353 = _3352[62:0];
    assign _3355 = { _3353,
                     _3354 };
    assign _3356 = _3355 < _22192;
    assign _3357 = ~ _3356;
    assign _3345 = _2929[17:17];
    assign _3342 = _3337 - _22192;
    assign _3343 = _3339 ? _3342 : _3337;
    assign _3344 = _3343[62:0];
    assign _3346 = { _3344,
                     _3345 };
    assign _3347 = _3346 < _22192;
    assign _3348 = ~ _3347;
    assign _3336 = _2929[18:18];
    assign _3333 = _3328 - _22192;
    assign _3334 = _3330 ? _3333 : _3328;
    assign _3335 = _3334[62:0];
    assign _3337 = { _3335,
                     _3336 };
    assign _3338 = _3337 < _22192;
    assign _3339 = ~ _3338;
    assign _3327 = _2929[19:19];
    assign _3324 = _3319 - _22192;
    assign _3325 = _3321 ? _3324 : _3319;
    assign _3326 = _3325[62:0];
    assign _3328 = { _3326,
                     _3327 };
    assign _3329 = _3328 < _22192;
    assign _3330 = ~ _3329;
    assign _3318 = _2929[20:20];
    assign _3315 = _3310 - _22192;
    assign _3316 = _3312 ? _3315 : _3310;
    assign _3317 = _3316[62:0];
    assign _3319 = { _3317,
                     _3318 };
    assign _3320 = _3319 < _22192;
    assign _3321 = ~ _3320;
    assign _3309 = _2929[21:21];
    assign _3306 = _3301 - _22192;
    assign _3307 = _3303 ? _3306 : _3301;
    assign _3308 = _3307[62:0];
    assign _3310 = { _3308,
                     _3309 };
    assign _3311 = _3310 < _22192;
    assign _3312 = ~ _3311;
    assign _3300 = _2929[22:22];
    assign _3297 = _3292 - _22192;
    assign _3298 = _3294 ? _3297 : _3292;
    assign _3299 = _3298[62:0];
    assign _3301 = { _3299,
                     _3300 };
    assign _3302 = _3301 < _22192;
    assign _3303 = ~ _3302;
    assign _3291 = _2929[23:23];
    assign _3288 = _3283 - _22192;
    assign _3289 = _3285 ? _3288 : _3283;
    assign _3290 = _3289[62:0];
    assign _3292 = { _3290,
                     _3291 };
    assign _3293 = _3292 < _22192;
    assign _3294 = ~ _3293;
    assign _3282 = _2929[24:24];
    assign _3279 = _3274 - _22192;
    assign _3280 = _3276 ? _3279 : _3274;
    assign _3281 = _3280[62:0];
    assign _3283 = { _3281,
                     _3282 };
    assign _3284 = _3283 < _22192;
    assign _3285 = ~ _3284;
    assign _3273 = _2929[25:25];
    assign _3270 = _3265 - _22192;
    assign _3271 = _3267 ? _3270 : _3265;
    assign _3272 = _3271[62:0];
    assign _3274 = { _3272,
                     _3273 };
    assign _3275 = _3274 < _22192;
    assign _3276 = ~ _3275;
    assign _3264 = _2929[26:26];
    assign _3261 = _3256 - _22192;
    assign _3262 = _3258 ? _3261 : _3256;
    assign _3263 = _3262[62:0];
    assign _3265 = { _3263,
                     _3264 };
    assign _3266 = _3265 < _22192;
    assign _3267 = ~ _3266;
    assign _3255 = _2929[27:27];
    assign _3252 = _3247 - _22192;
    assign _3253 = _3249 ? _3252 : _3247;
    assign _3254 = _3253[62:0];
    assign _3256 = { _3254,
                     _3255 };
    assign _3257 = _3256 < _22192;
    assign _3258 = ~ _3257;
    assign _3246 = _2929[28:28];
    assign _3243 = _3238 - _22192;
    assign _3244 = _3240 ? _3243 : _3238;
    assign _3245 = _3244[62:0];
    assign _3247 = { _3245,
                     _3246 };
    assign _3248 = _3247 < _22192;
    assign _3249 = ~ _3248;
    assign _3237 = _2929[29:29];
    assign _3234 = _3229 - _22192;
    assign _3235 = _3231 ? _3234 : _3229;
    assign _3236 = _3235[62:0];
    assign _3238 = { _3236,
                     _3237 };
    assign _3239 = _3238 < _22192;
    assign _3240 = ~ _3239;
    assign _3228 = _2929[30:30];
    assign _3225 = _3220 - _22192;
    assign _3226 = _3222 ? _3225 : _3220;
    assign _3227 = _3226[62:0];
    assign _3229 = { _3227,
                     _3228 };
    assign _3230 = _3229 < _22192;
    assign _3231 = ~ _3230;
    assign _3219 = _2929[31:31];
    assign _3216 = _3211 - _22192;
    assign _3217 = _3213 ? _3216 : _3211;
    assign _3218 = _3217[62:0];
    assign _3220 = { _3218,
                     _3219 };
    assign _3221 = _3220 < _22192;
    assign _3222 = ~ _3221;
    assign _3210 = _2929[32:32];
    assign _3207 = _3202 - _22192;
    assign _3208 = _3204 ? _3207 : _3202;
    assign _3209 = _3208[62:0];
    assign _3211 = { _3209,
                     _3210 };
    assign _3212 = _3211 < _22192;
    assign _3213 = ~ _3212;
    assign _3201 = _2929[33:33];
    assign _3198 = _3193 - _22192;
    assign _3199 = _3195 ? _3198 : _3193;
    assign _3200 = _3199[62:0];
    assign _3202 = { _3200,
                     _3201 };
    assign _3203 = _3202 < _22192;
    assign _3204 = ~ _3203;
    assign _3192 = _2929[34:34];
    assign _3189 = _3184 - _22192;
    assign _3190 = _3186 ? _3189 : _3184;
    assign _3191 = _3190[62:0];
    assign _3193 = { _3191,
                     _3192 };
    assign _3194 = _3193 < _22192;
    assign _3195 = ~ _3194;
    assign _3183 = _2929[35:35];
    assign _3180 = _3175 - _22192;
    assign _3181 = _3177 ? _3180 : _3175;
    assign _3182 = _3181[62:0];
    assign _3184 = { _3182,
                     _3183 };
    assign _3185 = _3184 < _22192;
    assign _3186 = ~ _3185;
    assign _3174 = _2929[36:36];
    assign _3171 = _3166 - _22192;
    assign _3172 = _3168 ? _3171 : _3166;
    assign _3173 = _3172[62:0];
    assign _3175 = { _3173,
                     _3174 };
    assign _3176 = _3175 < _22192;
    assign _3177 = ~ _3176;
    assign _3165 = _2929[37:37];
    assign _3162 = _3157 - _22192;
    assign _3163 = _3159 ? _3162 : _3157;
    assign _3164 = _3163[62:0];
    assign _3166 = { _3164,
                     _3165 };
    assign _3167 = _3166 < _22192;
    assign _3168 = ~ _3167;
    assign _3156 = _2929[38:38];
    assign _3153 = _3148 - _22192;
    assign _3154 = _3150 ? _3153 : _3148;
    assign _3155 = _3154[62:0];
    assign _3157 = { _3155,
                     _3156 };
    assign _3158 = _3157 < _22192;
    assign _3159 = ~ _3158;
    assign _3147 = _2929[39:39];
    assign _3144 = _3139 - _22192;
    assign _3145 = _3141 ? _3144 : _3139;
    assign _3146 = _3145[62:0];
    assign _3148 = { _3146,
                     _3147 };
    assign _3149 = _3148 < _22192;
    assign _3150 = ~ _3149;
    assign _3138 = _2929[40:40];
    assign _3135 = _3130 - _22192;
    assign _3136 = _3132 ? _3135 : _3130;
    assign _3137 = _3136[62:0];
    assign _3139 = { _3137,
                     _3138 };
    assign _3140 = _3139 < _22192;
    assign _3141 = ~ _3140;
    assign _3129 = _2929[41:41];
    assign _3126 = _3121 - _22192;
    assign _3127 = _3123 ? _3126 : _3121;
    assign _3128 = _3127[62:0];
    assign _3130 = { _3128,
                     _3129 };
    assign _3131 = _3130 < _22192;
    assign _3132 = ~ _3131;
    assign _3120 = _2929[42:42];
    assign _3117 = _3112 - _22192;
    assign _3118 = _3114 ? _3117 : _3112;
    assign _3119 = _3118[62:0];
    assign _3121 = { _3119,
                     _3120 };
    assign _3122 = _3121 < _22192;
    assign _3123 = ~ _3122;
    assign _3111 = _2929[43:43];
    assign _3108 = _3103 - _22192;
    assign _3109 = _3105 ? _3108 : _3103;
    assign _3110 = _3109[62:0];
    assign _3112 = { _3110,
                     _3111 };
    assign _3113 = _3112 < _22192;
    assign _3114 = ~ _3113;
    assign _3102 = _2929[44:44];
    assign _3099 = _3094 - _22192;
    assign _3100 = _3096 ? _3099 : _3094;
    assign _3101 = _3100[62:0];
    assign _3103 = { _3101,
                     _3102 };
    assign _3104 = _3103 < _22192;
    assign _3105 = ~ _3104;
    assign _3093 = _2929[45:45];
    assign _3090 = _3085 - _22192;
    assign _3091 = _3087 ? _3090 : _3085;
    assign _3092 = _3091[62:0];
    assign _3094 = { _3092,
                     _3093 };
    assign _3095 = _3094 < _22192;
    assign _3096 = ~ _3095;
    assign _3084 = _2929[46:46];
    assign _3081 = _3076 - _22192;
    assign _3082 = _3078 ? _3081 : _3076;
    assign _3083 = _3082[62:0];
    assign _3085 = { _3083,
                     _3084 };
    assign _3086 = _3085 < _22192;
    assign _3087 = ~ _3086;
    assign _3075 = _2929[47:47];
    assign _3072 = _3067 - _22192;
    assign _3073 = _3069 ? _3072 : _3067;
    assign _3074 = _3073[62:0];
    assign _3076 = { _3074,
                     _3075 };
    assign _3077 = _3076 < _22192;
    assign _3078 = ~ _3077;
    assign _3066 = _2929[48:48];
    assign _3063 = _3058 - _22192;
    assign _3064 = _3060 ? _3063 : _3058;
    assign _3065 = _3064[62:0];
    assign _3067 = { _3065,
                     _3066 };
    assign _3068 = _3067 < _22192;
    assign _3069 = ~ _3068;
    assign _3057 = _2929[49:49];
    assign _3054 = _3049 - _22192;
    assign _3055 = _3051 ? _3054 : _3049;
    assign _3056 = _3055[62:0];
    assign _3058 = { _3056,
                     _3057 };
    assign _3059 = _3058 < _22192;
    assign _3060 = ~ _3059;
    assign _3048 = _2929[50:50];
    assign _3045 = _3040 - _22192;
    assign _3046 = _3042 ? _3045 : _3040;
    assign _3047 = _3046[62:0];
    assign _3049 = { _3047,
                     _3048 };
    assign _3050 = _3049 < _22192;
    assign _3051 = ~ _3050;
    assign _3039 = _2929[51:51];
    assign _3036 = _3031 - _22192;
    assign _3037 = _3033 ? _3036 : _3031;
    assign _3038 = _3037[62:0];
    assign _3040 = { _3038,
                     _3039 };
    assign _3041 = _3040 < _22192;
    assign _3042 = ~ _3041;
    assign _3030 = _2929[52:52];
    assign _3027 = _3022 - _22192;
    assign _3028 = _3024 ? _3027 : _3022;
    assign _3029 = _3028[62:0];
    assign _3031 = { _3029,
                     _3030 };
    assign _3032 = _3031 < _22192;
    assign _3033 = ~ _3032;
    assign _3021 = _2929[53:53];
    assign _3018 = _3013 - _22192;
    assign _3019 = _3015 ? _3018 : _3013;
    assign _3020 = _3019[62:0];
    assign _3022 = { _3020,
                     _3021 };
    assign _3023 = _3022 < _22192;
    assign _3024 = ~ _3023;
    assign _3012 = _2929[54:54];
    assign _3009 = _3004 - _22192;
    assign _3010 = _3006 ? _3009 : _3004;
    assign _3011 = _3010[62:0];
    assign _3013 = { _3011,
                     _3012 };
    assign _3014 = _3013 < _22192;
    assign _3015 = ~ _3014;
    assign _3003 = _2929[55:55];
    assign _3000 = _2995 - _22192;
    assign _3001 = _2997 ? _3000 : _2995;
    assign _3002 = _3001[62:0];
    assign _3004 = { _3002,
                     _3003 };
    assign _3005 = _3004 < _22192;
    assign _3006 = ~ _3005;
    assign _2994 = _2929[56:56];
    assign _2991 = _2986 - _22192;
    assign _2992 = _2988 ? _2991 : _2986;
    assign _2993 = _2992[62:0];
    assign _2995 = { _2993,
                     _2994 };
    assign _2996 = _2995 < _22192;
    assign _2997 = ~ _2996;
    assign _2985 = _2929[57:57];
    assign _2982 = _2977 - _22192;
    assign _2983 = _2979 ? _2982 : _2977;
    assign _2984 = _2983[62:0];
    assign _2986 = { _2984,
                     _2985 };
    assign _2987 = _2986 < _22192;
    assign _2988 = ~ _2987;
    assign _2976 = _2929[58:58];
    assign _2973 = _2968 - _22192;
    assign _2974 = _2970 ? _2973 : _2968;
    assign _2975 = _2974[62:0];
    assign _2977 = { _2975,
                     _2976 };
    assign _2978 = _2977 < _22192;
    assign _2979 = ~ _2978;
    assign _2967 = _2929[59:59];
    assign _2964 = _2959 - _22192;
    assign _2965 = _2961 ? _2964 : _2959;
    assign _2966 = _2965[62:0];
    assign _2968 = { _2966,
                     _2967 };
    assign _2969 = _2968 < _22192;
    assign _2970 = ~ _2969;
    assign _2958 = _2929[60:60];
    assign _2955 = _2950 - _22192;
    assign _2956 = _2952 ? _2955 : _2950;
    assign _2957 = _2956[62:0];
    assign _2959 = { _2957,
                     _2958 };
    assign _2960 = _2959 < _22192;
    assign _2961 = ~ _2960;
    assign _2949 = _2929[61:61];
    assign _2946 = _2941 - _22192;
    assign _2947 = _2943 ? _2946 : _2941;
    assign _2948 = _2947[62:0];
    assign _2950 = { _2948,
                     _2949 };
    assign _2951 = _2950 < _22192;
    assign _2952 = ~ _2951;
    assign _2940 = _2929[62:62];
    assign _2937 = _2931 - _22192;
    assign _2938 = _2934 ? _2937 : _2931;
    assign _2939 = _2938[62:0];
    assign _2941 = { _2939,
                     _2940 };
    assign _2942 = _2941 < _22192;
    assign _2943 = ~ _2942;
    assign _2927 = _2919 + _22186;
    assign _2928 = _2919 * _2927;
    assign _2929 = _2928[63:0];
    assign _2930 = _2929[63:63];
    assign _2931 = { _22185,
                     _2930 };
    assign _2933 = _2931 < _22192;
    assign _2934 = ~ _2933;
    assign _2935 = { _22185,
                     _2934 };
    assign _2936 = _2935[62:0];
    assign _2944 = { _2936,
                     _2943 };
    assign _2945 = _2944[62:0];
    assign _2953 = { _2945,
                     _2952 };
    assign _2954 = _2953[62:0];
    assign _2962 = { _2954,
                     _2961 };
    assign _2963 = _2962[62:0];
    assign _2971 = { _2963,
                     _2970 };
    assign _2972 = _2971[62:0];
    assign _2980 = { _2972,
                     _2979 };
    assign _2981 = _2980[62:0];
    assign _2989 = { _2981,
                     _2988 };
    assign _2990 = _2989[62:0];
    assign _2998 = { _2990,
                     _2997 };
    assign _2999 = _2998[62:0];
    assign _3007 = { _2999,
                     _3006 };
    assign _3008 = _3007[62:0];
    assign _3016 = { _3008,
                     _3015 };
    assign _3017 = _3016[62:0];
    assign _3025 = { _3017,
                     _3024 };
    assign _3026 = _3025[62:0];
    assign _3034 = { _3026,
                     _3033 };
    assign _3035 = _3034[62:0];
    assign _3043 = { _3035,
                     _3042 };
    assign _3044 = _3043[62:0];
    assign _3052 = { _3044,
                     _3051 };
    assign _3053 = _3052[62:0];
    assign _3061 = { _3053,
                     _3060 };
    assign _3062 = _3061[62:0];
    assign _3070 = { _3062,
                     _3069 };
    assign _3071 = _3070[62:0];
    assign _3079 = { _3071,
                     _3078 };
    assign _3080 = _3079[62:0];
    assign _3088 = { _3080,
                     _3087 };
    assign _3089 = _3088[62:0];
    assign _3097 = { _3089,
                     _3096 };
    assign _3098 = _3097[62:0];
    assign _3106 = { _3098,
                     _3105 };
    assign _3107 = _3106[62:0];
    assign _3115 = { _3107,
                     _3114 };
    assign _3116 = _3115[62:0];
    assign _3124 = { _3116,
                     _3123 };
    assign _3125 = _3124[62:0];
    assign _3133 = { _3125,
                     _3132 };
    assign _3134 = _3133[62:0];
    assign _3142 = { _3134,
                     _3141 };
    assign _3143 = _3142[62:0];
    assign _3151 = { _3143,
                     _3150 };
    assign _3152 = _3151[62:0];
    assign _3160 = { _3152,
                     _3159 };
    assign _3161 = _3160[62:0];
    assign _3169 = { _3161,
                     _3168 };
    assign _3170 = _3169[62:0];
    assign _3178 = { _3170,
                     _3177 };
    assign _3179 = _3178[62:0];
    assign _3187 = { _3179,
                     _3186 };
    assign _3188 = _3187[62:0];
    assign _3196 = { _3188,
                     _3195 };
    assign _3197 = _3196[62:0];
    assign _3205 = { _3197,
                     _3204 };
    assign _3206 = _3205[62:0];
    assign _3214 = { _3206,
                     _3213 };
    assign _3215 = _3214[62:0];
    assign _3223 = { _3215,
                     _3222 };
    assign _3224 = _3223[62:0];
    assign _3232 = { _3224,
                     _3231 };
    assign _3233 = _3232[62:0];
    assign _3241 = { _3233,
                     _3240 };
    assign _3242 = _3241[62:0];
    assign _3250 = { _3242,
                     _3249 };
    assign _3251 = _3250[62:0];
    assign _3259 = { _3251,
                     _3258 };
    assign _3260 = _3259[62:0];
    assign _3268 = { _3260,
                     _3267 };
    assign _3269 = _3268[62:0];
    assign _3277 = { _3269,
                     _3276 };
    assign _3278 = _3277[62:0];
    assign _3286 = { _3278,
                     _3285 };
    assign _3287 = _3286[62:0];
    assign _3295 = { _3287,
                     _3294 };
    assign _3296 = _3295[62:0];
    assign _3304 = { _3296,
                     _3303 };
    assign _3305 = _3304[62:0];
    assign _3313 = { _3305,
                     _3312 };
    assign _3314 = _3313[62:0];
    assign _3322 = { _3314,
                     _3321 };
    assign _3323 = _3322[62:0];
    assign _3331 = { _3323,
                     _3330 };
    assign _3332 = _3331[62:0];
    assign _3340 = { _3332,
                     _3339 };
    assign _3341 = _3340[62:0];
    assign _3349 = { _3341,
                     _3348 };
    assign _3350 = _3349[62:0];
    assign _3358 = { _3350,
                     _3357 };
    assign _3359 = _3358[62:0];
    assign _3367 = { _3359,
                     _3366 };
    assign _3368 = _3367[62:0];
    assign _3376 = { _3368,
                     _3375 };
    assign _3377 = _3376[62:0];
    assign _3385 = { _3377,
                     _3384 };
    assign _3386 = _3385[62:0];
    assign _3394 = { _3386,
                     _3393 };
    assign _3395 = _3394[62:0];
    assign _3403 = { _3395,
                     _3402 };
    assign _3404 = _3403[62:0];
    assign _3412 = { _3404,
                     _3411 };
    assign _3413 = _3412[62:0];
    assign _3421 = { _3413,
                     _3420 };
    assign _3422 = _3421[62:0];
    assign _3430 = { _3422,
                     _3429 };
    assign _3431 = _3430[62:0];
    assign _3439 = { _3431,
                     _3438 };
    assign _3440 = _3439[62:0];
    assign _3448 = { _3440,
                     _3447 };
    assign _3449 = _3448[62:0];
    assign _3457 = { _3449,
                     _3456 };
    assign _3458 = _3457[62:0];
    assign _3466 = { _3458,
                     _3465 };
    assign _3467 = _3466[62:0];
    assign _3475 = { _3467,
                     _3474 };
    assign _3476 = _3475[62:0];
    assign _3484 = { _3476,
                     _3483 };
    assign _3485 = _3484[62:0];
    assign _3493 = { _3485,
                     _3492 };
    assign _3494 = _3493[62:0];
    assign _3502 = { _3494,
                     _3501 };
    assign _3503 = _1767 * _3502;
    assign _3504 = _3503[63:0];
    assign _2915 = _2347[0:0];
    assign _2912 = _2907 - _1767;
    assign _2913 = _2909 ? _2912 : _2907;
    assign _2914 = _2913[62:0];
    assign _2916 = { _2914,
                     _2915 };
    assign _2917 = _2916 < _1767;
    assign _2918 = ~ _2917;
    assign _2906 = _2347[1:1];
    assign _2903 = _2898 - _1767;
    assign _2904 = _2900 ? _2903 : _2898;
    assign _2905 = _2904[62:0];
    assign _2907 = { _2905,
                     _2906 };
    assign _2908 = _2907 < _1767;
    assign _2909 = ~ _2908;
    assign _2897 = _2347[2:2];
    assign _2894 = _2889 - _1767;
    assign _2895 = _2891 ? _2894 : _2889;
    assign _2896 = _2895[62:0];
    assign _2898 = { _2896,
                     _2897 };
    assign _2899 = _2898 < _1767;
    assign _2900 = ~ _2899;
    assign _2888 = _2347[3:3];
    assign _2885 = _2880 - _1767;
    assign _2886 = _2882 ? _2885 : _2880;
    assign _2887 = _2886[62:0];
    assign _2889 = { _2887,
                     _2888 };
    assign _2890 = _2889 < _1767;
    assign _2891 = ~ _2890;
    assign _2879 = _2347[4:4];
    assign _2876 = _2871 - _1767;
    assign _2877 = _2873 ? _2876 : _2871;
    assign _2878 = _2877[62:0];
    assign _2880 = { _2878,
                     _2879 };
    assign _2881 = _2880 < _1767;
    assign _2882 = ~ _2881;
    assign _2870 = _2347[5:5];
    assign _2867 = _2862 - _1767;
    assign _2868 = _2864 ? _2867 : _2862;
    assign _2869 = _2868[62:0];
    assign _2871 = { _2869,
                     _2870 };
    assign _2872 = _2871 < _1767;
    assign _2873 = ~ _2872;
    assign _2861 = _2347[6:6];
    assign _2858 = _2853 - _1767;
    assign _2859 = _2855 ? _2858 : _2853;
    assign _2860 = _2859[62:0];
    assign _2862 = { _2860,
                     _2861 };
    assign _2863 = _2862 < _1767;
    assign _2864 = ~ _2863;
    assign _2852 = _2347[7:7];
    assign _2849 = _2844 - _1767;
    assign _2850 = _2846 ? _2849 : _2844;
    assign _2851 = _2850[62:0];
    assign _2853 = { _2851,
                     _2852 };
    assign _2854 = _2853 < _1767;
    assign _2855 = ~ _2854;
    assign _2843 = _2347[8:8];
    assign _2840 = _2835 - _1767;
    assign _2841 = _2837 ? _2840 : _2835;
    assign _2842 = _2841[62:0];
    assign _2844 = { _2842,
                     _2843 };
    assign _2845 = _2844 < _1767;
    assign _2846 = ~ _2845;
    assign _2834 = _2347[9:9];
    assign _2831 = _2826 - _1767;
    assign _2832 = _2828 ? _2831 : _2826;
    assign _2833 = _2832[62:0];
    assign _2835 = { _2833,
                     _2834 };
    assign _2836 = _2835 < _1767;
    assign _2837 = ~ _2836;
    assign _2825 = _2347[10:10];
    assign _2822 = _2817 - _1767;
    assign _2823 = _2819 ? _2822 : _2817;
    assign _2824 = _2823[62:0];
    assign _2826 = { _2824,
                     _2825 };
    assign _2827 = _2826 < _1767;
    assign _2828 = ~ _2827;
    assign _2816 = _2347[11:11];
    assign _2813 = _2808 - _1767;
    assign _2814 = _2810 ? _2813 : _2808;
    assign _2815 = _2814[62:0];
    assign _2817 = { _2815,
                     _2816 };
    assign _2818 = _2817 < _1767;
    assign _2819 = ~ _2818;
    assign _2807 = _2347[12:12];
    assign _2804 = _2799 - _1767;
    assign _2805 = _2801 ? _2804 : _2799;
    assign _2806 = _2805[62:0];
    assign _2808 = { _2806,
                     _2807 };
    assign _2809 = _2808 < _1767;
    assign _2810 = ~ _2809;
    assign _2798 = _2347[13:13];
    assign _2795 = _2790 - _1767;
    assign _2796 = _2792 ? _2795 : _2790;
    assign _2797 = _2796[62:0];
    assign _2799 = { _2797,
                     _2798 };
    assign _2800 = _2799 < _1767;
    assign _2801 = ~ _2800;
    assign _2789 = _2347[14:14];
    assign _2786 = _2781 - _1767;
    assign _2787 = _2783 ? _2786 : _2781;
    assign _2788 = _2787[62:0];
    assign _2790 = { _2788,
                     _2789 };
    assign _2791 = _2790 < _1767;
    assign _2792 = ~ _2791;
    assign _2780 = _2347[15:15];
    assign _2777 = _2772 - _1767;
    assign _2778 = _2774 ? _2777 : _2772;
    assign _2779 = _2778[62:0];
    assign _2781 = { _2779,
                     _2780 };
    assign _2782 = _2781 < _1767;
    assign _2783 = ~ _2782;
    assign _2771 = _2347[16:16];
    assign _2768 = _2763 - _1767;
    assign _2769 = _2765 ? _2768 : _2763;
    assign _2770 = _2769[62:0];
    assign _2772 = { _2770,
                     _2771 };
    assign _2773 = _2772 < _1767;
    assign _2774 = ~ _2773;
    assign _2762 = _2347[17:17];
    assign _2759 = _2754 - _1767;
    assign _2760 = _2756 ? _2759 : _2754;
    assign _2761 = _2760[62:0];
    assign _2763 = { _2761,
                     _2762 };
    assign _2764 = _2763 < _1767;
    assign _2765 = ~ _2764;
    assign _2753 = _2347[18:18];
    assign _2750 = _2745 - _1767;
    assign _2751 = _2747 ? _2750 : _2745;
    assign _2752 = _2751[62:0];
    assign _2754 = { _2752,
                     _2753 };
    assign _2755 = _2754 < _1767;
    assign _2756 = ~ _2755;
    assign _2744 = _2347[19:19];
    assign _2741 = _2736 - _1767;
    assign _2742 = _2738 ? _2741 : _2736;
    assign _2743 = _2742[62:0];
    assign _2745 = { _2743,
                     _2744 };
    assign _2746 = _2745 < _1767;
    assign _2747 = ~ _2746;
    assign _2735 = _2347[20:20];
    assign _2732 = _2727 - _1767;
    assign _2733 = _2729 ? _2732 : _2727;
    assign _2734 = _2733[62:0];
    assign _2736 = { _2734,
                     _2735 };
    assign _2737 = _2736 < _1767;
    assign _2738 = ~ _2737;
    assign _2726 = _2347[21:21];
    assign _2723 = _2718 - _1767;
    assign _2724 = _2720 ? _2723 : _2718;
    assign _2725 = _2724[62:0];
    assign _2727 = { _2725,
                     _2726 };
    assign _2728 = _2727 < _1767;
    assign _2729 = ~ _2728;
    assign _2717 = _2347[22:22];
    assign _2714 = _2709 - _1767;
    assign _2715 = _2711 ? _2714 : _2709;
    assign _2716 = _2715[62:0];
    assign _2718 = { _2716,
                     _2717 };
    assign _2719 = _2718 < _1767;
    assign _2720 = ~ _2719;
    assign _2708 = _2347[23:23];
    assign _2705 = _2700 - _1767;
    assign _2706 = _2702 ? _2705 : _2700;
    assign _2707 = _2706[62:0];
    assign _2709 = { _2707,
                     _2708 };
    assign _2710 = _2709 < _1767;
    assign _2711 = ~ _2710;
    assign _2699 = _2347[24:24];
    assign _2696 = _2691 - _1767;
    assign _2697 = _2693 ? _2696 : _2691;
    assign _2698 = _2697[62:0];
    assign _2700 = { _2698,
                     _2699 };
    assign _2701 = _2700 < _1767;
    assign _2702 = ~ _2701;
    assign _2690 = _2347[25:25];
    assign _2687 = _2682 - _1767;
    assign _2688 = _2684 ? _2687 : _2682;
    assign _2689 = _2688[62:0];
    assign _2691 = { _2689,
                     _2690 };
    assign _2692 = _2691 < _1767;
    assign _2693 = ~ _2692;
    assign _2681 = _2347[26:26];
    assign _2678 = _2673 - _1767;
    assign _2679 = _2675 ? _2678 : _2673;
    assign _2680 = _2679[62:0];
    assign _2682 = { _2680,
                     _2681 };
    assign _2683 = _2682 < _1767;
    assign _2684 = ~ _2683;
    assign _2672 = _2347[27:27];
    assign _2669 = _2664 - _1767;
    assign _2670 = _2666 ? _2669 : _2664;
    assign _2671 = _2670[62:0];
    assign _2673 = { _2671,
                     _2672 };
    assign _2674 = _2673 < _1767;
    assign _2675 = ~ _2674;
    assign _2663 = _2347[28:28];
    assign _2660 = _2655 - _1767;
    assign _2661 = _2657 ? _2660 : _2655;
    assign _2662 = _2661[62:0];
    assign _2664 = { _2662,
                     _2663 };
    assign _2665 = _2664 < _1767;
    assign _2666 = ~ _2665;
    assign _2654 = _2347[29:29];
    assign _2651 = _2646 - _1767;
    assign _2652 = _2648 ? _2651 : _2646;
    assign _2653 = _2652[62:0];
    assign _2655 = { _2653,
                     _2654 };
    assign _2656 = _2655 < _1767;
    assign _2657 = ~ _2656;
    assign _2645 = _2347[30:30];
    assign _2642 = _2637 - _1767;
    assign _2643 = _2639 ? _2642 : _2637;
    assign _2644 = _2643[62:0];
    assign _2646 = { _2644,
                     _2645 };
    assign _2647 = _2646 < _1767;
    assign _2648 = ~ _2647;
    assign _2636 = _2347[31:31];
    assign _2633 = _2628 - _1767;
    assign _2634 = _2630 ? _2633 : _2628;
    assign _2635 = _2634[62:0];
    assign _2637 = { _2635,
                     _2636 };
    assign _2638 = _2637 < _1767;
    assign _2639 = ~ _2638;
    assign _2627 = _2347[32:32];
    assign _2624 = _2619 - _1767;
    assign _2625 = _2621 ? _2624 : _2619;
    assign _2626 = _2625[62:0];
    assign _2628 = { _2626,
                     _2627 };
    assign _2629 = _2628 < _1767;
    assign _2630 = ~ _2629;
    assign _2618 = _2347[33:33];
    assign _2615 = _2610 - _1767;
    assign _2616 = _2612 ? _2615 : _2610;
    assign _2617 = _2616[62:0];
    assign _2619 = { _2617,
                     _2618 };
    assign _2620 = _2619 < _1767;
    assign _2621 = ~ _2620;
    assign _2609 = _2347[34:34];
    assign _2606 = _2601 - _1767;
    assign _2607 = _2603 ? _2606 : _2601;
    assign _2608 = _2607[62:0];
    assign _2610 = { _2608,
                     _2609 };
    assign _2611 = _2610 < _1767;
    assign _2612 = ~ _2611;
    assign _2600 = _2347[35:35];
    assign _2597 = _2592 - _1767;
    assign _2598 = _2594 ? _2597 : _2592;
    assign _2599 = _2598[62:0];
    assign _2601 = { _2599,
                     _2600 };
    assign _2602 = _2601 < _1767;
    assign _2603 = ~ _2602;
    assign _2591 = _2347[36:36];
    assign _2588 = _2583 - _1767;
    assign _2589 = _2585 ? _2588 : _2583;
    assign _2590 = _2589[62:0];
    assign _2592 = { _2590,
                     _2591 };
    assign _2593 = _2592 < _1767;
    assign _2594 = ~ _2593;
    assign _2582 = _2347[37:37];
    assign _2579 = _2574 - _1767;
    assign _2580 = _2576 ? _2579 : _2574;
    assign _2581 = _2580[62:0];
    assign _2583 = { _2581,
                     _2582 };
    assign _2584 = _2583 < _1767;
    assign _2585 = ~ _2584;
    assign _2573 = _2347[38:38];
    assign _2570 = _2565 - _1767;
    assign _2571 = _2567 ? _2570 : _2565;
    assign _2572 = _2571[62:0];
    assign _2574 = { _2572,
                     _2573 };
    assign _2575 = _2574 < _1767;
    assign _2576 = ~ _2575;
    assign _2564 = _2347[39:39];
    assign _2561 = _2556 - _1767;
    assign _2562 = _2558 ? _2561 : _2556;
    assign _2563 = _2562[62:0];
    assign _2565 = { _2563,
                     _2564 };
    assign _2566 = _2565 < _1767;
    assign _2567 = ~ _2566;
    assign _2555 = _2347[40:40];
    assign _2552 = _2547 - _1767;
    assign _2553 = _2549 ? _2552 : _2547;
    assign _2554 = _2553[62:0];
    assign _2556 = { _2554,
                     _2555 };
    assign _2557 = _2556 < _1767;
    assign _2558 = ~ _2557;
    assign _2546 = _2347[41:41];
    assign _2543 = _2538 - _1767;
    assign _2544 = _2540 ? _2543 : _2538;
    assign _2545 = _2544[62:0];
    assign _2547 = { _2545,
                     _2546 };
    assign _2548 = _2547 < _1767;
    assign _2549 = ~ _2548;
    assign _2537 = _2347[42:42];
    assign _2534 = _2529 - _1767;
    assign _2535 = _2531 ? _2534 : _2529;
    assign _2536 = _2535[62:0];
    assign _2538 = { _2536,
                     _2537 };
    assign _2539 = _2538 < _1767;
    assign _2540 = ~ _2539;
    assign _2528 = _2347[43:43];
    assign _2525 = _2520 - _1767;
    assign _2526 = _2522 ? _2525 : _2520;
    assign _2527 = _2526[62:0];
    assign _2529 = { _2527,
                     _2528 };
    assign _2530 = _2529 < _1767;
    assign _2531 = ~ _2530;
    assign _2519 = _2347[44:44];
    assign _2516 = _2511 - _1767;
    assign _2517 = _2513 ? _2516 : _2511;
    assign _2518 = _2517[62:0];
    assign _2520 = { _2518,
                     _2519 };
    assign _2521 = _2520 < _1767;
    assign _2522 = ~ _2521;
    assign _2510 = _2347[45:45];
    assign _2507 = _2502 - _1767;
    assign _2508 = _2504 ? _2507 : _2502;
    assign _2509 = _2508[62:0];
    assign _2511 = { _2509,
                     _2510 };
    assign _2512 = _2511 < _1767;
    assign _2513 = ~ _2512;
    assign _2501 = _2347[46:46];
    assign _2498 = _2493 - _1767;
    assign _2499 = _2495 ? _2498 : _2493;
    assign _2500 = _2499[62:0];
    assign _2502 = { _2500,
                     _2501 };
    assign _2503 = _2502 < _1767;
    assign _2504 = ~ _2503;
    assign _2492 = _2347[47:47];
    assign _2489 = _2484 - _1767;
    assign _2490 = _2486 ? _2489 : _2484;
    assign _2491 = _2490[62:0];
    assign _2493 = { _2491,
                     _2492 };
    assign _2494 = _2493 < _1767;
    assign _2495 = ~ _2494;
    assign _2483 = _2347[48:48];
    assign _2480 = _2475 - _1767;
    assign _2481 = _2477 ? _2480 : _2475;
    assign _2482 = _2481[62:0];
    assign _2484 = { _2482,
                     _2483 };
    assign _2485 = _2484 < _1767;
    assign _2486 = ~ _2485;
    assign _2474 = _2347[49:49];
    assign _2471 = _2466 - _1767;
    assign _2472 = _2468 ? _2471 : _2466;
    assign _2473 = _2472[62:0];
    assign _2475 = { _2473,
                     _2474 };
    assign _2476 = _2475 < _1767;
    assign _2477 = ~ _2476;
    assign _2465 = _2347[50:50];
    assign _2462 = _2457 - _1767;
    assign _2463 = _2459 ? _2462 : _2457;
    assign _2464 = _2463[62:0];
    assign _2466 = { _2464,
                     _2465 };
    assign _2467 = _2466 < _1767;
    assign _2468 = ~ _2467;
    assign _2456 = _2347[51:51];
    assign _2453 = _2448 - _1767;
    assign _2454 = _2450 ? _2453 : _2448;
    assign _2455 = _2454[62:0];
    assign _2457 = { _2455,
                     _2456 };
    assign _2458 = _2457 < _1767;
    assign _2459 = ~ _2458;
    assign _2447 = _2347[52:52];
    assign _2444 = _2439 - _1767;
    assign _2445 = _2441 ? _2444 : _2439;
    assign _2446 = _2445[62:0];
    assign _2448 = { _2446,
                     _2447 };
    assign _2449 = _2448 < _1767;
    assign _2450 = ~ _2449;
    assign _2438 = _2347[53:53];
    assign _2435 = _2430 - _1767;
    assign _2436 = _2432 ? _2435 : _2430;
    assign _2437 = _2436[62:0];
    assign _2439 = { _2437,
                     _2438 };
    assign _2440 = _2439 < _1767;
    assign _2441 = ~ _2440;
    assign _2429 = _2347[54:54];
    assign _2426 = _2421 - _1767;
    assign _2427 = _2423 ? _2426 : _2421;
    assign _2428 = _2427[62:0];
    assign _2430 = { _2428,
                     _2429 };
    assign _2431 = _2430 < _1767;
    assign _2432 = ~ _2431;
    assign _2420 = _2347[55:55];
    assign _2417 = _2412 - _1767;
    assign _2418 = _2414 ? _2417 : _2412;
    assign _2419 = _2418[62:0];
    assign _2421 = { _2419,
                     _2420 };
    assign _2422 = _2421 < _1767;
    assign _2423 = ~ _2422;
    assign _2411 = _2347[56:56];
    assign _2408 = _2403 - _1767;
    assign _2409 = _2405 ? _2408 : _2403;
    assign _2410 = _2409[62:0];
    assign _2412 = { _2410,
                     _2411 };
    assign _2413 = _2412 < _1767;
    assign _2414 = ~ _2413;
    assign _2402 = _2347[57:57];
    assign _2399 = _2394 - _1767;
    assign _2400 = _2396 ? _2399 : _2394;
    assign _2401 = _2400[62:0];
    assign _2403 = { _2401,
                     _2402 };
    assign _2404 = _2403 < _1767;
    assign _2405 = ~ _2404;
    assign _2393 = _2347[58:58];
    assign _2390 = _2385 - _1767;
    assign _2391 = _2387 ? _2390 : _2385;
    assign _2392 = _2391[62:0];
    assign _2394 = { _2392,
                     _2393 };
    assign _2395 = _2394 < _1767;
    assign _2396 = ~ _2395;
    assign _2384 = _2347[59:59];
    assign _2381 = _2376 - _1767;
    assign _2382 = _2378 ? _2381 : _2376;
    assign _2383 = _2382[62:0];
    assign _2385 = { _2383,
                     _2384 };
    assign _2386 = _2385 < _1767;
    assign _2387 = ~ _2386;
    assign _2375 = _2347[60:60];
    assign _2372 = _2367 - _1767;
    assign _2373 = _2369 ? _2372 : _2367;
    assign _2374 = _2373[62:0];
    assign _2376 = { _2374,
                     _2375 };
    assign _2377 = _2376 < _1767;
    assign _2378 = ~ _2377;
    assign _2366 = _2347[61:61];
    assign _2363 = _2358 - _1767;
    assign _2364 = _2360 ? _2363 : _2358;
    assign _2365 = _2364[62:0];
    assign _2367 = { _2365,
                     _2366 };
    assign _2368 = _2367 < _1767;
    assign _2369 = ~ _2368;
    assign _2357 = _2347[62:62];
    assign _2354 = _2349 - _1767;
    assign _2355 = _2351 ? _2354 : _2349;
    assign _2356 = _2355[62:0];
    assign _2358 = { _2356,
                     _2357 };
    assign _2359 = _2358 < _1767;
    assign _2360 = ~ _2359;
    assign _2347 = _1759 - _2341;
    assign _2348 = _2347[63:63];
    assign _2349 = { _22185,
                     _2348 };
    assign _2350 = _2349 < _1767;
    assign _2351 = ~ _2350;
    assign _2352 = { _22185,
                     _2351 };
    assign _2353 = _2352[62:0];
    assign _2361 = { _2353,
                     _2360 };
    assign _2362 = _2361[62:0];
    assign _2370 = { _2362,
                     _2369 };
    assign _2371 = _2370[62:0];
    assign _2379 = { _2371,
                     _2378 };
    assign _2380 = _2379[62:0];
    assign _2388 = { _2380,
                     _2387 };
    assign _2389 = _2388[62:0];
    assign _2397 = { _2389,
                     _2396 };
    assign _2398 = _2397[62:0];
    assign _2406 = { _2398,
                     _2405 };
    assign _2407 = _2406[62:0];
    assign _2415 = { _2407,
                     _2414 };
    assign _2416 = _2415[62:0];
    assign _2424 = { _2416,
                     _2423 };
    assign _2425 = _2424[62:0];
    assign _2433 = { _2425,
                     _2432 };
    assign _2434 = _2433[62:0];
    assign _2442 = { _2434,
                     _2441 };
    assign _2443 = _2442[62:0];
    assign _2451 = { _2443,
                     _2450 };
    assign _2452 = _2451[62:0];
    assign _2460 = { _2452,
                     _2459 };
    assign _2461 = _2460[62:0];
    assign _2469 = { _2461,
                     _2468 };
    assign _2470 = _2469[62:0];
    assign _2478 = { _2470,
                     _2477 };
    assign _2479 = _2478[62:0];
    assign _2487 = { _2479,
                     _2486 };
    assign _2488 = _2487[62:0];
    assign _2496 = { _2488,
                     _2495 };
    assign _2497 = _2496[62:0];
    assign _2505 = { _2497,
                     _2504 };
    assign _2506 = _2505[62:0];
    assign _2514 = { _2506,
                     _2513 };
    assign _2515 = _2514[62:0];
    assign _2523 = { _2515,
                     _2522 };
    assign _2524 = _2523[62:0];
    assign _2532 = { _2524,
                     _2531 };
    assign _2533 = _2532[62:0];
    assign _2541 = { _2533,
                     _2540 };
    assign _2542 = _2541[62:0];
    assign _2550 = { _2542,
                     _2549 };
    assign _2551 = _2550[62:0];
    assign _2559 = { _2551,
                     _2558 };
    assign _2560 = _2559[62:0];
    assign _2568 = { _2560,
                     _2567 };
    assign _2569 = _2568[62:0];
    assign _2577 = { _2569,
                     _2576 };
    assign _2578 = _2577[62:0];
    assign _2586 = { _2578,
                     _2585 };
    assign _2587 = _2586[62:0];
    assign _2595 = { _2587,
                     _2594 };
    assign _2596 = _2595[62:0];
    assign _2604 = { _2596,
                     _2603 };
    assign _2605 = _2604[62:0];
    assign _2613 = { _2605,
                     _2612 };
    assign _2614 = _2613[62:0];
    assign _2622 = { _2614,
                     _2621 };
    assign _2623 = _2622[62:0];
    assign _2631 = { _2623,
                     _2630 };
    assign _2632 = _2631[62:0];
    assign _2640 = { _2632,
                     _2639 };
    assign _2641 = _2640[62:0];
    assign _2649 = { _2641,
                     _2648 };
    assign _2650 = _2649[62:0];
    assign _2658 = { _2650,
                     _2657 };
    assign _2659 = _2658[62:0];
    assign _2667 = { _2659,
                     _2666 };
    assign _2668 = _2667[62:0];
    assign _2676 = { _2668,
                     _2675 };
    assign _2677 = _2676[62:0];
    assign _2685 = { _2677,
                     _2684 };
    assign _2686 = _2685[62:0];
    assign _2694 = { _2686,
                     _2693 };
    assign _2695 = _2694[62:0];
    assign _2703 = { _2695,
                     _2702 };
    assign _2704 = _2703[62:0];
    assign _2712 = { _2704,
                     _2711 };
    assign _2713 = _2712[62:0];
    assign _2721 = { _2713,
                     _2720 };
    assign _2722 = _2721[62:0];
    assign _2730 = { _2722,
                     _2729 };
    assign _2731 = _2730[62:0];
    assign _2739 = { _2731,
                     _2738 };
    assign _2740 = _2739[62:0];
    assign _2748 = { _2740,
                     _2747 };
    assign _2749 = _2748[62:0];
    assign _2757 = { _2749,
                     _2756 };
    assign _2758 = _2757[62:0];
    assign _2766 = { _2758,
                     _2765 };
    assign _2767 = _2766[62:0];
    assign _2775 = { _2767,
                     _2774 };
    assign _2776 = _2775[62:0];
    assign _2784 = { _2776,
                     _2783 };
    assign _2785 = _2784[62:0];
    assign _2793 = { _2785,
                     _2792 };
    assign _2794 = _2793[62:0];
    assign _2802 = { _2794,
                     _2801 };
    assign _2803 = _2802[62:0];
    assign _2811 = { _2803,
                     _2810 };
    assign _2812 = _2811[62:0];
    assign _2820 = { _2812,
                     _2819 };
    assign _2821 = _2820[62:0];
    assign _2829 = { _2821,
                     _2828 };
    assign _2830 = _2829[62:0];
    assign _2838 = { _2830,
                     _2837 };
    assign _2839 = _2838[62:0];
    assign _2847 = { _2839,
                     _2846 };
    assign _2848 = _2847[62:0];
    assign _2856 = { _2848,
                     _2855 };
    assign _2857 = _2856[62:0];
    assign _2865 = { _2857,
                     _2864 };
    assign _2866 = _2865[62:0];
    assign _2874 = { _2866,
                     _2873 };
    assign _2875 = _2874[62:0];
    assign _2883 = { _2875,
                     _2882 };
    assign _2884 = _2883[62:0];
    assign _2892 = { _2884,
                     _2891 };
    assign _2893 = _2892[62:0];
    assign _2901 = { _2893,
                     _2900 };
    assign _2902 = _2901[62:0];
    assign _2910 = { _2902,
                     _2909 };
    assign _2911 = _2910[62:0];
    assign _2919 = { _2911,
                     _2918 };
    assign _2921 = _2919 + _22186;
    assign _2922 = _2921 * _2341;
    assign _2923 = _2922[63:0];
    assign _3505 = _2923 + _3504;
    assign _2333 = _1764[0:0];
    assign _2330 = _2325 - _1767;
    assign _2331 = _2327 ? _2330 : _2325;
    assign _2332 = _2331[62:0];
    assign _2334 = { _2332,
                     _2333 };
    assign _2335 = _2334 < _1767;
    assign _2336 = ~ _2335;
    assign _2324 = _1764[1:1];
    assign _2321 = _2316 - _1767;
    assign _2322 = _2318 ? _2321 : _2316;
    assign _2323 = _2322[62:0];
    assign _2325 = { _2323,
                     _2324 };
    assign _2326 = _2325 < _1767;
    assign _2327 = ~ _2326;
    assign _2315 = _1764[2:2];
    assign _2312 = _2307 - _1767;
    assign _2313 = _2309 ? _2312 : _2307;
    assign _2314 = _2313[62:0];
    assign _2316 = { _2314,
                     _2315 };
    assign _2317 = _2316 < _1767;
    assign _2318 = ~ _2317;
    assign _2306 = _1764[3:3];
    assign _2303 = _2298 - _1767;
    assign _2304 = _2300 ? _2303 : _2298;
    assign _2305 = _2304[62:0];
    assign _2307 = { _2305,
                     _2306 };
    assign _2308 = _2307 < _1767;
    assign _2309 = ~ _2308;
    assign _2297 = _1764[4:4];
    assign _2294 = _2289 - _1767;
    assign _2295 = _2291 ? _2294 : _2289;
    assign _2296 = _2295[62:0];
    assign _2298 = { _2296,
                     _2297 };
    assign _2299 = _2298 < _1767;
    assign _2300 = ~ _2299;
    assign _2288 = _1764[5:5];
    assign _2285 = _2280 - _1767;
    assign _2286 = _2282 ? _2285 : _2280;
    assign _2287 = _2286[62:0];
    assign _2289 = { _2287,
                     _2288 };
    assign _2290 = _2289 < _1767;
    assign _2291 = ~ _2290;
    assign _2279 = _1764[6:6];
    assign _2276 = _2271 - _1767;
    assign _2277 = _2273 ? _2276 : _2271;
    assign _2278 = _2277[62:0];
    assign _2280 = { _2278,
                     _2279 };
    assign _2281 = _2280 < _1767;
    assign _2282 = ~ _2281;
    assign _2270 = _1764[7:7];
    assign _2267 = _2262 - _1767;
    assign _2268 = _2264 ? _2267 : _2262;
    assign _2269 = _2268[62:0];
    assign _2271 = { _2269,
                     _2270 };
    assign _2272 = _2271 < _1767;
    assign _2273 = ~ _2272;
    assign _2261 = _1764[8:8];
    assign _2258 = _2253 - _1767;
    assign _2259 = _2255 ? _2258 : _2253;
    assign _2260 = _2259[62:0];
    assign _2262 = { _2260,
                     _2261 };
    assign _2263 = _2262 < _1767;
    assign _2264 = ~ _2263;
    assign _2252 = _1764[9:9];
    assign _2249 = _2244 - _1767;
    assign _2250 = _2246 ? _2249 : _2244;
    assign _2251 = _2250[62:0];
    assign _2253 = { _2251,
                     _2252 };
    assign _2254 = _2253 < _1767;
    assign _2255 = ~ _2254;
    assign _2243 = _1764[10:10];
    assign _2240 = _2235 - _1767;
    assign _2241 = _2237 ? _2240 : _2235;
    assign _2242 = _2241[62:0];
    assign _2244 = { _2242,
                     _2243 };
    assign _2245 = _2244 < _1767;
    assign _2246 = ~ _2245;
    assign _2234 = _1764[11:11];
    assign _2231 = _2226 - _1767;
    assign _2232 = _2228 ? _2231 : _2226;
    assign _2233 = _2232[62:0];
    assign _2235 = { _2233,
                     _2234 };
    assign _2236 = _2235 < _1767;
    assign _2237 = ~ _2236;
    assign _2225 = _1764[12:12];
    assign _2222 = _2217 - _1767;
    assign _2223 = _2219 ? _2222 : _2217;
    assign _2224 = _2223[62:0];
    assign _2226 = { _2224,
                     _2225 };
    assign _2227 = _2226 < _1767;
    assign _2228 = ~ _2227;
    assign _2216 = _1764[13:13];
    assign _2213 = _2208 - _1767;
    assign _2214 = _2210 ? _2213 : _2208;
    assign _2215 = _2214[62:0];
    assign _2217 = { _2215,
                     _2216 };
    assign _2218 = _2217 < _1767;
    assign _2219 = ~ _2218;
    assign _2207 = _1764[14:14];
    assign _2204 = _2199 - _1767;
    assign _2205 = _2201 ? _2204 : _2199;
    assign _2206 = _2205[62:0];
    assign _2208 = { _2206,
                     _2207 };
    assign _2209 = _2208 < _1767;
    assign _2210 = ~ _2209;
    assign _2198 = _1764[15:15];
    assign _2195 = _2190 - _1767;
    assign _2196 = _2192 ? _2195 : _2190;
    assign _2197 = _2196[62:0];
    assign _2199 = { _2197,
                     _2198 };
    assign _2200 = _2199 < _1767;
    assign _2201 = ~ _2200;
    assign _2189 = _1764[16:16];
    assign _2186 = _2181 - _1767;
    assign _2187 = _2183 ? _2186 : _2181;
    assign _2188 = _2187[62:0];
    assign _2190 = { _2188,
                     _2189 };
    assign _2191 = _2190 < _1767;
    assign _2192 = ~ _2191;
    assign _2180 = _1764[17:17];
    assign _2177 = _2172 - _1767;
    assign _2178 = _2174 ? _2177 : _2172;
    assign _2179 = _2178[62:0];
    assign _2181 = { _2179,
                     _2180 };
    assign _2182 = _2181 < _1767;
    assign _2183 = ~ _2182;
    assign _2171 = _1764[18:18];
    assign _2168 = _2163 - _1767;
    assign _2169 = _2165 ? _2168 : _2163;
    assign _2170 = _2169[62:0];
    assign _2172 = { _2170,
                     _2171 };
    assign _2173 = _2172 < _1767;
    assign _2174 = ~ _2173;
    assign _2162 = _1764[19:19];
    assign _2159 = _2154 - _1767;
    assign _2160 = _2156 ? _2159 : _2154;
    assign _2161 = _2160[62:0];
    assign _2163 = { _2161,
                     _2162 };
    assign _2164 = _2163 < _1767;
    assign _2165 = ~ _2164;
    assign _2153 = _1764[20:20];
    assign _2150 = _2145 - _1767;
    assign _2151 = _2147 ? _2150 : _2145;
    assign _2152 = _2151[62:0];
    assign _2154 = { _2152,
                     _2153 };
    assign _2155 = _2154 < _1767;
    assign _2156 = ~ _2155;
    assign _2144 = _1764[21:21];
    assign _2141 = _2136 - _1767;
    assign _2142 = _2138 ? _2141 : _2136;
    assign _2143 = _2142[62:0];
    assign _2145 = { _2143,
                     _2144 };
    assign _2146 = _2145 < _1767;
    assign _2147 = ~ _2146;
    assign _2135 = _1764[22:22];
    assign _2132 = _2127 - _1767;
    assign _2133 = _2129 ? _2132 : _2127;
    assign _2134 = _2133[62:0];
    assign _2136 = { _2134,
                     _2135 };
    assign _2137 = _2136 < _1767;
    assign _2138 = ~ _2137;
    assign _2126 = _1764[23:23];
    assign _2123 = _2118 - _1767;
    assign _2124 = _2120 ? _2123 : _2118;
    assign _2125 = _2124[62:0];
    assign _2127 = { _2125,
                     _2126 };
    assign _2128 = _2127 < _1767;
    assign _2129 = ~ _2128;
    assign _2117 = _1764[24:24];
    assign _2114 = _2109 - _1767;
    assign _2115 = _2111 ? _2114 : _2109;
    assign _2116 = _2115[62:0];
    assign _2118 = { _2116,
                     _2117 };
    assign _2119 = _2118 < _1767;
    assign _2120 = ~ _2119;
    assign _2108 = _1764[25:25];
    assign _2105 = _2100 - _1767;
    assign _2106 = _2102 ? _2105 : _2100;
    assign _2107 = _2106[62:0];
    assign _2109 = { _2107,
                     _2108 };
    assign _2110 = _2109 < _1767;
    assign _2111 = ~ _2110;
    assign _2099 = _1764[26:26];
    assign _2096 = _2091 - _1767;
    assign _2097 = _2093 ? _2096 : _2091;
    assign _2098 = _2097[62:0];
    assign _2100 = { _2098,
                     _2099 };
    assign _2101 = _2100 < _1767;
    assign _2102 = ~ _2101;
    assign _2090 = _1764[27:27];
    assign _2087 = _2082 - _1767;
    assign _2088 = _2084 ? _2087 : _2082;
    assign _2089 = _2088[62:0];
    assign _2091 = { _2089,
                     _2090 };
    assign _2092 = _2091 < _1767;
    assign _2093 = ~ _2092;
    assign _2081 = _1764[28:28];
    assign _2078 = _2073 - _1767;
    assign _2079 = _2075 ? _2078 : _2073;
    assign _2080 = _2079[62:0];
    assign _2082 = { _2080,
                     _2081 };
    assign _2083 = _2082 < _1767;
    assign _2084 = ~ _2083;
    assign _2072 = _1764[29:29];
    assign _2069 = _2064 - _1767;
    assign _2070 = _2066 ? _2069 : _2064;
    assign _2071 = _2070[62:0];
    assign _2073 = { _2071,
                     _2072 };
    assign _2074 = _2073 < _1767;
    assign _2075 = ~ _2074;
    assign _2063 = _1764[30:30];
    assign _2060 = _2055 - _1767;
    assign _2061 = _2057 ? _2060 : _2055;
    assign _2062 = _2061[62:0];
    assign _2064 = { _2062,
                     _2063 };
    assign _2065 = _2064 < _1767;
    assign _2066 = ~ _2065;
    assign _2054 = _1764[31:31];
    assign _2051 = _2046 - _1767;
    assign _2052 = _2048 ? _2051 : _2046;
    assign _2053 = _2052[62:0];
    assign _2055 = { _2053,
                     _2054 };
    assign _2056 = _2055 < _1767;
    assign _2057 = ~ _2056;
    assign _2045 = _1764[32:32];
    assign _2042 = _2037 - _1767;
    assign _2043 = _2039 ? _2042 : _2037;
    assign _2044 = _2043[62:0];
    assign _2046 = { _2044,
                     _2045 };
    assign _2047 = _2046 < _1767;
    assign _2048 = ~ _2047;
    assign _2036 = _1764[33:33];
    assign _2033 = _2028 - _1767;
    assign _2034 = _2030 ? _2033 : _2028;
    assign _2035 = _2034[62:0];
    assign _2037 = { _2035,
                     _2036 };
    assign _2038 = _2037 < _1767;
    assign _2039 = ~ _2038;
    assign _2027 = _1764[34:34];
    assign _2024 = _2019 - _1767;
    assign _2025 = _2021 ? _2024 : _2019;
    assign _2026 = _2025[62:0];
    assign _2028 = { _2026,
                     _2027 };
    assign _2029 = _2028 < _1767;
    assign _2030 = ~ _2029;
    assign _2018 = _1764[35:35];
    assign _2015 = _2010 - _1767;
    assign _2016 = _2012 ? _2015 : _2010;
    assign _2017 = _2016[62:0];
    assign _2019 = { _2017,
                     _2018 };
    assign _2020 = _2019 < _1767;
    assign _2021 = ~ _2020;
    assign _2009 = _1764[36:36];
    assign _2006 = _2001 - _1767;
    assign _2007 = _2003 ? _2006 : _2001;
    assign _2008 = _2007[62:0];
    assign _2010 = { _2008,
                     _2009 };
    assign _2011 = _2010 < _1767;
    assign _2012 = ~ _2011;
    assign _2000 = _1764[37:37];
    assign _1997 = _1992 - _1767;
    assign _1998 = _1994 ? _1997 : _1992;
    assign _1999 = _1998[62:0];
    assign _2001 = { _1999,
                     _2000 };
    assign _2002 = _2001 < _1767;
    assign _2003 = ~ _2002;
    assign _1991 = _1764[38:38];
    assign _1988 = _1983 - _1767;
    assign _1989 = _1985 ? _1988 : _1983;
    assign _1990 = _1989[62:0];
    assign _1992 = { _1990,
                     _1991 };
    assign _1993 = _1992 < _1767;
    assign _1994 = ~ _1993;
    assign _1982 = _1764[39:39];
    assign _1979 = _1974 - _1767;
    assign _1980 = _1976 ? _1979 : _1974;
    assign _1981 = _1980[62:0];
    assign _1983 = { _1981,
                     _1982 };
    assign _1984 = _1983 < _1767;
    assign _1985 = ~ _1984;
    assign _1973 = _1764[40:40];
    assign _1970 = _1965 - _1767;
    assign _1971 = _1967 ? _1970 : _1965;
    assign _1972 = _1971[62:0];
    assign _1974 = { _1972,
                     _1973 };
    assign _1975 = _1974 < _1767;
    assign _1976 = ~ _1975;
    assign _1964 = _1764[41:41];
    assign _1961 = _1956 - _1767;
    assign _1962 = _1958 ? _1961 : _1956;
    assign _1963 = _1962[62:0];
    assign _1965 = { _1963,
                     _1964 };
    assign _1966 = _1965 < _1767;
    assign _1967 = ~ _1966;
    assign _1955 = _1764[42:42];
    assign _1952 = _1947 - _1767;
    assign _1953 = _1949 ? _1952 : _1947;
    assign _1954 = _1953[62:0];
    assign _1956 = { _1954,
                     _1955 };
    assign _1957 = _1956 < _1767;
    assign _1958 = ~ _1957;
    assign _1946 = _1764[43:43];
    assign _1943 = _1938 - _1767;
    assign _1944 = _1940 ? _1943 : _1938;
    assign _1945 = _1944[62:0];
    assign _1947 = { _1945,
                     _1946 };
    assign _1948 = _1947 < _1767;
    assign _1949 = ~ _1948;
    assign _1937 = _1764[44:44];
    assign _1934 = _1929 - _1767;
    assign _1935 = _1931 ? _1934 : _1929;
    assign _1936 = _1935[62:0];
    assign _1938 = { _1936,
                     _1937 };
    assign _1939 = _1938 < _1767;
    assign _1940 = ~ _1939;
    assign _1928 = _1764[45:45];
    assign _1925 = _1920 - _1767;
    assign _1926 = _1922 ? _1925 : _1920;
    assign _1927 = _1926[62:0];
    assign _1929 = { _1927,
                     _1928 };
    assign _1930 = _1929 < _1767;
    assign _1931 = ~ _1930;
    assign _1919 = _1764[46:46];
    assign _1916 = _1911 - _1767;
    assign _1917 = _1913 ? _1916 : _1911;
    assign _1918 = _1917[62:0];
    assign _1920 = { _1918,
                     _1919 };
    assign _1921 = _1920 < _1767;
    assign _1922 = ~ _1921;
    assign _1910 = _1764[47:47];
    assign _1907 = _1902 - _1767;
    assign _1908 = _1904 ? _1907 : _1902;
    assign _1909 = _1908[62:0];
    assign _1911 = { _1909,
                     _1910 };
    assign _1912 = _1911 < _1767;
    assign _1913 = ~ _1912;
    assign _1901 = _1764[48:48];
    assign _1898 = _1893 - _1767;
    assign _1899 = _1895 ? _1898 : _1893;
    assign _1900 = _1899[62:0];
    assign _1902 = { _1900,
                     _1901 };
    assign _1903 = _1902 < _1767;
    assign _1904 = ~ _1903;
    assign _1892 = _1764[49:49];
    assign _1889 = _1884 - _1767;
    assign _1890 = _1886 ? _1889 : _1884;
    assign _1891 = _1890[62:0];
    assign _1893 = { _1891,
                     _1892 };
    assign _1894 = _1893 < _1767;
    assign _1895 = ~ _1894;
    assign _1883 = _1764[50:50];
    assign _1880 = _1875 - _1767;
    assign _1881 = _1877 ? _1880 : _1875;
    assign _1882 = _1881[62:0];
    assign _1884 = { _1882,
                     _1883 };
    assign _1885 = _1884 < _1767;
    assign _1886 = ~ _1885;
    assign _1874 = _1764[51:51];
    assign _1871 = _1866 - _1767;
    assign _1872 = _1868 ? _1871 : _1866;
    assign _1873 = _1872[62:0];
    assign _1875 = { _1873,
                     _1874 };
    assign _1876 = _1875 < _1767;
    assign _1877 = ~ _1876;
    assign _1865 = _1764[52:52];
    assign _1862 = _1857 - _1767;
    assign _1863 = _1859 ? _1862 : _1857;
    assign _1864 = _1863[62:0];
    assign _1866 = { _1864,
                     _1865 };
    assign _1867 = _1866 < _1767;
    assign _1868 = ~ _1867;
    assign _1856 = _1764[53:53];
    assign _1853 = _1848 - _1767;
    assign _1854 = _1850 ? _1853 : _1848;
    assign _1855 = _1854[62:0];
    assign _1857 = { _1855,
                     _1856 };
    assign _1858 = _1857 < _1767;
    assign _1859 = ~ _1858;
    assign _1847 = _1764[54:54];
    assign _1844 = _1839 - _1767;
    assign _1845 = _1841 ? _1844 : _1839;
    assign _1846 = _1845[62:0];
    assign _1848 = { _1846,
                     _1847 };
    assign _1849 = _1848 < _1767;
    assign _1850 = ~ _1849;
    assign _1838 = _1764[55:55];
    assign _1835 = _1830 - _1767;
    assign _1836 = _1832 ? _1835 : _1830;
    assign _1837 = _1836[62:0];
    assign _1839 = { _1837,
                     _1838 };
    assign _1840 = _1839 < _1767;
    assign _1841 = ~ _1840;
    assign _1829 = _1764[56:56];
    assign _1826 = _1821 - _1767;
    assign _1827 = _1823 ? _1826 : _1821;
    assign _1828 = _1827[62:0];
    assign _1830 = { _1828,
                     _1829 };
    assign _1831 = _1830 < _1767;
    assign _1832 = ~ _1831;
    assign _1820 = _1764[57:57];
    assign _1817 = _1812 - _1767;
    assign _1818 = _1814 ? _1817 : _1812;
    assign _1819 = _1818[62:0];
    assign _1821 = { _1819,
                     _1820 };
    assign _1822 = _1821 < _1767;
    assign _1823 = ~ _1822;
    assign _1811 = _1764[58:58];
    assign _1808 = _1803 - _1767;
    assign _1809 = _1805 ? _1808 : _1803;
    assign _1810 = _1809[62:0];
    assign _1812 = { _1810,
                     _1811 };
    assign _1813 = _1812 < _1767;
    assign _1814 = ~ _1813;
    assign _1802 = _1764[59:59];
    assign _1799 = _1794 - _1767;
    assign _1800 = _1796 ? _1799 : _1794;
    assign _1801 = _1800[62:0];
    assign _1803 = { _1801,
                     _1802 };
    assign _1804 = _1803 < _1767;
    assign _1805 = ~ _1804;
    assign _1793 = _1764[60:60];
    assign _1790 = _1785 - _1767;
    assign _1791 = _1787 ? _1790 : _1785;
    assign _1792 = _1791[62:0];
    assign _1794 = { _1792,
                     _1793 };
    assign _1795 = _1794 < _1767;
    assign _1796 = ~ _1795;
    assign _1784 = _1764[61:61];
    assign _1781 = _1776 - _1767;
    assign _1782 = _1778 ? _1781 : _1776;
    assign _1783 = _1782[62:0];
    assign _1785 = { _1783,
                     _1784 };
    assign _1786 = _1785 < _1767;
    assign _1787 = ~ _1786;
    assign _1775 = _1764[62:62];
    assign _1772 = _1766 - _1767;
    assign _1773 = _1769 ? _1772 : _1766;
    assign _1774 = _1773[62:0];
    assign _1776 = { _1774,
                     _1775 };
    assign _1777 = _1776 < _1767;
    assign _1778 = ~ _1777;
    assign _1767 = 64'b0000000000000000000000000000000000000000000000000000000001100101;
    assign _1763 = 64'b0000000000000000000000000000000000000000000000000000000001100100;
    assign _1764 = _3 + _1763;
    assign _1765 = _1764[63:63];
    assign _1766 = { _22185,
                     _1765 };
    assign _1768 = _1766 < _1767;
    assign _1769 = ~ _1768;
    assign _1770 = { _22185,
                     _1769 };
    assign _1771 = _1770[62:0];
    assign _1779 = { _1771,
                     _1778 };
    assign _1780 = _1779[62:0];
    assign _1788 = { _1780,
                     _1787 };
    assign _1789 = _1788[62:0];
    assign _1797 = { _1789,
                     _1796 };
    assign _1798 = _1797[62:0];
    assign _1806 = { _1798,
                     _1805 };
    assign _1807 = _1806[62:0];
    assign _1815 = { _1807,
                     _1814 };
    assign _1816 = _1815[62:0];
    assign _1824 = { _1816,
                     _1823 };
    assign _1825 = _1824[62:0];
    assign _1833 = { _1825,
                     _1832 };
    assign _1834 = _1833[62:0];
    assign _1842 = { _1834,
                     _1841 };
    assign _1843 = _1842[62:0];
    assign _1851 = { _1843,
                     _1850 };
    assign _1852 = _1851[62:0];
    assign _1860 = { _1852,
                     _1859 };
    assign _1861 = _1860[62:0];
    assign _1869 = { _1861,
                     _1868 };
    assign _1870 = _1869[62:0];
    assign _1878 = { _1870,
                     _1877 };
    assign _1879 = _1878[62:0];
    assign _1887 = { _1879,
                     _1886 };
    assign _1888 = _1887[62:0];
    assign _1896 = { _1888,
                     _1895 };
    assign _1897 = _1896[62:0];
    assign _1905 = { _1897,
                     _1904 };
    assign _1906 = _1905[62:0];
    assign _1914 = { _1906,
                     _1913 };
    assign _1915 = _1914[62:0];
    assign _1923 = { _1915,
                     _1922 };
    assign _1924 = _1923[62:0];
    assign _1932 = { _1924,
                     _1931 };
    assign _1933 = _1932[62:0];
    assign _1941 = { _1933,
                     _1940 };
    assign _1942 = _1941[62:0];
    assign _1950 = { _1942,
                     _1949 };
    assign _1951 = _1950[62:0];
    assign _1959 = { _1951,
                     _1958 };
    assign _1960 = _1959[62:0];
    assign _1968 = { _1960,
                     _1967 };
    assign _1969 = _1968[62:0];
    assign _1977 = { _1969,
                     _1976 };
    assign _1978 = _1977[62:0];
    assign _1986 = { _1978,
                     _1985 };
    assign _1987 = _1986[62:0];
    assign _1995 = { _1987,
                     _1994 };
    assign _1996 = _1995[62:0];
    assign _2004 = { _1996,
                     _2003 };
    assign _2005 = _2004[62:0];
    assign _2013 = { _2005,
                     _2012 };
    assign _2014 = _2013[62:0];
    assign _2022 = { _2014,
                     _2021 };
    assign _2023 = _2022[62:0];
    assign _2031 = { _2023,
                     _2030 };
    assign _2032 = _2031[62:0];
    assign _2040 = { _2032,
                     _2039 };
    assign _2041 = _2040[62:0];
    assign _2049 = { _2041,
                     _2048 };
    assign _2050 = _2049[62:0];
    assign _2058 = { _2050,
                     _2057 };
    assign _2059 = _2058[62:0];
    assign _2067 = { _2059,
                     _2066 };
    assign _2068 = _2067[62:0];
    assign _2076 = { _2068,
                     _2075 };
    assign _2077 = _2076[62:0];
    assign _2085 = { _2077,
                     _2084 };
    assign _2086 = _2085[62:0];
    assign _2094 = { _2086,
                     _2093 };
    assign _2095 = _2094[62:0];
    assign _2103 = { _2095,
                     _2102 };
    assign _2104 = _2103[62:0];
    assign _2112 = { _2104,
                     _2111 };
    assign _2113 = _2112[62:0];
    assign _2121 = { _2113,
                     _2120 };
    assign _2122 = _2121[62:0];
    assign _2130 = { _2122,
                     _2129 };
    assign _2131 = _2130[62:0];
    assign _2139 = { _2131,
                     _2138 };
    assign _2140 = _2139[62:0];
    assign _2148 = { _2140,
                     _2147 };
    assign _2149 = _2148[62:0];
    assign _2157 = { _2149,
                     _2156 };
    assign _2158 = _2157[62:0];
    assign _2166 = { _2158,
                     _2165 };
    assign _2167 = _2166[62:0];
    assign _2175 = { _2167,
                     _2174 };
    assign _2176 = _2175[62:0];
    assign _2184 = { _2176,
                     _2183 };
    assign _2185 = _2184[62:0];
    assign _2193 = { _2185,
                     _2192 };
    assign _2194 = _2193[62:0];
    assign _2202 = { _2194,
                     _2201 };
    assign _2203 = _2202[62:0];
    assign _2211 = { _2203,
                     _2210 };
    assign _2212 = _2211[62:0];
    assign _2220 = { _2212,
                     _2219 };
    assign _2221 = _2220[62:0];
    assign _2229 = { _2221,
                     _2228 };
    assign _2230 = _2229[62:0];
    assign _2238 = { _2230,
                     _2237 };
    assign _2239 = _2238[62:0];
    assign _2247 = { _2239,
                     _2246 };
    assign _2248 = _2247[62:0];
    assign _2256 = { _2248,
                     _2255 };
    assign _2257 = _2256[62:0];
    assign _2265 = { _2257,
                     _2264 };
    assign _2266 = _2265[62:0];
    assign _2274 = { _2266,
                     _2273 };
    assign _2275 = _2274[62:0];
    assign _2283 = { _2275,
                     _2282 };
    assign _2284 = _2283[62:0];
    assign _2292 = { _2284,
                     _2291 };
    assign _2293 = _2292[62:0];
    assign _2301 = { _2293,
                     _2300 };
    assign _2302 = _2301[62:0];
    assign _2310 = { _2302,
                     _2309 };
    assign _2311 = _2310[62:0];
    assign _2319 = { _2311,
                     _2318 };
    assign _2320 = _2319[62:0];
    assign _2328 = { _2320,
                     _2327 };
    assign _2329 = _2328[62:0];
    assign _2337 = { _2329,
                     _2336 };
    assign _2338 = _2337 * _1767;
    assign _2339 = _2338[63:0];
    assign _1760 = 64'b0000000000000000000000000000000000000000000000000000001111110010;
    assign _2340 = _1760 < _2339;
    assign _2341 = _2340 ? _2339 : _1760;
    assign _1757 = 64'b0000000000000000000000000000000000000000000000000010011100001111;
    assign _1758 = _5 < _1757;
    assign _1759 = _1758 ? _5 : _1757;
    assign _2342 = _1759 < _2341;
    assign _2343 = ~ _2342;
    assign _3506 = _2343 ? _3505 : _21604;
    assign _1748 = _1179[0:0];
    assign _1745 = _1740 - _22192;
    assign _1746 = _1742 ? _1745 : _1740;
    assign _1747 = _1746[62:0];
    assign _1749 = { _1747,
                     _1748 };
    assign _1750 = _1749 < _22192;
    assign _1751 = ~ _1750;
    assign _1739 = _1179[1:1];
    assign _1736 = _1731 - _22192;
    assign _1737 = _1733 ? _1736 : _1731;
    assign _1738 = _1737[62:0];
    assign _1740 = { _1738,
                     _1739 };
    assign _1741 = _1740 < _22192;
    assign _1742 = ~ _1741;
    assign _1730 = _1179[2:2];
    assign _1727 = _1722 - _22192;
    assign _1728 = _1724 ? _1727 : _1722;
    assign _1729 = _1728[62:0];
    assign _1731 = { _1729,
                     _1730 };
    assign _1732 = _1731 < _22192;
    assign _1733 = ~ _1732;
    assign _1721 = _1179[3:3];
    assign _1718 = _1713 - _22192;
    assign _1719 = _1715 ? _1718 : _1713;
    assign _1720 = _1719[62:0];
    assign _1722 = { _1720,
                     _1721 };
    assign _1723 = _1722 < _22192;
    assign _1724 = ~ _1723;
    assign _1712 = _1179[4:4];
    assign _1709 = _1704 - _22192;
    assign _1710 = _1706 ? _1709 : _1704;
    assign _1711 = _1710[62:0];
    assign _1713 = { _1711,
                     _1712 };
    assign _1714 = _1713 < _22192;
    assign _1715 = ~ _1714;
    assign _1703 = _1179[5:5];
    assign _1700 = _1695 - _22192;
    assign _1701 = _1697 ? _1700 : _1695;
    assign _1702 = _1701[62:0];
    assign _1704 = { _1702,
                     _1703 };
    assign _1705 = _1704 < _22192;
    assign _1706 = ~ _1705;
    assign _1694 = _1179[6:6];
    assign _1691 = _1686 - _22192;
    assign _1692 = _1688 ? _1691 : _1686;
    assign _1693 = _1692[62:0];
    assign _1695 = { _1693,
                     _1694 };
    assign _1696 = _1695 < _22192;
    assign _1697 = ~ _1696;
    assign _1685 = _1179[7:7];
    assign _1682 = _1677 - _22192;
    assign _1683 = _1679 ? _1682 : _1677;
    assign _1684 = _1683[62:0];
    assign _1686 = { _1684,
                     _1685 };
    assign _1687 = _1686 < _22192;
    assign _1688 = ~ _1687;
    assign _1676 = _1179[8:8];
    assign _1673 = _1668 - _22192;
    assign _1674 = _1670 ? _1673 : _1668;
    assign _1675 = _1674[62:0];
    assign _1677 = { _1675,
                     _1676 };
    assign _1678 = _1677 < _22192;
    assign _1679 = ~ _1678;
    assign _1667 = _1179[9:9];
    assign _1664 = _1659 - _22192;
    assign _1665 = _1661 ? _1664 : _1659;
    assign _1666 = _1665[62:0];
    assign _1668 = { _1666,
                     _1667 };
    assign _1669 = _1668 < _22192;
    assign _1670 = ~ _1669;
    assign _1658 = _1179[10:10];
    assign _1655 = _1650 - _22192;
    assign _1656 = _1652 ? _1655 : _1650;
    assign _1657 = _1656[62:0];
    assign _1659 = { _1657,
                     _1658 };
    assign _1660 = _1659 < _22192;
    assign _1661 = ~ _1660;
    assign _1649 = _1179[11:11];
    assign _1646 = _1641 - _22192;
    assign _1647 = _1643 ? _1646 : _1641;
    assign _1648 = _1647[62:0];
    assign _1650 = { _1648,
                     _1649 };
    assign _1651 = _1650 < _22192;
    assign _1652 = ~ _1651;
    assign _1640 = _1179[12:12];
    assign _1637 = _1632 - _22192;
    assign _1638 = _1634 ? _1637 : _1632;
    assign _1639 = _1638[62:0];
    assign _1641 = { _1639,
                     _1640 };
    assign _1642 = _1641 < _22192;
    assign _1643 = ~ _1642;
    assign _1631 = _1179[13:13];
    assign _1628 = _1623 - _22192;
    assign _1629 = _1625 ? _1628 : _1623;
    assign _1630 = _1629[62:0];
    assign _1632 = { _1630,
                     _1631 };
    assign _1633 = _1632 < _22192;
    assign _1634 = ~ _1633;
    assign _1622 = _1179[14:14];
    assign _1619 = _1614 - _22192;
    assign _1620 = _1616 ? _1619 : _1614;
    assign _1621 = _1620[62:0];
    assign _1623 = { _1621,
                     _1622 };
    assign _1624 = _1623 < _22192;
    assign _1625 = ~ _1624;
    assign _1613 = _1179[15:15];
    assign _1610 = _1605 - _22192;
    assign _1611 = _1607 ? _1610 : _1605;
    assign _1612 = _1611[62:0];
    assign _1614 = { _1612,
                     _1613 };
    assign _1615 = _1614 < _22192;
    assign _1616 = ~ _1615;
    assign _1604 = _1179[16:16];
    assign _1601 = _1596 - _22192;
    assign _1602 = _1598 ? _1601 : _1596;
    assign _1603 = _1602[62:0];
    assign _1605 = { _1603,
                     _1604 };
    assign _1606 = _1605 < _22192;
    assign _1607 = ~ _1606;
    assign _1595 = _1179[17:17];
    assign _1592 = _1587 - _22192;
    assign _1593 = _1589 ? _1592 : _1587;
    assign _1594 = _1593[62:0];
    assign _1596 = { _1594,
                     _1595 };
    assign _1597 = _1596 < _22192;
    assign _1598 = ~ _1597;
    assign _1586 = _1179[18:18];
    assign _1583 = _1578 - _22192;
    assign _1584 = _1580 ? _1583 : _1578;
    assign _1585 = _1584[62:0];
    assign _1587 = { _1585,
                     _1586 };
    assign _1588 = _1587 < _22192;
    assign _1589 = ~ _1588;
    assign _1577 = _1179[19:19];
    assign _1574 = _1569 - _22192;
    assign _1575 = _1571 ? _1574 : _1569;
    assign _1576 = _1575[62:0];
    assign _1578 = { _1576,
                     _1577 };
    assign _1579 = _1578 < _22192;
    assign _1580 = ~ _1579;
    assign _1568 = _1179[20:20];
    assign _1565 = _1560 - _22192;
    assign _1566 = _1562 ? _1565 : _1560;
    assign _1567 = _1566[62:0];
    assign _1569 = { _1567,
                     _1568 };
    assign _1570 = _1569 < _22192;
    assign _1571 = ~ _1570;
    assign _1559 = _1179[21:21];
    assign _1556 = _1551 - _22192;
    assign _1557 = _1553 ? _1556 : _1551;
    assign _1558 = _1557[62:0];
    assign _1560 = { _1558,
                     _1559 };
    assign _1561 = _1560 < _22192;
    assign _1562 = ~ _1561;
    assign _1550 = _1179[22:22];
    assign _1547 = _1542 - _22192;
    assign _1548 = _1544 ? _1547 : _1542;
    assign _1549 = _1548[62:0];
    assign _1551 = { _1549,
                     _1550 };
    assign _1552 = _1551 < _22192;
    assign _1553 = ~ _1552;
    assign _1541 = _1179[23:23];
    assign _1538 = _1533 - _22192;
    assign _1539 = _1535 ? _1538 : _1533;
    assign _1540 = _1539[62:0];
    assign _1542 = { _1540,
                     _1541 };
    assign _1543 = _1542 < _22192;
    assign _1544 = ~ _1543;
    assign _1532 = _1179[24:24];
    assign _1529 = _1524 - _22192;
    assign _1530 = _1526 ? _1529 : _1524;
    assign _1531 = _1530[62:0];
    assign _1533 = { _1531,
                     _1532 };
    assign _1534 = _1533 < _22192;
    assign _1535 = ~ _1534;
    assign _1523 = _1179[25:25];
    assign _1520 = _1515 - _22192;
    assign _1521 = _1517 ? _1520 : _1515;
    assign _1522 = _1521[62:0];
    assign _1524 = { _1522,
                     _1523 };
    assign _1525 = _1524 < _22192;
    assign _1526 = ~ _1525;
    assign _1514 = _1179[26:26];
    assign _1511 = _1506 - _22192;
    assign _1512 = _1508 ? _1511 : _1506;
    assign _1513 = _1512[62:0];
    assign _1515 = { _1513,
                     _1514 };
    assign _1516 = _1515 < _22192;
    assign _1517 = ~ _1516;
    assign _1505 = _1179[27:27];
    assign _1502 = _1497 - _22192;
    assign _1503 = _1499 ? _1502 : _1497;
    assign _1504 = _1503[62:0];
    assign _1506 = { _1504,
                     _1505 };
    assign _1507 = _1506 < _22192;
    assign _1508 = ~ _1507;
    assign _1496 = _1179[28:28];
    assign _1493 = _1488 - _22192;
    assign _1494 = _1490 ? _1493 : _1488;
    assign _1495 = _1494[62:0];
    assign _1497 = { _1495,
                     _1496 };
    assign _1498 = _1497 < _22192;
    assign _1499 = ~ _1498;
    assign _1487 = _1179[29:29];
    assign _1484 = _1479 - _22192;
    assign _1485 = _1481 ? _1484 : _1479;
    assign _1486 = _1485[62:0];
    assign _1488 = { _1486,
                     _1487 };
    assign _1489 = _1488 < _22192;
    assign _1490 = ~ _1489;
    assign _1478 = _1179[30:30];
    assign _1475 = _1470 - _22192;
    assign _1476 = _1472 ? _1475 : _1470;
    assign _1477 = _1476[62:0];
    assign _1479 = { _1477,
                     _1478 };
    assign _1480 = _1479 < _22192;
    assign _1481 = ~ _1480;
    assign _1469 = _1179[31:31];
    assign _1466 = _1461 - _22192;
    assign _1467 = _1463 ? _1466 : _1461;
    assign _1468 = _1467[62:0];
    assign _1470 = { _1468,
                     _1469 };
    assign _1471 = _1470 < _22192;
    assign _1472 = ~ _1471;
    assign _1460 = _1179[32:32];
    assign _1457 = _1452 - _22192;
    assign _1458 = _1454 ? _1457 : _1452;
    assign _1459 = _1458[62:0];
    assign _1461 = { _1459,
                     _1460 };
    assign _1462 = _1461 < _22192;
    assign _1463 = ~ _1462;
    assign _1451 = _1179[33:33];
    assign _1448 = _1443 - _22192;
    assign _1449 = _1445 ? _1448 : _1443;
    assign _1450 = _1449[62:0];
    assign _1452 = { _1450,
                     _1451 };
    assign _1453 = _1452 < _22192;
    assign _1454 = ~ _1453;
    assign _1442 = _1179[34:34];
    assign _1439 = _1434 - _22192;
    assign _1440 = _1436 ? _1439 : _1434;
    assign _1441 = _1440[62:0];
    assign _1443 = { _1441,
                     _1442 };
    assign _1444 = _1443 < _22192;
    assign _1445 = ~ _1444;
    assign _1433 = _1179[35:35];
    assign _1430 = _1425 - _22192;
    assign _1431 = _1427 ? _1430 : _1425;
    assign _1432 = _1431[62:0];
    assign _1434 = { _1432,
                     _1433 };
    assign _1435 = _1434 < _22192;
    assign _1436 = ~ _1435;
    assign _1424 = _1179[36:36];
    assign _1421 = _1416 - _22192;
    assign _1422 = _1418 ? _1421 : _1416;
    assign _1423 = _1422[62:0];
    assign _1425 = { _1423,
                     _1424 };
    assign _1426 = _1425 < _22192;
    assign _1427 = ~ _1426;
    assign _1415 = _1179[37:37];
    assign _1412 = _1407 - _22192;
    assign _1413 = _1409 ? _1412 : _1407;
    assign _1414 = _1413[62:0];
    assign _1416 = { _1414,
                     _1415 };
    assign _1417 = _1416 < _22192;
    assign _1418 = ~ _1417;
    assign _1406 = _1179[38:38];
    assign _1403 = _1398 - _22192;
    assign _1404 = _1400 ? _1403 : _1398;
    assign _1405 = _1404[62:0];
    assign _1407 = { _1405,
                     _1406 };
    assign _1408 = _1407 < _22192;
    assign _1409 = ~ _1408;
    assign _1397 = _1179[39:39];
    assign _1394 = _1389 - _22192;
    assign _1395 = _1391 ? _1394 : _1389;
    assign _1396 = _1395[62:0];
    assign _1398 = { _1396,
                     _1397 };
    assign _1399 = _1398 < _22192;
    assign _1400 = ~ _1399;
    assign _1388 = _1179[40:40];
    assign _1385 = _1380 - _22192;
    assign _1386 = _1382 ? _1385 : _1380;
    assign _1387 = _1386[62:0];
    assign _1389 = { _1387,
                     _1388 };
    assign _1390 = _1389 < _22192;
    assign _1391 = ~ _1390;
    assign _1379 = _1179[41:41];
    assign _1376 = _1371 - _22192;
    assign _1377 = _1373 ? _1376 : _1371;
    assign _1378 = _1377[62:0];
    assign _1380 = { _1378,
                     _1379 };
    assign _1381 = _1380 < _22192;
    assign _1382 = ~ _1381;
    assign _1370 = _1179[42:42];
    assign _1367 = _1362 - _22192;
    assign _1368 = _1364 ? _1367 : _1362;
    assign _1369 = _1368[62:0];
    assign _1371 = { _1369,
                     _1370 };
    assign _1372 = _1371 < _22192;
    assign _1373 = ~ _1372;
    assign _1361 = _1179[43:43];
    assign _1358 = _1353 - _22192;
    assign _1359 = _1355 ? _1358 : _1353;
    assign _1360 = _1359[62:0];
    assign _1362 = { _1360,
                     _1361 };
    assign _1363 = _1362 < _22192;
    assign _1364 = ~ _1363;
    assign _1352 = _1179[44:44];
    assign _1349 = _1344 - _22192;
    assign _1350 = _1346 ? _1349 : _1344;
    assign _1351 = _1350[62:0];
    assign _1353 = { _1351,
                     _1352 };
    assign _1354 = _1353 < _22192;
    assign _1355 = ~ _1354;
    assign _1343 = _1179[45:45];
    assign _1340 = _1335 - _22192;
    assign _1341 = _1337 ? _1340 : _1335;
    assign _1342 = _1341[62:0];
    assign _1344 = { _1342,
                     _1343 };
    assign _1345 = _1344 < _22192;
    assign _1346 = ~ _1345;
    assign _1334 = _1179[46:46];
    assign _1331 = _1326 - _22192;
    assign _1332 = _1328 ? _1331 : _1326;
    assign _1333 = _1332[62:0];
    assign _1335 = { _1333,
                     _1334 };
    assign _1336 = _1335 < _22192;
    assign _1337 = ~ _1336;
    assign _1325 = _1179[47:47];
    assign _1322 = _1317 - _22192;
    assign _1323 = _1319 ? _1322 : _1317;
    assign _1324 = _1323[62:0];
    assign _1326 = { _1324,
                     _1325 };
    assign _1327 = _1326 < _22192;
    assign _1328 = ~ _1327;
    assign _1316 = _1179[48:48];
    assign _1313 = _1308 - _22192;
    assign _1314 = _1310 ? _1313 : _1308;
    assign _1315 = _1314[62:0];
    assign _1317 = { _1315,
                     _1316 };
    assign _1318 = _1317 < _22192;
    assign _1319 = ~ _1318;
    assign _1307 = _1179[49:49];
    assign _1304 = _1299 - _22192;
    assign _1305 = _1301 ? _1304 : _1299;
    assign _1306 = _1305[62:0];
    assign _1308 = { _1306,
                     _1307 };
    assign _1309 = _1308 < _22192;
    assign _1310 = ~ _1309;
    assign _1298 = _1179[50:50];
    assign _1295 = _1290 - _22192;
    assign _1296 = _1292 ? _1295 : _1290;
    assign _1297 = _1296[62:0];
    assign _1299 = { _1297,
                     _1298 };
    assign _1300 = _1299 < _22192;
    assign _1301 = ~ _1300;
    assign _1289 = _1179[51:51];
    assign _1286 = _1281 - _22192;
    assign _1287 = _1283 ? _1286 : _1281;
    assign _1288 = _1287[62:0];
    assign _1290 = { _1288,
                     _1289 };
    assign _1291 = _1290 < _22192;
    assign _1292 = ~ _1291;
    assign _1280 = _1179[52:52];
    assign _1277 = _1272 - _22192;
    assign _1278 = _1274 ? _1277 : _1272;
    assign _1279 = _1278[62:0];
    assign _1281 = { _1279,
                     _1280 };
    assign _1282 = _1281 < _22192;
    assign _1283 = ~ _1282;
    assign _1271 = _1179[53:53];
    assign _1268 = _1263 - _22192;
    assign _1269 = _1265 ? _1268 : _1263;
    assign _1270 = _1269[62:0];
    assign _1272 = { _1270,
                     _1271 };
    assign _1273 = _1272 < _22192;
    assign _1274 = ~ _1273;
    assign _1262 = _1179[54:54];
    assign _1259 = _1254 - _22192;
    assign _1260 = _1256 ? _1259 : _1254;
    assign _1261 = _1260[62:0];
    assign _1263 = { _1261,
                     _1262 };
    assign _1264 = _1263 < _22192;
    assign _1265 = ~ _1264;
    assign _1253 = _1179[55:55];
    assign _1250 = _1245 - _22192;
    assign _1251 = _1247 ? _1250 : _1245;
    assign _1252 = _1251[62:0];
    assign _1254 = { _1252,
                     _1253 };
    assign _1255 = _1254 < _22192;
    assign _1256 = ~ _1255;
    assign _1244 = _1179[56:56];
    assign _1241 = _1236 - _22192;
    assign _1242 = _1238 ? _1241 : _1236;
    assign _1243 = _1242[62:0];
    assign _1245 = { _1243,
                     _1244 };
    assign _1246 = _1245 < _22192;
    assign _1247 = ~ _1246;
    assign _1235 = _1179[57:57];
    assign _1232 = _1227 - _22192;
    assign _1233 = _1229 ? _1232 : _1227;
    assign _1234 = _1233[62:0];
    assign _1236 = { _1234,
                     _1235 };
    assign _1237 = _1236 < _22192;
    assign _1238 = ~ _1237;
    assign _1226 = _1179[58:58];
    assign _1223 = _1218 - _22192;
    assign _1224 = _1220 ? _1223 : _1218;
    assign _1225 = _1224[62:0];
    assign _1227 = { _1225,
                     _1226 };
    assign _1228 = _1227 < _22192;
    assign _1229 = ~ _1228;
    assign _1217 = _1179[59:59];
    assign _1214 = _1209 - _22192;
    assign _1215 = _1211 ? _1214 : _1209;
    assign _1216 = _1215[62:0];
    assign _1218 = { _1216,
                     _1217 };
    assign _1219 = _1218 < _22192;
    assign _1220 = ~ _1219;
    assign _1208 = _1179[60:60];
    assign _1205 = _1200 - _22192;
    assign _1206 = _1202 ? _1205 : _1200;
    assign _1207 = _1206[62:0];
    assign _1209 = { _1207,
                     _1208 };
    assign _1210 = _1209 < _22192;
    assign _1211 = ~ _1210;
    assign _1199 = _1179[61:61];
    assign _1196 = _1191 - _22192;
    assign _1197 = _1193 ? _1196 : _1191;
    assign _1198 = _1197[62:0];
    assign _1200 = { _1198,
                     _1199 };
    assign _1201 = _1200 < _22192;
    assign _1202 = ~ _1201;
    assign _1190 = _1179[62:62];
    assign _1187 = _1181 - _22192;
    assign _1188 = _1184 ? _1187 : _1181;
    assign _1189 = _1188[62:0];
    assign _1191 = { _1189,
                     _1190 };
    assign _1192 = _1191 < _22192;
    assign _1193 = ~ _1192;
    assign _1177 = _1169 + _22186;
    assign _1178 = _1169 * _1177;
    assign _1179 = _1178[63:0];
    assign _1180 = _1179[63:63];
    assign _1181 = { _22185,
                     _1180 };
    assign _1183 = _1181 < _22192;
    assign _1184 = ~ _1183;
    assign _1185 = { _22185,
                     _1184 };
    assign _1186 = _1185[62:0];
    assign _1194 = { _1186,
                     _1193 };
    assign _1195 = _1194[62:0];
    assign _1203 = { _1195,
                     _1202 };
    assign _1204 = _1203[62:0];
    assign _1212 = { _1204,
                     _1211 };
    assign _1213 = _1212[62:0];
    assign _1221 = { _1213,
                     _1220 };
    assign _1222 = _1221[62:0];
    assign _1230 = { _1222,
                     _1229 };
    assign _1231 = _1230[62:0];
    assign _1239 = { _1231,
                     _1238 };
    assign _1240 = _1239[62:0];
    assign _1248 = { _1240,
                     _1247 };
    assign _1249 = _1248[62:0];
    assign _1257 = { _1249,
                     _1256 };
    assign _1258 = _1257[62:0];
    assign _1266 = { _1258,
                     _1265 };
    assign _1267 = _1266[62:0];
    assign _1275 = { _1267,
                     _1274 };
    assign _1276 = _1275[62:0];
    assign _1284 = { _1276,
                     _1283 };
    assign _1285 = _1284[62:0];
    assign _1293 = { _1285,
                     _1292 };
    assign _1294 = _1293[62:0];
    assign _1302 = { _1294,
                     _1301 };
    assign _1303 = _1302[62:0];
    assign _1311 = { _1303,
                     _1310 };
    assign _1312 = _1311[62:0];
    assign _1320 = { _1312,
                     _1319 };
    assign _1321 = _1320[62:0];
    assign _1329 = { _1321,
                     _1328 };
    assign _1330 = _1329[62:0];
    assign _1338 = { _1330,
                     _1337 };
    assign _1339 = _1338[62:0];
    assign _1347 = { _1339,
                     _1346 };
    assign _1348 = _1347[62:0];
    assign _1356 = { _1348,
                     _1355 };
    assign _1357 = _1356[62:0];
    assign _1365 = { _1357,
                     _1364 };
    assign _1366 = _1365[62:0];
    assign _1374 = { _1366,
                     _1373 };
    assign _1375 = _1374[62:0];
    assign _1383 = { _1375,
                     _1382 };
    assign _1384 = _1383[62:0];
    assign _1392 = { _1384,
                     _1391 };
    assign _1393 = _1392[62:0];
    assign _1401 = { _1393,
                     _1400 };
    assign _1402 = _1401[62:0];
    assign _1410 = { _1402,
                     _1409 };
    assign _1411 = _1410[62:0];
    assign _1419 = { _1411,
                     _1418 };
    assign _1420 = _1419[62:0];
    assign _1428 = { _1420,
                     _1427 };
    assign _1429 = _1428[62:0];
    assign _1437 = { _1429,
                     _1436 };
    assign _1438 = _1437[62:0];
    assign _1446 = { _1438,
                     _1445 };
    assign _1447 = _1446[62:0];
    assign _1455 = { _1447,
                     _1454 };
    assign _1456 = _1455[62:0];
    assign _1464 = { _1456,
                     _1463 };
    assign _1465 = _1464[62:0];
    assign _1473 = { _1465,
                     _1472 };
    assign _1474 = _1473[62:0];
    assign _1482 = { _1474,
                     _1481 };
    assign _1483 = _1482[62:0];
    assign _1491 = { _1483,
                     _1490 };
    assign _1492 = _1491[62:0];
    assign _1500 = { _1492,
                     _1499 };
    assign _1501 = _1500[62:0];
    assign _1509 = { _1501,
                     _1508 };
    assign _1510 = _1509[62:0];
    assign _1518 = { _1510,
                     _1517 };
    assign _1519 = _1518[62:0];
    assign _1527 = { _1519,
                     _1526 };
    assign _1528 = _1527[62:0];
    assign _1536 = { _1528,
                     _1535 };
    assign _1537 = _1536[62:0];
    assign _1545 = { _1537,
                     _1544 };
    assign _1546 = _1545[62:0];
    assign _1554 = { _1546,
                     _1553 };
    assign _1555 = _1554[62:0];
    assign _1563 = { _1555,
                     _1562 };
    assign _1564 = _1563[62:0];
    assign _1572 = { _1564,
                     _1571 };
    assign _1573 = _1572[62:0];
    assign _1581 = { _1573,
                     _1580 };
    assign _1582 = _1581[62:0];
    assign _1590 = { _1582,
                     _1589 };
    assign _1591 = _1590[62:0];
    assign _1599 = { _1591,
                     _1598 };
    assign _1600 = _1599[62:0];
    assign _1608 = { _1600,
                     _1607 };
    assign _1609 = _1608[62:0];
    assign _1617 = { _1609,
                     _1616 };
    assign _1618 = _1617[62:0];
    assign _1626 = { _1618,
                     _1625 };
    assign _1627 = _1626[62:0];
    assign _1635 = { _1627,
                     _1634 };
    assign _1636 = _1635[62:0];
    assign _1644 = { _1636,
                     _1643 };
    assign _1645 = _1644[62:0];
    assign _1653 = { _1645,
                     _1652 };
    assign _1654 = _1653[62:0];
    assign _1662 = { _1654,
                     _1661 };
    assign _1663 = _1662[62:0];
    assign _1671 = { _1663,
                     _1670 };
    assign _1672 = _1671[62:0];
    assign _1680 = { _1672,
                     _1679 };
    assign _1681 = _1680[62:0];
    assign _1689 = { _1681,
                     _1688 };
    assign _1690 = _1689[62:0];
    assign _1698 = { _1690,
                     _1697 };
    assign _1699 = _1698[62:0];
    assign _1707 = { _1699,
                     _1706 };
    assign _1708 = _1707[62:0];
    assign _1716 = { _1708,
                     _1715 };
    assign _1717 = _1716[62:0];
    assign _1725 = { _1717,
                     _1724 };
    assign _1726 = _1725[62:0];
    assign _1734 = { _1726,
                     _1733 };
    assign _1735 = _1734[62:0];
    assign _1743 = { _1735,
                     _1742 };
    assign _1744 = _1743[62:0];
    assign _1752 = { _1744,
                     _1751 };
    assign _1753 = _17 * _1752;
    assign _1754 = _1753[63:0];
    assign _1165 = _597[0:0];
    assign _1162 = _1157 - _17;
    assign _1163 = _1159 ? _1162 : _1157;
    assign _1164 = _1163[62:0];
    assign _1166 = { _1164,
                     _1165 };
    assign _1167 = _1166 < _17;
    assign _1168 = ~ _1167;
    assign _1156 = _597[1:1];
    assign _1153 = _1148 - _17;
    assign _1154 = _1150 ? _1153 : _1148;
    assign _1155 = _1154[62:0];
    assign _1157 = { _1155,
                     _1156 };
    assign _1158 = _1157 < _17;
    assign _1159 = ~ _1158;
    assign _1147 = _597[2:2];
    assign _1144 = _1139 - _17;
    assign _1145 = _1141 ? _1144 : _1139;
    assign _1146 = _1145[62:0];
    assign _1148 = { _1146,
                     _1147 };
    assign _1149 = _1148 < _17;
    assign _1150 = ~ _1149;
    assign _1138 = _597[3:3];
    assign _1135 = _1130 - _17;
    assign _1136 = _1132 ? _1135 : _1130;
    assign _1137 = _1136[62:0];
    assign _1139 = { _1137,
                     _1138 };
    assign _1140 = _1139 < _17;
    assign _1141 = ~ _1140;
    assign _1129 = _597[4:4];
    assign _1126 = _1121 - _17;
    assign _1127 = _1123 ? _1126 : _1121;
    assign _1128 = _1127[62:0];
    assign _1130 = { _1128,
                     _1129 };
    assign _1131 = _1130 < _17;
    assign _1132 = ~ _1131;
    assign _1120 = _597[5:5];
    assign _1117 = _1112 - _17;
    assign _1118 = _1114 ? _1117 : _1112;
    assign _1119 = _1118[62:0];
    assign _1121 = { _1119,
                     _1120 };
    assign _1122 = _1121 < _17;
    assign _1123 = ~ _1122;
    assign _1111 = _597[6:6];
    assign _1108 = _1103 - _17;
    assign _1109 = _1105 ? _1108 : _1103;
    assign _1110 = _1109[62:0];
    assign _1112 = { _1110,
                     _1111 };
    assign _1113 = _1112 < _17;
    assign _1114 = ~ _1113;
    assign _1102 = _597[7:7];
    assign _1099 = _1094 - _17;
    assign _1100 = _1096 ? _1099 : _1094;
    assign _1101 = _1100[62:0];
    assign _1103 = { _1101,
                     _1102 };
    assign _1104 = _1103 < _17;
    assign _1105 = ~ _1104;
    assign _1093 = _597[8:8];
    assign _1090 = _1085 - _17;
    assign _1091 = _1087 ? _1090 : _1085;
    assign _1092 = _1091[62:0];
    assign _1094 = { _1092,
                     _1093 };
    assign _1095 = _1094 < _17;
    assign _1096 = ~ _1095;
    assign _1084 = _597[9:9];
    assign _1081 = _1076 - _17;
    assign _1082 = _1078 ? _1081 : _1076;
    assign _1083 = _1082[62:0];
    assign _1085 = { _1083,
                     _1084 };
    assign _1086 = _1085 < _17;
    assign _1087 = ~ _1086;
    assign _1075 = _597[10:10];
    assign _1072 = _1067 - _17;
    assign _1073 = _1069 ? _1072 : _1067;
    assign _1074 = _1073[62:0];
    assign _1076 = { _1074,
                     _1075 };
    assign _1077 = _1076 < _17;
    assign _1078 = ~ _1077;
    assign _1066 = _597[11:11];
    assign _1063 = _1058 - _17;
    assign _1064 = _1060 ? _1063 : _1058;
    assign _1065 = _1064[62:0];
    assign _1067 = { _1065,
                     _1066 };
    assign _1068 = _1067 < _17;
    assign _1069 = ~ _1068;
    assign _1057 = _597[12:12];
    assign _1054 = _1049 - _17;
    assign _1055 = _1051 ? _1054 : _1049;
    assign _1056 = _1055[62:0];
    assign _1058 = { _1056,
                     _1057 };
    assign _1059 = _1058 < _17;
    assign _1060 = ~ _1059;
    assign _1048 = _597[13:13];
    assign _1045 = _1040 - _17;
    assign _1046 = _1042 ? _1045 : _1040;
    assign _1047 = _1046[62:0];
    assign _1049 = { _1047,
                     _1048 };
    assign _1050 = _1049 < _17;
    assign _1051 = ~ _1050;
    assign _1039 = _597[14:14];
    assign _1036 = _1031 - _17;
    assign _1037 = _1033 ? _1036 : _1031;
    assign _1038 = _1037[62:0];
    assign _1040 = { _1038,
                     _1039 };
    assign _1041 = _1040 < _17;
    assign _1042 = ~ _1041;
    assign _1030 = _597[15:15];
    assign _1027 = _1022 - _17;
    assign _1028 = _1024 ? _1027 : _1022;
    assign _1029 = _1028[62:0];
    assign _1031 = { _1029,
                     _1030 };
    assign _1032 = _1031 < _17;
    assign _1033 = ~ _1032;
    assign _1021 = _597[16:16];
    assign _1018 = _1013 - _17;
    assign _1019 = _1015 ? _1018 : _1013;
    assign _1020 = _1019[62:0];
    assign _1022 = { _1020,
                     _1021 };
    assign _1023 = _1022 < _17;
    assign _1024 = ~ _1023;
    assign _1012 = _597[17:17];
    assign _1009 = _1004 - _17;
    assign _1010 = _1006 ? _1009 : _1004;
    assign _1011 = _1010[62:0];
    assign _1013 = { _1011,
                     _1012 };
    assign _1014 = _1013 < _17;
    assign _1015 = ~ _1014;
    assign _1003 = _597[18:18];
    assign _1000 = _995 - _17;
    assign _1001 = _997 ? _1000 : _995;
    assign _1002 = _1001[62:0];
    assign _1004 = { _1002,
                     _1003 };
    assign _1005 = _1004 < _17;
    assign _1006 = ~ _1005;
    assign _994 = _597[19:19];
    assign _991 = _986 - _17;
    assign _992 = _988 ? _991 : _986;
    assign _993 = _992[62:0];
    assign _995 = { _993,
                    _994 };
    assign _996 = _995 < _17;
    assign _997 = ~ _996;
    assign _985 = _597[20:20];
    assign _982 = _977 - _17;
    assign _983 = _979 ? _982 : _977;
    assign _984 = _983[62:0];
    assign _986 = { _984,
                    _985 };
    assign _987 = _986 < _17;
    assign _988 = ~ _987;
    assign _976 = _597[21:21];
    assign _973 = _968 - _17;
    assign _974 = _970 ? _973 : _968;
    assign _975 = _974[62:0];
    assign _977 = { _975,
                    _976 };
    assign _978 = _977 < _17;
    assign _979 = ~ _978;
    assign _967 = _597[22:22];
    assign _964 = _959 - _17;
    assign _965 = _961 ? _964 : _959;
    assign _966 = _965[62:0];
    assign _968 = { _966,
                    _967 };
    assign _969 = _968 < _17;
    assign _970 = ~ _969;
    assign _958 = _597[23:23];
    assign _955 = _950 - _17;
    assign _956 = _952 ? _955 : _950;
    assign _957 = _956[62:0];
    assign _959 = { _957,
                    _958 };
    assign _960 = _959 < _17;
    assign _961 = ~ _960;
    assign _949 = _597[24:24];
    assign _946 = _941 - _17;
    assign _947 = _943 ? _946 : _941;
    assign _948 = _947[62:0];
    assign _950 = { _948,
                    _949 };
    assign _951 = _950 < _17;
    assign _952 = ~ _951;
    assign _940 = _597[25:25];
    assign _937 = _932 - _17;
    assign _938 = _934 ? _937 : _932;
    assign _939 = _938[62:0];
    assign _941 = { _939,
                    _940 };
    assign _942 = _941 < _17;
    assign _943 = ~ _942;
    assign _931 = _597[26:26];
    assign _928 = _923 - _17;
    assign _929 = _925 ? _928 : _923;
    assign _930 = _929[62:0];
    assign _932 = { _930,
                    _931 };
    assign _933 = _932 < _17;
    assign _934 = ~ _933;
    assign _922 = _597[27:27];
    assign _919 = _914 - _17;
    assign _920 = _916 ? _919 : _914;
    assign _921 = _920[62:0];
    assign _923 = { _921,
                    _922 };
    assign _924 = _923 < _17;
    assign _925 = ~ _924;
    assign _913 = _597[28:28];
    assign _910 = _905 - _17;
    assign _911 = _907 ? _910 : _905;
    assign _912 = _911[62:0];
    assign _914 = { _912,
                    _913 };
    assign _915 = _914 < _17;
    assign _916 = ~ _915;
    assign _904 = _597[29:29];
    assign _901 = _896 - _17;
    assign _902 = _898 ? _901 : _896;
    assign _903 = _902[62:0];
    assign _905 = { _903,
                    _904 };
    assign _906 = _905 < _17;
    assign _907 = ~ _906;
    assign _895 = _597[30:30];
    assign _892 = _887 - _17;
    assign _893 = _889 ? _892 : _887;
    assign _894 = _893[62:0];
    assign _896 = { _894,
                    _895 };
    assign _897 = _896 < _17;
    assign _898 = ~ _897;
    assign _886 = _597[31:31];
    assign _883 = _878 - _17;
    assign _884 = _880 ? _883 : _878;
    assign _885 = _884[62:0];
    assign _887 = { _885,
                    _886 };
    assign _888 = _887 < _17;
    assign _889 = ~ _888;
    assign _877 = _597[32:32];
    assign _874 = _869 - _17;
    assign _875 = _871 ? _874 : _869;
    assign _876 = _875[62:0];
    assign _878 = { _876,
                    _877 };
    assign _879 = _878 < _17;
    assign _880 = ~ _879;
    assign _868 = _597[33:33];
    assign _865 = _860 - _17;
    assign _866 = _862 ? _865 : _860;
    assign _867 = _866[62:0];
    assign _869 = { _867,
                    _868 };
    assign _870 = _869 < _17;
    assign _871 = ~ _870;
    assign _859 = _597[34:34];
    assign _856 = _851 - _17;
    assign _857 = _853 ? _856 : _851;
    assign _858 = _857[62:0];
    assign _860 = { _858,
                    _859 };
    assign _861 = _860 < _17;
    assign _862 = ~ _861;
    assign _850 = _597[35:35];
    assign _847 = _842 - _17;
    assign _848 = _844 ? _847 : _842;
    assign _849 = _848[62:0];
    assign _851 = { _849,
                    _850 };
    assign _852 = _851 < _17;
    assign _853 = ~ _852;
    assign _841 = _597[36:36];
    assign _838 = _833 - _17;
    assign _839 = _835 ? _838 : _833;
    assign _840 = _839[62:0];
    assign _842 = { _840,
                    _841 };
    assign _843 = _842 < _17;
    assign _844 = ~ _843;
    assign _832 = _597[37:37];
    assign _829 = _824 - _17;
    assign _830 = _826 ? _829 : _824;
    assign _831 = _830[62:0];
    assign _833 = { _831,
                    _832 };
    assign _834 = _833 < _17;
    assign _835 = ~ _834;
    assign _823 = _597[38:38];
    assign _820 = _815 - _17;
    assign _821 = _817 ? _820 : _815;
    assign _822 = _821[62:0];
    assign _824 = { _822,
                    _823 };
    assign _825 = _824 < _17;
    assign _826 = ~ _825;
    assign _814 = _597[39:39];
    assign _811 = _806 - _17;
    assign _812 = _808 ? _811 : _806;
    assign _813 = _812[62:0];
    assign _815 = { _813,
                    _814 };
    assign _816 = _815 < _17;
    assign _817 = ~ _816;
    assign _805 = _597[40:40];
    assign _802 = _797 - _17;
    assign _803 = _799 ? _802 : _797;
    assign _804 = _803[62:0];
    assign _806 = { _804,
                    _805 };
    assign _807 = _806 < _17;
    assign _808 = ~ _807;
    assign _796 = _597[41:41];
    assign _793 = _788 - _17;
    assign _794 = _790 ? _793 : _788;
    assign _795 = _794[62:0];
    assign _797 = { _795,
                    _796 };
    assign _798 = _797 < _17;
    assign _799 = ~ _798;
    assign _787 = _597[42:42];
    assign _784 = _779 - _17;
    assign _785 = _781 ? _784 : _779;
    assign _786 = _785[62:0];
    assign _788 = { _786,
                    _787 };
    assign _789 = _788 < _17;
    assign _790 = ~ _789;
    assign _778 = _597[43:43];
    assign _775 = _770 - _17;
    assign _776 = _772 ? _775 : _770;
    assign _777 = _776[62:0];
    assign _779 = { _777,
                    _778 };
    assign _780 = _779 < _17;
    assign _781 = ~ _780;
    assign _769 = _597[44:44];
    assign _766 = _761 - _17;
    assign _767 = _763 ? _766 : _761;
    assign _768 = _767[62:0];
    assign _770 = { _768,
                    _769 };
    assign _771 = _770 < _17;
    assign _772 = ~ _771;
    assign _760 = _597[45:45];
    assign _757 = _752 - _17;
    assign _758 = _754 ? _757 : _752;
    assign _759 = _758[62:0];
    assign _761 = { _759,
                    _760 };
    assign _762 = _761 < _17;
    assign _763 = ~ _762;
    assign _751 = _597[46:46];
    assign _748 = _743 - _17;
    assign _749 = _745 ? _748 : _743;
    assign _750 = _749[62:0];
    assign _752 = { _750,
                    _751 };
    assign _753 = _752 < _17;
    assign _754 = ~ _753;
    assign _742 = _597[47:47];
    assign _739 = _734 - _17;
    assign _740 = _736 ? _739 : _734;
    assign _741 = _740[62:0];
    assign _743 = { _741,
                    _742 };
    assign _744 = _743 < _17;
    assign _745 = ~ _744;
    assign _733 = _597[48:48];
    assign _730 = _725 - _17;
    assign _731 = _727 ? _730 : _725;
    assign _732 = _731[62:0];
    assign _734 = { _732,
                    _733 };
    assign _735 = _734 < _17;
    assign _736 = ~ _735;
    assign _724 = _597[49:49];
    assign _721 = _716 - _17;
    assign _722 = _718 ? _721 : _716;
    assign _723 = _722[62:0];
    assign _725 = { _723,
                    _724 };
    assign _726 = _725 < _17;
    assign _727 = ~ _726;
    assign _715 = _597[50:50];
    assign _712 = _707 - _17;
    assign _713 = _709 ? _712 : _707;
    assign _714 = _713[62:0];
    assign _716 = { _714,
                    _715 };
    assign _717 = _716 < _17;
    assign _718 = ~ _717;
    assign _706 = _597[51:51];
    assign _703 = _698 - _17;
    assign _704 = _700 ? _703 : _698;
    assign _705 = _704[62:0];
    assign _707 = { _705,
                    _706 };
    assign _708 = _707 < _17;
    assign _709 = ~ _708;
    assign _697 = _597[52:52];
    assign _694 = _689 - _17;
    assign _695 = _691 ? _694 : _689;
    assign _696 = _695[62:0];
    assign _698 = { _696,
                    _697 };
    assign _699 = _698 < _17;
    assign _700 = ~ _699;
    assign _688 = _597[53:53];
    assign _685 = _680 - _17;
    assign _686 = _682 ? _685 : _680;
    assign _687 = _686[62:0];
    assign _689 = { _687,
                    _688 };
    assign _690 = _689 < _17;
    assign _691 = ~ _690;
    assign _679 = _597[54:54];
    assign _676 = _671 - _17;
    assign _677 = _673 ? _676 : _671;
    assign _678 = _677[62:0];
    assign _680 = { _678,
                    _679 };
    assign _681 = _680 < _17;
    assign _682 = ~ _681;
    assign _670 = _597[55:55];
    assign _667 = _662 - _17;
    assign _668 = _664 ? _667 : _662;
    assign _669 = _668[62:0];
    assign _671 = { _669,
                    _670 };
    assign _672 = _671 < _17;
    assign _673 = ~ _672;
    assign _661 = _597[56:56];
    assign _658 = _653 - _17;
    assign _659 = _655 ? _658 : _653;
    assign _660 = _659[62:0];
    assign _662 = { _660,
                    _661 };
    assign _663 = _662 < _17;
    assign _664 = ~ _663;
    assign _652 = _597[57:57];
    assign _649 = _644 - _17;
    assign _650 = _646 ? _649 : _644;
    assign _651 = _650[62:0];
    assign _653 = { _651,
                    _652 };
    assign _654 = _653 < _17;
    assign _655 = ~ _654;
    assign _643 = _597[58:58];
    assign _640 = _635 - _17;
    assign _641 = _637 ? _640 : _635;
    assign _642 = _641[62:0];
    assign _644 = { _642,
                    _643 };
    assign _645 = _644 < _17;
    assign _646 = ~ _645;
    assign _634 = _597[59:59];
    assign _631 = _626 - _17;
    assign _632 = _628 ? _631 : _626;
    assign _633 = _632[62:0];
    assign _635 = { _633,
                    _634 };
    assign _636 = _635 < _17;
    assign _637 = ~ _636;
    assign _625 = _597[60:60];
    assign _622 = _617 - _17;
    assign _623 = _619 ? _622 : _617;
    assign _624 = _623[62:0];
    assign _626 = { _624,
                    _625 };
    assign _627 = _626 < _17;
    assign _628 = ~ _627;
    assign _616 = _597[61:61];
    assign _613 = _608 - _17;
    assign _614 = _610 ? _613 : _608;
    assign _615 = _614[62:0];
    assign _617 = { _615,
                    _616 };
    assign _618 = _617 < _17;
    assign _619 = ~ _618;
    assign _607 = _597[62:62];
    assign _604 = _599 - _17;
    assign _605 = _601 ? _604 : _599;
    assign _606 = _605[62:0];
    assign _608 = { _606,
                    _607 };
    assign _609 = _608 < _17;
    assign _610 = ~ _609;
    assign _597 = _9 - _591;
    assign _598 = _597[63:63];
    assign _599 = { _22185,
                    _598 };
    assign _600 = _599 < _17;
    assign _601 = ~ _600;
    assign _602 = { _22185,
                    _601 };
    assign _603 = _602[62:0];
    assign _611 = { _603,
                    _610 };
    assign _612 = _611[62:0];
    assign _620 = { _612,
                    _619 };
    assign _621 = _620[62:0];
    assign _629 = { _621,
                    _628 };
    assign _630 = _629[62:0];
    assign _638 = { _630,
                    _637 };
    assign _639 = _638[62:0];
    assign _647 = { _639,
                    _646 };
    assign _648 = _647[62:0];
    assign _656 = { _648,
                    _655 };
    assign _657 = _656[62:0];
    assign _665 = { _657,
                    _664 };
    assign _666 = _665[62:0];
    assign _674 = { _666,
                    _673 };
    assign _675 = _674[62:0];
    assign _683 = { _675,
                    _682 };
    assign _684 = _683[62:0];
    assign _692 = { _684,
                    _691 };
    assign _693 = _692[62:0];
    assign _701 = { _693,
                    _700 };
    assign _702 = _701[62:0];
    assign _710 = { _702,
                    _709 };
    assign _711 = _710[62:0];
    assign _719 = { _711,
                    _718 };
    assign _720 = _719[62:0];
    assign _728 = { _720,
                    _727 };
    assign _729 = _728[62:0];
    assign _737 = { _729,
                    _736 };
    assign _738 = _737[62:0];
    assign _746 = { _738,
                    _745 };
    assign _747 = _746[62:0];
    assign _755 = { _747,
                    _754 };
    assign _756 = _755[62:0];
    assign _764 = { _756,
                    _763 };
    assign _765 = _764[62:0];
    assign _773 = { _765,
                    _772 };
    assign _774 = _773[62:0];
    assign _782 = { _774,
                    _781 };
    assign _783 = _782[62:0];
    assign _791 = { _783,
                    _790 };
    assign _792 = _791[62:0];
    assign _800 = { _792,
                    _799 };
    assign _801 = _800[62:0];
    assign _809 = { _801,
                    _808 };
    assign _810 = _809[62:0];
    assign _818 = { _810,
                    _817 };
    assign _819 = _818[62:0];
    assign _827 = { _819,
                    _826 };
    assign _828 = _827[62:0];
    assign _836 = { _828,
                    _835 };
    assign _837 = _836[62:0];
    assign _845 = { _837,
                    _844 };
    assign _846 = _845[62:0];
    assign _854 = { _846,
                    _853 };
    assign _855 = _854[62:0];
    assign _863 = { _855,
                    _862 };
    assign _864 = _863[62:0];
    assign _872 = { _864,
                    _871 };
    assign _873 = _872[62:0];
    assign _881 = { _873,
                    _880 };
    assign _882 = _881[62:0];
    assign _890 = { _882,
                    _889 };
    assign _891 = _890[62:0];
    assign _899 = { _891,
                    _898 };
    assign _900 = _899[62:0];
    assign _908 = { _900,
                    _907 };
    assign _909 = _908[62:0];
    assign _917 = { _909,
                    _916 };
    assign _918 = _917[62:0];
    assign _926 = { _918,
                    _925 };
    assign _927 = _926[62:0];
    assign _935 = { _927,
                    _934 };
    assign _936 = _935[62:0];
    assign _944 = { _936,
                    _943 };
    assign _945 = _944[62:0];
    assign _953 = { _945,
                    _952 };
    assign _954 = _953[62:0];
    assign _962 = { _954,
                    _961 };
    assign _963 = _962[62:0];
    assign _971 = { _963,
                    _970 };
    assign _972 = _971[62:0];
    assign _980 = { _972,
                    _979 };
    assign _981 = _980[62:0];
    assign _989 = { _981,
                    _988 };
    assign _990 = _989[62:0];
    assign _998 = { _990,
                    _997 };
    assign _999 = _998[62:0];
    assign _1007 = { _999,
                     _1006 };
    assign _1008 = _1007[62:0];
    assign _1016 = { _1008,
                     _1015 };
    assign _1017 = _1016[62:0];
    assign _1025 = { _1017,
                     _1024 };
    assign _1026 = _1025[62:0];
    assign _1034 = { _1026,
                     _1033 };
    assign _1035 = _1034[62:0];
    assign _1043 = { _1035,
                     _1042 };
    assign _1044 = _1043[62:0];
    assign _1052 = { _1044,
                     _1051 };
    assign _1053 = _1052[62:0];
    assign _1061 = { _1053,
                     _1060 };
    assign _1062 = _1061[62:0];
    assign _1070 = { _1062,
                     _1069 };
    assign _1071 = _1070[62:0];
    assign _1079 = { _1071,
                     _1078 };
    assign _1080 = _1079[62:0];
    assign _1088 = { _1080,
                     _1087 };
    assign _1089 = _1088[62:0];
    assign _1097 = { _1089,
                     _1096 };
    assign _1098 = _1097[62:0];
    assign _1106 = { _1098,
                     _1105 };
    assign _1107 = _1106[62:0];
    assign _1115 = { _1107,
                     _1114 };
    assign _1116 = _1115[62:0];
    assign _1124 = { _1116,
                     _1123 };
    assign _1125 = _1124[62:0];
    assign _1133 = { _1125,
                     _1132 };
    assign _1134 = _1133[62:0];
    assign _1142 = { _1134,
                     _1141 };
    assign _1143 = _1142[62:0];
    assign _1151 = { _1143,
                     _1150 };
    assign _1152 = _1151[62:0];
    assign _1160 = { _1152,
                     _1159 };
    assign _1161 = _1160[62:0];
    assign _1169 = { _1161,
                     _1168 };
    assign _1171 = _1169 + _22186;
    assign _1172 = _1171 * _591;
    assign _1173 = _1172[63:0];
    assign _1755 = _1173 + _1754;
    assign _583 = _14[0:0];
    assign _580 = _575 - _17;
    assign _581 = _577 ? _580 : _575;
    assign _582 = _581[62:0];
    assign _584 = { _582,
                    _583 };
    assign _585 = _584 < _17;
    assign _586 = ~ _585;
    assign _574 = _14[1:1];
    assign _571 = _566 - _17;
    assign _572 = _568 ? _571 : _566;
    assign _573 = _572[62:0];
    assign _575 = { _573,
                    _574 };
    assign _576 = _575 < _17;
    assign _577 = ~ _576;
    assign _565 = _14[2:2];
    assign _562 = _557 - _17;
    assign _563 = _559 ? _562 : _557;
    assign _564 = _563[62:0];
    assign _566 = { _564,
                    _565 };
    assign _567 = _566 < _17;
    assign _568 = ~ _567;
    assign _556 = _14[3:3];
    assign _553 = _548 - _17;
    assign _554 = _550 ? _553 : _548;
    assign _555 = _554[62:0];
    assign _557 = { _555,
                    _556 };
    assign _558 = _557 < _17;
    assign _559 = ~ _558;
    assign _547 = _14[4:4];
    assign _544 = _539 - _17;
    assign _545 = _541 ? _544 : _539;
    assign _546 = _545[62:0];
    assign _548 = { _546,
                    _547 };
    assign _549 = _548 < _17;
    assign _550 = ~ _549;
    assign _538 = _14[5:5];
    assign _535 = _530 - _17;
    assign _536 = _532 ? _535 : _530;
    assign _537 = _536[62:0];
    assign _539 = { _537,
                    _538 };
    assign _540 = _539 < _17;
    assign _541 = ~ _540;
    assign _529 = _14[6:6];
    assign _526 = _521 - _17;
    assign _527 = _523 ? _526 : _521;
    assign _528 = _527[62:0];
    assign _530 = { _528,
                    _529 };
    assign _531 = _530 < _17;
    assign _532 = ~ _531;
    assign _520 = _14[7:7];
    assign _517 = _512 - _17;
    assign _518 = _514 ? _517 : _512;
    assign _519 = _518[62:0];
    assign _521 = { _519,
                    _520 };
    assign _522 = _521 < _17;
    assign _523 = ~ _522;
    assign _511 = _14[8:8];
    assign _508 = _503 - _17;
    assign _509 = _505 ? _508 : _503;
    assign _510 = _509[62:0];
    assign _512 = { _510,
                    _511 };
    assign _513 = _512 < _17;
    assign _514 = ~ _513;
    assign _502 = _14[9:9];
    assign _499 = _494 - _17;
    assign _500 = _496 ? _499 : _494;
    assign _501 = _500[62:0];
    assign _503 = { _501,
                    _502 };
    assign _504 = _503 < _17;
    assign _505 = ~ _504;
    assign _493 = _14[10:10];
    assign _490 = _485 - _17;
    assign _491 = _487 ? _490 : _485;
    assign _492 = _491[62:0];
    assign _494 = { _492,
                    _493 };
    assign _495 = _494 < _17;
    assign _496 = ~ _495;
    assign _484 = _14[11:11];
    assign _481 = _476 - _17;
    assign _482 = _478 ? _481 : _476;
    assign _483 = _482[62:0];
    assign _485 = { _483,
                    _484 };
    assign _486 = _485 < _17;
    assign _487 = ~ _486;
    assign _475 = _14[12:12];
    assign _472 = _467 - _17;
    assign _473 = _469 ? _472 : _467;
    assign _474 = _473[62:0];
    assign _476 = { _474,
                    _475 };
    assign _477 = _476 < _17;
    assign _478 = ~ _477;
    assign _466 = _14[13:13];
    assign _463 = _458 - _17;
    assign _464 = _460 ? _463 : _458;
    assign _465 = _464[62:0];
    assign _467 = { _465,
                    _466 };
    assign _468 = _467 < _17;
    assign _469 = ~ _468;
    assign _457 = _14[14:14];
    assign _454 = _449 - _17;
    assign _455 = _451 ? _454 : _449;
    assign _456 = _455[62:0];
    assign _458 = { _456,
                    _457 };
    assign _459 = _458 < _17;
    assign _460 = ~ _459;
    assign _448 = _14[15:15];
    assign _445 = _440 - _17;
    assign _446 = _442 ? _445 : _440;
    assign _447 = _446[62:0];
    assign _449 = { _447,
                    _448 };
    assign _450 = _449 < _17;
    assign _451 = ~ _450;
    assign _439 = _14[16:16];
    assign _436 = _431 - _17;
    assign _437 = _433 ? _436 : _431;
    assign _438 = _437[62:0];
    assign _440 = { _438,
                    _439 };
    assign _441 = _440 < _17;
    assign _442 = ~ _441;
    assign _430 = _14[17:17];
    assign _427 = _422 - _17;
    assign _428 = _424 ? _427 : _422;
    assign _429 = _428[62:0];
    assign _431 = { _429,
                    _430 };
    assign _432 = _431 < _17;
    assign _433 = ~ _432;
    assign _421 = _14[18:18];
    assign _418 = _413 - _17;
    assign _419 = _415 ? _418 : _413;
    assign _420 = _419[62:0];
    assign _422 = { _420,
                    _421 };
    assign _423 = _422 < _17;
    assign _424 = ~ _423;
    assign _412 = _14[19:19];
    assign _409 = _404 - _17;
    assign _410 = _406 ? _409 : _404;
    assign _411 = _410[62:0];
    assign _413 = { _411,
                    _412 };
    assign _414 = _413 < _17;
    assign _415 = ~ _414;
    assign _403 = _14[20:20];
    assign _400 = _395 - _17;
    assign _401 = _397 ? _400 : _395;
    assign _402 = _401[62:0];
    assign _404 = { _402,
                    _403 };
    assign _405 = _404 < _17;
    assign _406 = ~ _405;
    assign _394 = _14[21:21];
    assign _391 = _386 - _17;
    assign _392 = _388 ? _391 : _386;
    assign _393 = _392[62:0];
    assign _395 = { _393,
                    _394 };
    assign _396 = _395 < _17;
    assign _397 = ~ _396;
    assign _385 = _14[22:22];
    assign _382 = _377 - _17;
    assign _383 = _379 ? _382 : _377;
    assign _384 = _383[62:0];
    assign _386 = { _384,
                    _385 };
    assign _387 = _386 < _17;
    assign _388 = ~ _387;
    assign _376 = _14[23:23];
    assign _373 = _368 - _17;
    assign _374 = _370 ? _373 : _368;
    assign _375 = _374[62:0];
    assign _377 = { _375,
                    _376 };
    assign _378 = _377 < _17;
    assign _379 = ~ _378;
    assign _367 = _14[24:24];
    assign _364 = _359 - _17;
    assign _365 = _361 ? _364 : _359;
    assign _366 = _365[62:0];
    assign _368 = { _366,
                    _367 };
    assign _369 = _368 < _17;
    assign _370 = ~ _369;
    assign _358 = _14[25:25];
    assign _355 = _350 - _17;
    assign _356 = _352 ? _355 : _350;
    assign _357 = _356[62:0];
    assign _359 = { _357,
                    _358 };
    assign _360 = _359 < _17;
    assign _361 = ~ _360;
    assign _349 = _14[26:26];
    assign _346 = _341 - _17;
    assign _347 = _343 ? _346 : _341;
    assign _348 = _347[62:0];
    assign _350 = { _348,
                    _349 };
    assign _351 = _350 < _17;
    assign _352 = ~ _351;
    assign _340 = _14[27:27];
    assign _337 = _332 - _17;
    assign _338 = _334 ? _337 : _332;
    assign _339 = _338[62:0];
    assign _341 = { _339,
                    _340 };
    assign _342 = _341 < _17;
    assign _343 = ~ _342;
    assign _331 = _14[28:28];
    assign _328 = _323 - _17;
    assign _329 = _325 ? _328 : _323;
    assign _330 = _329[62:0];
    assign _332 = { _330,
                    _331 };
    assign _333 = _332 < _17;
    assign _334 = ~ _333;
    assign _322 = _14[29:29];
    assign _319 = _314 - _17;
    assign _320 = _316 ? _319 : _314;
    assign _321 = _320[62:0];
    assign _323 = { _321,
                    _322 };
    assign _324 = _323 < _17;
    assign _325 = ~ _324;
    assign _313 = _14[30:30];
    assign _310 = _305 - _17;
    assign _311 = _307 ? _310 : _305;
    assign _312 = _311[62:0];
    assign _314 = { _312,
                    _313 };
    assign _315 = _314 < _17;
    assign _316 = ~ _315;
    assign _304 = _14[31:31];
    assign _301 = _296 - _17;
    assign _302 = _298 ? _301 : _296;
    assign _303 = _302[62:0];
    assign _305 = { _303,
                    _304 };
    assign _306 = _305 < _17;
    assign _307 = ~ _306;
    assign _295 = _14[32:32];
    assign _292 = _287 - _17;
    assign _293 = _289 ? _292 : _287;
    assign _294 = _293[62:0];
    assign _296 = { _294,
                    _295 };
    assign _297 = _296 < _17;
    assign _298 = ~ _297;
    assign _286 = _14[33:33];
    assign _283 = _278 - _17;
    assign _284 = _280 ? _283 : _278;
    assign _285 = _284[62:0];
    assign _287 = { _285,
                    _286 };
    assign _288 = _287 < _17;
    assign _289 = ~ _288;
    assign _277 = _14[34:34];
    assign _274 = _269 - _17;
    assign _275 = _271 ? _274 : _269;
    assign _276 = _275[62:0];
    assign _278 = { _276,
                    _277 };
    assign _279 = _278 < _17;
    assign _280 = ~ _279;
    assign _268 = _14[35:35];
    assign _265 = _260 - _17;
    assign _266 = _262 ? _265 : _260;
    assign _267 = _266[62:0];
    assign _269 = { _267,
                    _268 };
    assign _270 = _269 < _17;
    assign _271 = ~ _270;
    assign _259 = _14[36:36];
    assign _256 = _251 - _17;
    assign _257 = _253 ? _256 : _251;
    assign _258 = _257[62:0];
    assign _260 = { _258,
                    _259 };
    assign _261 = _260 < _17;
    assign _262 = ~ _261;
    assign _250 = _14[37:37];
    assign _247 = _242 - _17;
    assign _248 = _244 ? _247 : _242;
    assign _249 = _248[62:0];
    assign _251 = { _249,
                    _250 };
    assign _252 = _251 < _17;
    assign _253 = ~ _252;
    assign _241 = _14[38:38];
    assign _238 = _233 - _17;
    assign _239 = _235 ? _238 : _233;
    assign _240 = _239[62:0];
    assign _242 = { _240,
                    _241 };
    assign _243 = _242 < _17;
    assign _244 = ~ _243;
    assign _232 = _14[39:39];
    assign _229 = _224 - _17;
    assign _230 = _226 ? _229 : _224;
    assign _231 = _230[62:0];
    assign _233 = { _231,
                    _232 };
    assign _234 = _233 < _17;
    assign _235 = ~ _234;
    assign _223 = _14[40:40];
    assign _220 = _215 - _17;
    assign _221 = _217 ? _220 : _215;
    assign _222 = _221[62:0];
    assign _224 = { _222,
                    _223 };
    assign _225 = _224 < _17;
    assign _226 = ~ _225;
    assign _214 = _14[41:41];
    assign _211 = _206 - _17;
    assign _212 = _208 ? _211 : _206;
    assign _213 = _212[62:0];
    assign _215 = { _213,
                    _214 };
    assign _216 = _215 < _17;
    assign _217 = ~ _216;
    assign _205 = _14[42:42];
    assign _202 = _197 - _17;
    assign _203 = _199 ? _202 : _197;
    assign _204 = _203[62:0];
    assign _206 = { _204,
                    _205 };
    assign _207 = _206 < _17;
    assign _208 = ~ _207;
    assign _196 = _14[43:43];
    assign _193 = _188 - _17;
    assign _194 = _190 ? _193 : _188;
    assign _195 = _194[62:0];
    assign _197 = { _195,
                    _196 };
    assign _198 = _197 < _17;
    assign _199 = ~ _198;
    assign _187 = _14[44:44];
    assign _184 = _179 - _17;
    assign _185 = _181 ? _184 : _179;
    assign _186 = _185[62:0];
    assign _188 = { _186,
                    _187 };
    assign _189 = _188 < _17;
    assign _190 = ~ _189;
    assign _178 = _14[45:45];
    assign _175 = _170 - _17;
    assign _176 = _172 ? _175 : _170;
    assign _177 = _176[62:0];
    assign _179 = { _177,
                    _178 };
    assign _180 = _179 < _17;
    assign _181 = ~ _180;
    assign _169 = _14[46:46];
    assign _166 = _161 - _17;
    assign _167 = _163 ? _166 : _161;
    assign _168 = _167[62:0];
    assign _170 = { _168,
                    _169 };
    assign _171 = _170 < _17;
    assign _172 = ~ _171;
    assign _160 = _14[47:47];
    assign _157 = _152 - _17;
    assign _158 = _154 ? _157 : _152;
    assign _159 = _158[62:0];
    assign _161 = { _159,
                    _160 };
    assign _162 = _161 < _17;
    assign _163 = ~ _162;
    assign _151 = _14[48:48];
    assign _148 = _143 - _17;
    assign _149 = _145 ? _148 : _143;
    assign _150 = _149[62:0];
    assign _152 = { _150,
                    _151 };
    assign _153 = _152 < _17;
    assign _154 = ~ _153;
    assign _142 = _14[49:49];
    assign _139 = _134 - _17;
    assign _140 = _136 ? _139 : _134;
    assign _141 = _140[62:0];
    assign _143 = { _141,
                    _142 };
    assign _144 = _143 < _17;
    assign _145 = ~ _144;
    assign _133 = _14[50:50];
    assign _130 = _125 - _17;
    assign _131 = _127 ? _130 : _125;
    assign _132 = _131[62:0];
    assign _134 = { _132,
                    _133 };
    assign _135 = _134 < _17;
    assign _136 = ~ _135;
    assign _124 = _14[51:51];
    assign _121 = _116 - _17;
    assign _122 = _118 ? _121 : _116;
    assign _123 = _122[62:0];
    assign _125 = { _123,
                    _124 };
    assign _126 = _125 < _17;
    assign _127 = ~ _126;
    assign _115 = _14[52:52];
    assign _112 = _107 - _17;
    assign _113 = _109 ? _112 : _107;
    assign _114 = _113[62:0];
    assign _116 = { _114,
                    _115 };
    assign _117 = _116 < _17;
    assign _118 = ~ _117;
    assign _106 = _14[53:53];
    assign _103 = _98 - _17;
    assign _104 = _100 ? _103 : _98;
    assign _105 = _104[62:0];
    assign _107 = { _105,
                    _106 };
    assign _108 = _107 < _17;
    assign _109 = ~ _108;
    assign _97 = _14[54:54];
    assign _94 = _89 - _17;
    assign _95 = _91 ? _94 : _89;
    assign _96 = _95[62:0];
    assign _98 = { _96,
                   _97 };
    assign _99 = _98 < _17;
    assign _100 = ~ _99;
    assign _88 = _14[55:55];
    assign _85 = _80 - _17;
    assign _86 = _82 ? _85 : _80;
    assign _87 = _86[62:0];
    assign _89 = { _87,
                   _88 };
    assign _90 = _89 < _17;
    assign _91 = ~ _90;
    assign _79 = _14[56:56];
    assign _76 = _71 - _17;
    assign _77 = _73 ? _76 : _71;
    assign _78 = _77[62:0];
    assign _80 = { _78,
                   _79 };
    assign _81 = _80 < _17;
    assign _82 = ~ _81;
    assign _70 = _14[57:57];
    assign _67 = _62 - _17;
    assign _68 = _64 ? _67 : _62;
    assign _69 = _68[62:0];
    assign _71 = { _69,
                   _70 };
    assign _72 = _71 < _17;
    assign _73 = ~ _72;
    assign _61 = _14[58:58];
    assign _58 = _53 - _17;
    assign _59 = _55 ? _58 : _53;
    assign _60 = _59[62:0];
    assign _62 = { _60,
                   _61 };
    assign _63 = _62 < _17;
    assign _64 = ~ _63;
    assign _52 = _14[59:59];
    assign _49 = _44 - _17;
    assign _50 = _46 ? _49 : _44;
    assign _51 = _50[62:0];
    assign _53 = { _51,
                   _52 };
    assign _54 = _53 < _17;
    assign _55 = ~ _54;
    assign _43 = _14[60:60];
    assign _40 = _35 - _17;
    assign _41 = _37 ? _40 : _35;
    assign _42 = _41[62:0];
    assign _44 = { _42,
                   _43 };
    assign _45 = _44 < _17;
    assign _46 = ~ _45;
    assign _34 = _14[61:61];
    assign _31 = _26 - _17;
    assign _32 = _28 ? _31 : _26;
    assign _33 = _32[62:0];
    assign _35 = { _33,
                   _34 };
    assign _36 = _35 < _17;
    assign _37 = ~ _36;
    assign _25 = _14[62:62];
    assign _22 = _16 - _17;
    assign _23 = _19 ? _22 : _16;
    assign _24 = _23[62:0];
    assign _26 = { _24,
                   _25 };
    assign _27 = _26 < _17;
    assign _28 = ~ _27;
    assign _17 = 64'b0000000000000000000000000000000000000000000000000000000000001011;
    assign _13 = 64'b0000000000000000000000000000000000000000000000000000000000001010;
    assign _3 = from_;
    assign _14 = _3 + _13;
    assign _15 = _14[63:63];
    assign _16 = { _22185,
                   _15 };
    assign _18 = _16 < _17;
    assign _19 = ~ _18;
    assign _20 = { _22185,
                   _19 };
    assign _21 = _20[62:0];
    assign _29 = { _21,
                   _28 };
    assign _30 = _29[62:0];
    assign _38 = { _30,
                   _37 };
    assign _39 = _38[62:0];
    assign _47 = { _39,
                   _46 };
    assign _48 = _47[62:0];
    assign _56 = { _48,
                   _55 };
    assign _57 = _56[62:0];
    assign _65 = { _57,
                   _64 };
    assign _66 = _65[62:0];
    assign _74 = { _66,
                   _73 };
    assign _75 = _74[62:0];
    assign _83 = { _75,
                   _82 };
    assign _84 = _83[62:0];
    assign _92 = { _84,
                   _91 };
    assign _93 = _92[62:0];
    assign _101 = { _93,
                    _100 };
    assign _102 = _101[62:0];
    assign _110 = { _102,
                    _109 };
    assign _111 = _110[62:0];
    assign _119 = { _111,
                    _118 };
    assign _120 = _119[62:0];
    assign _128 = { _120,
                    _127 };
    assign _129 = _128[62:0];
    assign _137 = { _129,
                    _136 };
    assign _138 = _137[62:0];
    assign _146 = { _138,
                    _145 };
    assign _147 = _146[62:0];
    assign _155 = { _147,
                    _154 };
    assign _156 = _155[62:0];
    assign _164 = { _156,
                    _163 };
    assign _165 = _164[62:0];
    assign _173 = { _165,
                    _172 };
    assign _174 = _173[62:0];
    assign _182 = { _174,
                    _181 };
    assign _183 = _182[62:0];
    assign _191 = { _183,
                    _190 };
    assign _192 = _191[62:0];
    assign _200 = { _192,
                    _199 };
    assign _201 = _200[62:0];
    assign _209 = { _201,
                    _208 };
    assign _210 = _209[62:0];
    assign _218 = { _210,
                    _217 };
    assign _219 = _218[62:0];
    assign _227 = { _219,
                    _226 };
    assign _228 = _227[62:0];
    assign _236 = { _228,
                    _235 };
    assign _237 = _236[62:0];
    assign _245 = { _237,
                    _244 };
    assign _246 = _245[62:0];
    assign _254 = { _246,
                    _253 };
    assign _255 = _254[62:0];
    assign _263 = { _255,
                    _262 };
    assign _264 = _263[62:0];
    assign _272 = { _264,
                    _271 };
    assign _273 = _272[62:0];
    assign _281 = { _273,
                    _280 };
    assign _282 = _281[62:0];
    assign _290 = { _282,
                    _289 };
    assign _291 = _290[62:0];
    assign _299 = { _291,
                    _298 };
    assign _300 = _299[62:0];
    assign _308 = { _300,
                    _307 };
    assign _309 = _308[62:0];
    assign _317 = { _309,
                    _316 };
    assign _318 = _317[62:0];
    assign _326 = { _318,
                    _325 };
    assign _327 = _326[62:0];
    assign _335 = { _327,
                    _334 };
    assign _336 = _335[62:0];
    assign _344 = { _336,
                    _343 };
    assign _345 = _344[62:0];
    assign _353 = { _345,
                    _352 };
    assign _354 = _353[62:0];
    assign _362 = { _354,
                    _361 };
    assign _363 = _362[62:0];
    assign _371 = { _363,
                    _370 };
    assign _372 = _371[62:0];
    assign _380 = { _372,
                    _379 };
    assign _381 = _380[62:0];
    assign _389 = { _381,
                    _388 };
    assign _390 = _389[62:0];
    assign _398 = { _390,
                    _397 };
    assign _399 = _398[62:0];
    assign _407 = { _399,
                    _406 };
    assign _408 = _407[62:0];
    assign _416 = { _408,
                    _415 };
    assign _417 = _416[62:0];
    assign _425 = { _417,
                    _424 };
    assign _426 = _425[62:0];
    assign _434 = { _426,
                    _433 };
    assign _435 = _434[62:0];
    assign _443 = { _435,
                    _442 };
    assign _444 = _443[62:0];
    assign _452 = { _444,
                    _451 };
    assign _453 = _452[62:0];
    assign _461 = { _453,
                    _460 };
    assign _462 = _461[62:0];
    assign _470 = { _462,
                    _469 };
    assign _471 = _470[62:0];
    assign _479 = { _471,
                    _478 };
    assign _480 = _479[62:0];
    assign _488 = { _480,
                    _487 };
    assign _489 = _488[62:0];
    assign _497 = { _489,
                    _496 };
    assign _498 = _497[62:0];
    assign _506 = { _498,
                    _505 };
    assign _507 = _506[62:0];
    assign _515 = { _507,
                    _514 };
    assign _516 = _515[62:0];
    assign _524 = { _516,
                    _523 };
    assign _525 = _524[62:0];
    assign _533 = { _525,
                    _532 };
    assign _534 = _533[62:0];
    assign _542 = { _534,
                    _541 };
    assign _543 = _542[62:0];
    assign _551 = { _543,
                    _550 };
    assign _552 = _551[62:0];
    assign _560 = { _552,
                    _559 };
    assign _561 = _560[62:0];
    assign _569 = { _561,
                    _568 };
    assign _570 = _569[62:0];
    assign _578 = { _570,
                    _577 };
    assign _579 = _578[62:0];
    assign _587 = { _579,
                    _586 };
    assign _588 = _587 * _17;
    assign _589 = _588[63:0];
    assign _590 = _17 < _589;
    assign _591 = _590 ? _589 : _17;
    assign _7 = 64'b0000000000000000000000000000000000000000000000000000000001100011;
    assign _5 = to_;
    assign _8 = _5 < _7;
    assign _9 = _8 ? _5 : _7;
    assign _592 = _9 < _591;
    assign _593 = ~ _592;
    assign _1756 = _593 ? _1755 : _21604;
    assign _3507 = _1756 + _3506;
    assign _5258 = _3507 + _5257;
    assign _7009 = _5258 + _7008;
    assign _8760 = _7009 + _8759;
    assign sum_p1 = _8760;
    assign sum_p2 = _22768;

endmodule
