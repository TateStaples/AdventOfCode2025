module day3 (
    data,
    start,
    clear,
    clock,
    k,
    length,
    result,
    done_
);

    input [511:0] data;
    input start;
    input clear;
    input clock;
    input [3:0] k;
    input [7:0] length;
    output [63:0] result;
    output done_;

    wire _42;
    wire _45;
    wire _46;
    wire _1;
    reg _43;
    wire [3:0] _50;
    wire [3:0] _331;
    wire _332;
    wire _333;
    wire [3:0] _328;
    wire _329;
    wire _327;
    wire _330;
    wire _334;
    wire [3:0] _335;
    wire [7:0] _58;
    wire [7:0] _59;
    reg [3:0] _188;
    wire _53;
    wire [3:0] _189;
    wire [3:0] _190;
    wire [3:0] _336;
    wire [3:0] _3;
    reg [3:0] _51;
    wire [59:0] _565;
    wire [63:0] _566;
    wire [63:0] _562;
    wire [127:0] _563;
    wire [63:0] _564;
    wire [63:0] _567;
    wire [3:0] _320;
    wire _324;
    wire _325;
    wire [3:0] _191;
    wire _195;
    wire _318;
    wire _319;
    wire _326;
    wire [3:0] _345;
    wire [7:0] _340;
    wire [7:0] _341;
    reg [3:0] _342;
    wire _338;
    wire [3:0] _343;
    wire [3:0] _344;
    wire [3:0] _346;
    wire [3:0] _4;
    reg [3:0] _323;
    wire [63:0] _559;
    wire [127:0] _556;
    wire [63:0] _557;
    wire [63:0] _560;
    wire [3:0] _311;
    wire _315;
    wire _316;
    wire [3:0] _197;
    wire _198;
    wire _309;
    wire _310;
    wire _317;
    wire [3:0] _355;
    wire [7:0] _350;
    wire [7:0] _351;
    reg [3:0] _352;
    wire _348;
    wire [3:0] _353;
    wire [3:0] _354;
    wire [3:0] _356;
    wire [3:0] _5;
    reg [3:0] _314;
    wire [63:0] _552;
    wire [127:0] _549;
    wire [63:0] _550;
    wire [63:0] _553;
    wire [3:0] _302;
    wire _306;
    wire _307;
    wire [3:0] _200;
    wire _201;
    wire _300;
    wire _301;
    wire _308;
    wire [3:0] _365;
    wire [7:0] _360;
    wire [7:0] _361;
    reg [3:0] _362;
    wire _358;
    wire [3:0] _363;
    wire [3:0] _364;
    wire [3:0] _366;
    wire [3:0] _6;
    reg [3:0] _305;
    wire [63:0] _545;
    wire [127:0] _542;
    wire [63:0] _543;
    wire [63:0] _546;
    wire [3:0] _293;
    wire _297;
    wire _298;
    wire [3:0] _203;
    wire _204;
    wire _291;
    wire _292;
    wire _299;
    wire [3:0] _375;
    wire [7:0] _370;
    wire [7:0] _371;
    reg [3:0] _372;
    wire _368;
    wire [3:0] _373;
    wire [3:0] _374;
    wire [3:0] _376;
    wire [3:0] _7;
    reg [3:0] _296;
    wire [63:0] _538;
    wire [127:0] _535;
    wire [63:0] _536;
    wire [63:0] _539;
    wire [3:0] _284;
    wire _288;
    wire _289;
    wire [3:0] _206;
    wire _207;
    wire _282;
    wire _283;
    wire _290;
    wire [3:0] _385;
    wire [7:0] _380;
    wire [7:0] _381;
    reg [3:0] _382;
    wire _378;
    wire [3:0] _383;
    wire [3:0] _384;
    wire [3:0] _386;
    wire [3:0] _8;
    reg [3:0] _287;
    wire [63:0] _531;
    wire [127:0] _528;
    wire [63:0] _529;
    wire [63:0] _532;
    wire [3:0] _275;
    wire _279;
    wire _280;
    wire [3:0] _209;
    wire _210;
    wire _273;
    wire _274;
    wire _281;
    wire [3:0] _395;
    wire [7:0] _390;
    wire [7:0] _391;
    reg [3:0] _392;
    wire _388;
    wire [3:0] _393;
    wire [3:0] _394;
    wire [3:0] _396;
    wire [3:0] _9;
    reg [3:0] _278;
    wire [63:0] _524;
    wire [127:0] _521;
    wire [63:0] _522;
    wire [63:0] _525;
    wire [3:0] _266;
    wire _270;
    wire _271;
    wire [3:0] _212;
    wire _213;
    wire _264;
    wire _265;
    wire _272;
    wire [3:0] _405;
    wire [7:0] _400;
    wire [7:0] _401;
    reg [3:0] _402;
    wire _398;
    wire [3:0] _403;
    wire [3:0] _404;
    wire [3:0] _406;
    wire [3:0] _10;
    reg [3:0] _269;
    wire [63:0] _517;
    wire [127:0] _514;
    wire [63:0] _515;
    wire [63:0] _518;
    wire [3:0] _257;
    wire _261;
    wire _262;
    wire [3:0] _215;
    wire _216;
    wire _255;
    wire _256;
    wire _263;
    wire [3:0] _415;
    wire [7:0] _410;
    wire [7:0] _411;
    reg [3:0] _412;
    wire _408;
    wire [3:0] _413;
    wire [3:0] _414;
    wire [3:0] _416;
    wire [3:0] _11;
    reg [3:0] _260;
    wire [63:0] _510;
    wire [127:0] _507;
    wire [63:0] _508;
    wire [63:0] _511;
    wire [3:0] _248;
    wire _252;
    wire _253;
    wire [3:0] _218;
    wire _219;
    wire _246;
    wire _247;
    wire _254;
    wire [3:0] _425;
    wire [7:0] _420;
    wire [7:0] _421;
    reg [3:0] _422;
    wire _418;
    wire [3:0] _423;
    wire [3:0] _424;
    wire [3:0] _426;
    wire [3:0] _12;
    reg [3:0] _251;
    wire [63:0] _503;
    wire [127:0] _500;
    wire [63:0] _501;
    wire [63:0] _504;
    wire [3:0] _239;
    wire _243;
    wire _244;
    wire [3:0] _221;
    wire _222;
    wire _237;
    wire _238;
    wire _245;
    wire [3:0] _435;
    wire [7:0] _430;
    wire [7:0] _431;
    reg [3:0] _432;
    wire _428;
    wire [3:0] _433;
    wire [3:0] _434;
    wire [3:0] _436;
    wire [3:0] _13;
    reg [3:0] _242;
    wire [63:0] _496;
    wire [127:0] _493;
    wire [63:0] _494;
    wire [63:0] _497;
    reg [3:0] _230;
    wire _234;
    wire _235;
    wire _225;
    wire _236;
    wire [3:0] _443;
    wire [3:0] _187;
    wire [3:0] _186;
    wire [3:0] _185;
    wire [3:0] _184;
    wire [3:0] _183;
    wire [3:0] _182;
    wire [3:0] _181;
    wire [3:0] _180;
    wire [3:0] _179;
    wire [3:0] _178;
    wire [3:0] _177;
    wire [3:0] _176;
    wire [3:0] _175;
    wire [3:0] _174;
    wire [3:0] _173;
    wire [3:0] _172;
    wire [3:0] _171;
    wire [3:0] _170;
    wire [3:0] _169;
    wire [3:0] _168;
    wire [3:0] _167;
    wire [3:0] _166;
    wire [3:0] _165;
    wire [3:0] _164;
    wire [3:0] _163;
    wire [3:0] _162;
    wire [3:0] _161;
    wire [3:0] _160;
    wire [3:0] _159;
    wire [3:0] _158;
    wire [3:0] _157;
    wire [3:0] _156;
    wire [3:0] _155;
    wire [3:0] _154;
    wire [3:0] _153;
    wire [3:0] _152;
    wire [3:0] _151;
    wire [3:0] _150;
    wire [3:0] _149;
    wire [3:0] _148;
    wire [3:0] _147;
    wire [3:0] _146;
    wire [3:0] _145;
    wire [3:0] _144;
    wire [3:0] _143;
    wire [3:0] _142;
    wire [3:0] _141;
    wire [3:0] _140;
    wire [3:0] _139;
    wire [3:0] _138;
    wire [3:0] _137;
    wire [3:0] _136;
    wire [3:0] _135;
    wire [3:0] _134;
    wire [3:0] _133;
    wire [3:0] _132;
    wire [3:0] _131;
    wire [3:0] _130;
    wire [3:0] _129;
    wire [3:0] _128;
    wire [3:0] _127;
    wire [3:0] _126;
    wire [3:0] _125;
    wire [3:0] _124;
    wire [3:0] _123;
    wire [3:0] _122;
    wire [3:0] _121;
    wire [3:0] _120;
    wire [3:0] _119;
    wire [3:0] _118;
    wire [3:0] _117;
    wire [3:0] _116;
    wire [3:0] _115;
    wire [3:0] _114;
    wire [3:0] _113;
    wire [3:0] _112;
    wire [3:0] _111;
    wire [3:0] _110;
    wire [3:0] _109;
    wire [3:0] _108;
    wire [3:0] _107;
    wire [3:0] _106;
    wire [3:0] _105;
    wire [3:0] _104;
    wire [3:0] _103;
    wire [3:0] _102;
    wire [3:0] _101;
    wire [3:0] _100;
    wire [3:0] _99;
    wire [3:0] _98;
    wire [3:0] _97;
    wire [3:0] _96;
    wire [3:0] _95;
    wire [3:0] _94;
    wire [3:0] _93;
    wire [3:0] _92;
    wire [3:0] _91;
    wire [3:0] _90;
    wire [3:0] _89;
    wire [3:0] _88;
    wire [3:0] _87;
    wire [3:0] _86;
    wire [3:0] _85;
    wire [3:0] _84;
    wire [3:0] _83;
    wire [3:0] _82;
    wire [3:0] _81;
    wire [3:0] _80;
    wire [3:0] _79;
    wire [3:0] _78;
    wire [3:0] _77;
    wire [3:0] _76;
    wire [3:0] _75;
    wire [3:0] _74;
    wire [3:0] _73;
    wire [3:0] _72;
    wire [3:0] _71;
    wire [3:0] _70;
    wire [3:0] _69;
    wire [3:0] _68;
    wire [3:0] _67;
    wire [3:0] _66;
    wire [3:0] _65;
    wire [3:0] _64;
    wire [3:0] _63;
    wire [3:0] _62;
    wire [3:0] _61;
    wire [511:0] _15;
    wire [3:0] _60;
    reg [3:0] _440;
    wire _438;
    wire [3:0] _441;
    wire [3:0] _442;
    wire [3:0] _444;
    wire [3:0] _16;
    reg [3:0] _233;
    wire [63:0] _490;
    wire [63:0] _488;
    wire _487;
    wire [63:0] _491;
    wire _485;
    wire [63:0] _498;
    wire _483;
    wire [63:0] _505;
    wire _481;
    wire [63:0] _512;
    wire _479;
    wire [63:0] _519;
    wire _477;
    wire [63:0] _526;
    wire _475;
    wire [63:0] _533;
    wire _473;
    wire [63:0] _540;
    wire _471;
    wire [63:0] _547;
    wire _469;
    wire [63:0] _554;
    wire _467;
    wire [63:0] _561;
    wire _18;
    wire [1:0] _35;
    wire _36;
    wire [1:0] _37;
    wire [1:0] _459;
    wire [7:0] _457;
    wire vdd;
    wire _20;
    wire _22;
    wire [7:0] _449;
    wire [7:0] _446;
    wire [7:0] _447;
    wire [7:0] _450;
    wire [7:0] _23;
    reg [7:0] _229;
    wire _458;
    wire [1:0] _461;
    wire [3:0] _25;
    wire [7:0] _56;
    wire [7:0] _27;
    wire [7:0] _57;
    wire _452;
    wire [1:0] _455;
    wire [1:0] _456;
    wire _48;
    wire [1:0] _462;
    wire [1:0] _28;
    reg [1:0] _34;
    wire _38;
    wire _39;
    wire _40;
    wire [3:0] _463;
    wire [3:0] _29;
    reg [3:0] _194;
    wire _465;
    wire [63:0] _568;
    assign _42 = 1'b0;
    assign _45 = _40 ? _42 : _43;
    assign _46 = _36 ? vdd : _45;
    assign _1 = _46;
    always @(posedge _22) begin
        if (_20)
            _43 <= _42;
        else
            _43 <= _1;
    end
    assign _50 = 4'b0000;
    assign _331 = _326 ? _323 : _320;
    assign _332 = _331 < _51;
    assign _333 = ~ _332;
    assign _328 = 4'b1011;
    assign _329 = _328 < _194;
    assign _327 = _195 ? _326 : _42;
    assign _330 = _327 & _329;
    assign _334 = _330 & _333;
    assign _335 = _334 ? _331 : _51;
    assign _58 = 8'b00001011;
    assign _59 = _57 + _58;
    always @* begin
        case (_59)
        0:
            _188 <= _60;
        1:
            _188 <= _61;
        2:
            _188 <= _62;
        3:
            _188 <= _63;
        4:
            _188 <= _64;
        5:
            _188 <= _65;
        6:
            _188 <= _66;
        7:
            _188 <= _67;
        8:
            _188 <= _68;
        9:
            _188 <= _69;
        10:
            _188 <= _70;
        11:
            _188 <= _71;
        12:
            _188 <= _72;
        13:
            _188 <= _73;
        14:
            _188 <= _74;
        15:
            _188 <= _75;
        16:
            _188 <= _76;
        17:
            _188 <= _77;
        18:
            _188 <= _78;
        19:
            _188 <= _79;
        20:
            _188 <= _80;
        21:
            _188 <= _81;
        22:
            _188 <= _82;
        23:
            _188 <= _83;
        24:
            _188 <= _84;
        25:
            _188 <= _85;
        26:
            _188 <= _86;
        27:
            _188 <= _87;
        28:
            _188 <= _88;
        29:
            _188 <= _89;
        30:
            _188 <= _90;
        31:
            _188 <= _91;
        32:
            _188 <= _92;
        33:
            _188 <= _93;
        34:
            _188 <= _94;
        35:
            _188 <= _95;
        36:
            _188 <= _96;
        37:
            _188 <= _97;
        38:
            _188 <= _98;
        39:
            _188 <= _99;
        40:
            _188 <= _100;
        41:
            _188 <= _101;
        42:
            _188 <= _102;
        43:
            _188 <= _103;
        44:
            _188 <= _104;
        45:
            _188 <= _105;
        46:
            _188 <= _106;
        47:
            _188 <= _107;
        48:
            _188 <= _108;
        49:
            _188 <= _109;
        50:
            _188 <= _110;
        51:
            _188 <= _111;
        52:
            _188 <= _112;
        53:
            _188 <= _113;
        54:
            _188 <= _114;
        55:
            _188 <= _115;
        56:
            _188 <= _116;
        57:
            _188 <= _117;
        58:
            _188 <= _118;
        59:
            _188 <= _119;
        60:
            _188 <= _120;
        61:
            _188 <= _121;
        62:
            _188 <= _122;
        63:
            _188 <= _123;
        64:
            _188 <= _124;
        65:
            _188 <= _125;
        66:
            _188 <= _126;
        67:
            _188 <= _127;
        68:
            _188 <= _128;
        69:
            _188 <= _129;
        70:
            _188 <= _130;
        71:
            _188 <= _131;
        72:
            _188 <= _132;
        73:
            _188 <= _133;
        74:
            _188 <= _134;
        75:
            _188 <= _135;
        76:
            _188 <= _136;
        77:
            _188 <= _137;
        78:
            _188 <= _138;
        79:
            _188 <= _139;
        80:
            _188 <= _140;
        81:
            _188 <= _141;
        82:
            _188 <= _142;
        83:
            _188 <= _143;
        84:
            _188 <= _144;
        85:
            _188 <= _145;
        86:
            _188 <= _146;
        87:
            _188 <= _147;
        88:
            _188 <= _148;
        89:
            _188 <= _149;
        90:
            _188 <= _150;
        91:
            _188 <= _151;
        92:
            _188 <= _152;
        93:
            _188 <= _153;
        94:
            _188 <= _154;
        95:
            _188 <= _155;
        96:
            _188 <= _156;
        97:
            _188 <= _157;
        98:
            _188 <= _158;
        99:
            _188 <= _159;
        100:
            _188 <= _160;
        101:
            _188 <= _161;
        102:
            _188 <= _162;
        103:
            _188 <= _163;
        104:
            _188 <= _164;
        105:
            _188 <= _165;
        106:
            _188 <= _166;
        107:
            _188 <= _167;
        108:
            _188 <= _168;
        109:
            _188 <= _169;
        110:
            _188 <= _170;
        111:
            _188 <= _171;
        112:
            _188 <= _172;
        113:
            _188 <= _173;
        114:
            _188 <= _174;
        115:
            _188 <= _175;
        116:
            _188 <= _176;
        117:
            _188 <= _177;
        118:
            _188 <= _178;
        119:
            _188 <= _179;
        120:
            _188 <= _180;
        121:
            _188 <= _181;
        122:
            _188 <= _182;
        123:
            _188 <= _183;
        124:
            _188 <= _184;
        125:
            _188 <= _185;
        126:
            _188 <= _186;
        default:
            _188 <= _187;
        endcase
    end
    assign _53 = _328 < _25;
    assign _189 = _53 ? _188 : _50;
    assign _190 = _40 ? _189 : _51;
    assign _336 = _48 ? _335 : _190;
    assign _3 = _336;
    always @(posedge _22) begin
        if (_20)
            _51 <= _50;
        else
            _51 <= _3;
    end
    assign _565 = 60'b000000000000000000000000000000000000000000000000000000000000;
    assign _566 = { _565,
                    _51 };
    assign _562 = 64'b0000000000000000000000000000000000000000000000000000000000001010;
    assign _563 = _561 * _562;
    assign _564 = _563[63:0];
    assign _567 = _564 + _566;
    assign _320 = _317 ? _314 : _311;
    assign _324 = _320 < _323;
    assign _325 = ~ _324;
    assign _191 = 4'b1010;
    assign _195 = _191 < _194;
    assign _318 = _198 ? _317 : _42;
    assign _319 = _318 & _195;
    assign _326 = _319 & _325;
    assign _345 = _326 ? _320 : _323;
    assign _340 = 8'b00001010;
    assign _341 = _57 + _340;
    always @* begin
        case (_341)
        0:
            _342 <= _60;
        1:
            _342 <= _61;
        2:
            _342 <= _62;
        3:
            _342 <= _63;
        4:
            _342 <= _64;
        5:
            _342 <= _65;
        6:
            _342 <= _66;
        7:
            _342 <= _67;
        8:
            _342 <= _68;
        9:
            _342 <= _69;
        10:
            _342 <= _70;
        11:
            _342 <= _71;
        12:
            _342 <= _72;
        13:
            _342 <= _73;
        14:
            _342 <= _74;
        15:
            _342 <= _75;
        16:
            _342 <= _76;
        17:
            _342 <= _77;
        18:
            _342 <= _78;
        19:
            _342 <= _79;
        20:
            _342 <= _80;
        21:
            _342 <= _81;
        22:
            _342 <= _82;
        23:
            _342 <= _83;
        24:
            _342 <= _84;
        25:
            _342 <= _85;
        26:
            _342 <= _86;
        27:
            _342 <= _87;
        28:
            _342 <= _88;
        29:
            _342 <= _89;
        30:
            _342 <= _90;
        31:
            _342 <= _91;
        32:
            _342 <= _92;
        33:
            _342 <= _93;
        34:
            _342 <= _94;
        35:
            _342 <= _95;
        36:
            _342 <= _96;
        37:
            _342 <= _97;
        38:
            _342 <= _98;
        39:
            _342 <= _99;
        40:
            _342 <= _100;
        41:
            _342 <= _101;
        42:
            _342 <= _102;
        43:
            _342 <= _103;
        44:
            _342 <= _104;
        45:
            _342 <= _105;
        46:
            _342 <= _106;
        47:
            _342 <= _107;
        48:
            _342 <= _108;
        49:
            _342 <= _109;
        50:
            _342 <= _110;
        51:
            _342 <= _111;
        52:
            _342 <= _112;
        53:
            _342 <= _113;
        54:
            _342 <= _114;
        55:
            _342 <= _115;
        56:
            _342 <= _116;
        57:
            _342 <= _117;
        58:
            _342 <= _118;
        59:
            _342 <= _119;
        60:
            _342 <= _120;
        61:
            _342 <= _121;
        62:
            _342 <= _122;
        63:
            _342 <= _123;
        64:
            _342 <= _124;
        65:
            _342 <= _125;
        66:
            _342 <= _126;
        67:
            _342 <= _127;
        68:
            _342 <= _128;
        69:
            _342 <= _129;
        70:
            _342 <= _130;
        71:
            _342 <= _131;
        72:
            _342 <= _132;
        73:
            _342 <= _133;
        74:
            _342 <= _134;
        75:
            _342 <= _135;
        76:
            _342 <= _136;
        77:
            _342 <= _137;
        78:
            _342 <= _138;
        79:
            _342 <= _139;
        80:
            _342 <= _140;
        81:
            _342 <= _141;
        82:
            _342 <= _142;
        83:
            _342 <= _143;
        84:
            _342 <= _144;
        85:
            _342 <= _145;
        86:
            _342 <= _146;
        87:
            _342 <= _147;
        88:
            _342 <= _148;
        89:
            _342 <= _149;
        90:
            _342 <= _150;
        91:
            _342 <= _151;
        92:
            _342 <= _152;
        93:
            _342 <= _153;
        94:
            _342 <= _154;
        95:
            _342 <= _155;
        96:
            _342 <= _156;
        97:
            _342 <= _157;
        98:
            _342 <= _158;
        99:
            _342 <= _159;
        100:
            _342 <= _160;
        101:
            _342 <= _161;
        102:
            _342 <= _162;
        103:
            _342 <= _163;
        104:
            _342 <= _164;
        105:
            _342 <= _165;
        106:
            _342 <= _166;
        107:
            _342 <= _167;
        108:
            _342 <= _168;
        109:
            _342 <= _169;
        110:
            _342 <= _170;
        111:
            _342 <= _171;
        112:
            _342 <= _172;
        113:
            _342 <= _173;
        114:
            _342 <= _174;
        115:
            _342 <= _175;
        116:
            _342 <= _176;
        117:
            _342 <= _177;
        118:
            _342 <= _178;
        119:
            _342 <= _179;
        120:
            _342 <= _180;
        121:
            _342 <= _181;
        122:
            _342 <= _182;
        123:
            _342 <= _183;
        124:
            _342 <= _184;
        125:
            _342 <= _185;
        126:
            _342 <= _186;
        default:
            _342 <= _187;
        endcase
    end
    assign _338 = _191 < _25;
    assign _343 = _338 ? _342 : _50;
    assign _344 = _40 ? _343 : _323;
    assign _346 = _48 ? _345 : _344;
    assign _4 = _346;
    always @(posedge _22) begin
        if (_20)
            _323 <= _50;
        else
            _323 <= _4;
    end
    assign _559 = { _565,
                    _323 };
    assign _556 = _554 * _562;
    assign _557 = _556[63:0];
    assign _560 = _557 + _559;
    assign _311 = _308 ? _305 : _302;
    assign _315 = _311 < _314;
    assign _316 = ~ _315;
    assign _197 = 4'b1001;
    assign _198 = _197 < _194;
    assign _309 = _201 ? _308 : _42;
    assign _310 = _309 & _198;
    assign _317 = _310 & _316;
    assign _355 = _317 ? _311 : _314;
    assign _350 = 8'b00001001;
    assign _351 = _57 + _350;
    always @* begin
        case (_351)
        0:
            _352 <= _60;
        1:
            _352 <= _61;
        2:
            _352 <= _62;
        3:
            _352 <= _63;
        4:
            _352 <= _64;
        5:
            _352 <= _65;
        6:
            _352 <= _66;
        7:
            _352 <= _67;
        8:
            _352 <= _68;
        9:
            _352 <= _69;
        10:
            _352 <= _70;
        11:
            _352 <= _71;
        12:
            _352 <= _72;
        13:
            _352 <= _73;
        14:
            _352 <= _74;
        15:
            _352 <= _75;
        16:
            _352 <= _76;
        17:
            _352 <= _77;
        18:
            _352 <= _78;
        19:
            _352 <= _79;
        20:
            _352 <= _80;
        21:
            _352 <= _81;
        22:
            _352 <= _82;
        23:
            _352 <= _83;
        24:
            _352 <= _84;
        25:
            _352 <= _85;
        26:
            _352 <= _86;
        27:
            _352 <= _87;
        28:
            _352 <= _88;
        29:
            _352 <= _89;
        30:
            _352 <= _90;
        31:
            _352 <= _91;
        32:
            _352 <= _92;
        33:
            _352 <= _93;
        34:
            _352 <= _94;
        35:
            _352 <= _95;
        36:
            _352 <= _96;
        37:
            _352 <= _97;
        38:
            _352 <= _98;
        39:
            _352 <= _99;
        40:
            _352 <= _100;
        41:
            _352 <= _101;
        42:
            _352 <= _102;
        43:
            _352 <= _103;
        44:
            _352 <= _104;
        45:
            _352 <= _105;
        46:
            _352 <= _106;
        47:
            _352 <= _107;
        48:
            _352 <= _108;
        49:
            _352 <= _109;
        50:
            _352 <= _110;
        51:
            _352 <= _111;
        52:
            _352 <= _112;
        53:
            _352 <= _113;
        54:
            _352 <= _114;
        55:
            _352 <= _115;
        56:
            _352 <= _116;
        57:
            _352 <= _117;
        58:
            _352 <= _118;
        59:
            _352 <= _119;
        60:
            _352 <= _120;
        61:
            _352 <= _121;
        62:
            _352 <= _122;
        63:
            _352 <= _123;
        64:
            _352 <= _124;
        65:
            _352 <= _125;
        66:
            _352 <= _126;
        67:
            _352 <= _127;
        68:
            _352 <= _128;
        69:
            _352 <= _129;
        70:
            _352 <= _130;
        71:
            _352 <= _131;
        72:
            _352 <= _132;
        73:
            _352 <= _133;
        74:
            _352 <= _134;
        75:
            _352 <= _135;
        76:
            _352 <= _136;
        77:
            _352 <= _137;
        78:
            _352 <= _138;
        79:
            _352 <= _139;
        80:
            _352 <= _140;
        81:
            _352 <= _141;
        82:
            _352 <= _142;
        83:
            _352 <= _143;
        84:
            _352 <= _144;
        85:
            _352 <= _145;
        86:
            _352 <= _146;
        87:
            _352 <= _147;
        88:
            _352 <= _148;
        89:
            _352 <= _149;
        90:
            _352 <= _150;
        91:
            _352 <= _151;
        92:
            _352 <= _152;
        93:
            _352 <= _153;
        94:
            _352 <= _154;
        95:
            _352 <= _155;
        96:
            _352 <= _156;
        97:
            _352 <= _157;
        98:
            _352 <= _158;
        99:
            _352 <= _159;
        100:
            _352 <= _160;
        101:
            _352 <= _161;
        102:
            _352 <= _162;
        103:
            _352 <= _163;
        104:
            _352 <= _164;
        105:
            _352 <= _165;
        106:
            _352 <= _166;
        107:
            _352 <= _167;
        108:
            _352 <= _168;
        109:
            _352 <= _169;
        110:
            _352 <= _170;
        111:
            _352 <= _171;
        112:
            _352 <= _172;
        113:
            _352 <= _173;
        114:
            _352 <= _174;
        115:
            _352 <= _175;
        116:
            _352 <= _176;
        117:
            _352 <= _177;
        118:
            _352 <= _178;
        119:
            _352 <= _179;
        120:
            _352 <= _180;
        121:
            _352 <= _181;
        122:
            _352 <= _182;
        123:
            _352 <= _183;
        124:
            _352 <= _184;
        125:
            _352 <= _185;
        126:
            _352 <= _186;
        default:
            _352 <= _187;
        endcase
    end
    assign _348 = _197 < _25;
    assign _353 = _348 ? _352 : _50;
    assign _354 = _40 ? _353 : _314;
    assign _356 = _48 ? _355 : _354;
    assign _5 = _356;
    always @(posedge _22) begin
        if (_20)
            _314 <= _50;
        else
            _314 <= _5;
    end
    assign _552 = { _565,
                    _314 };
    assign _549 = _547 * _562;
    assign _550 = _549[63:0];
    assign _553 = _550 + _552;
    assign _302 = _299 ? _296 : _293;
    assign _306 = _302 < _305;
    assign _307 = ~ _306;
    assign _200 = 4'b1000;
    assign _201 = _200 < _194;
    assign _300 = _204 ? _299 : _42;
    assign _301 = _300 & _201;
    assign _308 = _301 & _307;
    assign _365 = _308 ? _302 : _305;
    assign _360 = 8'b00001000;
    assign _361 = _57 + _360;
    always @* begin
        case (_361)
        0:
            _362 <= _60;
        1:
            _362 <= _61;
        2:
            _362 <= _62;
        3:
            _362 <= _63;
        4:
            _362 <= _64;
        5:
            _362 <= _65;
        6:
            _362 <= _66;
        7:
            _362 <= _67;
        8:
            _362 <= _68;
        9:
            _362 <= _69;
        10:
            _362 <= _70;
        11:
            _362 <= _71;
        12:
            _362 <= _72;
        13:
            _362 <= _73;
        14:
            _362 <= _74;
        15:
            _362 <= _75;
        16:
            _362 <= _76;
        17:
            _362 <= _77;
        18:
            _362 <= _78;
        19:
            _362 <= _79;
        20:
            _362 <= _80;
        21:
            _362 <= _81;
        22:
            _362 <= _82;
        23:
            _362 <= _83;
        24:
            _362 <= _84;
        25:
            _362 <= _85;
        26:
            _362 <= _86;
        27:
            _362 <= _87;
        28:
            _362 <= _88;
        29:
            _362 <= _89;
        30:
            _362 <= _90;
        31:
            _362 <= _91;
        32:
            _362 <= _92;
        33:
            _362 <= _93;
        34:
            _362 <= _94;
        35:
            _362 <= _95;
        36:
            _362 <= _96;
        37:
            _362 <= _97;
        38:
            _362 <= _98;
        39:
            _362 <= _99;
        40:
            _362 <= _100;
        41:
            _362 <= _101;
        42:
            _362 <= _102;
        43:
            _362 <= _103;
        44:
            _362 <= _104;
        45:
            _362 <= _105;
        46:
            _362 <= _106;
        47:
            _362 <= _107;
        48:
            _362 <= _108;
        49:
            _362 <= _109;
        50:
            _362 <= _110;
        51:
            _362 <= _111;
        52:
            _362 <= _112;
        53:
            _362 <= _113;
        54:
            _362 <= _114;
        55:
            _362 <= _115;
        56:
            _362 <= _116;
        57:
            _362 <= _117;
        58:
            _362 <= _118;
        59:
            _362 <= _119;
        60:
            _362 <= _120;
        61:
            _362 <= _121;
        62:
            _362 <= _122;
        63:
            _362 <= _123;
        64:
            _362 <= _124;
        65:
            _362 <= _125;
        66:
            _362 <= _126;
        67:
            _362 <= _127;
        68:
            _362 <= _128;
        69:
            _362 <= _129;
        70:
            _362 <= _130;
        71:
            _362 <= _131;
        72:
            _362 <= _132;
        73:
            _362 <= _133;
        74:
            _362 <= _134;
        75:
            _362 <= _135;
        76:
            _362 <= _136;
        77:
            _362 <= _137;
        78:
            _362 <= _138;
        79:
            _362 <= _139;
        80:
            _362 <= _140;
        81:
            _362 <= _141;
        82:
            _362 <= _142;
        83:
            _362 <= _143;
        84:
            _362 <= _144;
        85:
            _362 <= _145;
        86:
            _362 <= _146;
        87:
            _362 <= _147;
        88:
            _362 <= _148;
        89:
            _362 <= _149;
        90:
            _362 <= _150;
        91:
            _362 <= _151;
        92:
            _362 <= _152;
        93:
            _362 <= _153;
        94:
            _362 <= _154;
        95:
            _362 <= _155;
        96:
            _362 <= _156;
        97:
            _362 <= _157;
        98:
            _362 <= _158;
        99:
            _362 <= _159;
        100:
            _362 <= _160;
        101:
            _362 <= _161;
        102:
            _362 <= _162;
        103:
            _362 <= _163;
        104:
            _362 <= _164;
        105:
            _362 <= _165;
        106:
            _362 <= _166;
        107:
            _362 <= _167;
        108:
            _362 <= _168;
        109:
            _362 <= _169;
        110:
            _362 <= _170;
        111:
            _362 <= _171;
        112:
            _362 <= _172;
        113:
            _362 <= _173;
        114:
            _362 <= _174;
        115:
            _362 <= _175;
        116:
            _362 <= _176;
        117:
            _362 <= _177;
        118:
            _362 <= _178;
        119:
            _362 <= _179;
        120:
            _362 <= _180;
        121:
            _362 <= _181;
        122:
            _362 <= _182;
        123:
            _362 <= _183;
        124:
            _362 <= _184;
        125:
            _362 <= _185;
        126:
            _362 <= _186;
        default:
            _362 <= _187;
        endcase
    end
    assign _358 = _200 < _25;
    assign _363 = _358 ? _362 : _50;
    assign _364 = _40 ? _363 : _305;
    assign _366 = _48 ? _365 : _364;
    assign _6 = _366;
    always @(posedge _22) begin
        if (_20)
            _305 <= _50;
        else
            _305 <= _6;
    end
    assign _545 = { _565,
                    _305 };
    assign _542 = _540 * _562;
    assign _543 = _542[63:0];
    assign _546 = _543 + _545;
    assign _293 = _290 ? _287 : _284;
    assign _297 = _293 < _296;
    assign _298 = ~ _297;
    assign _203 = 4'b0111;
    assign _204 = _203 < _194;
    assign _291 = _207 ? _290 : _42;
    assign _292 = _291 & _204;
    assign _299 = _292 & _298;
    assign _375 = _299 ? _293 : _296;
    assign _370 = 8'b00000111;
    assign _371 = _57 + _370;
    always @* begin
        case (_371)
        0:
            _372 <= _60;
        1:
            _372 <= _61;
        2:
            _372 <= _62;
        3:
            _372 <= _63;
        4:
            _372 <= _64;
        5:
            _372 <= _65;
        6:
            _372 <= _66;
        7:
            _372 <= _67;
        8:
            _372 <= _68;
        9:
            _372 <= _69;
        10:
            _372 <= _70;
        11:
            _372 <= _71;
        12:
            _372 <= _72;
        13:
            _372 <= _73;
        14:
            _372 <= _74;
        15:
            _372 <= _75;
        16:
            _372 <= _76;
        17:
            _372 <= _77;
        18:
            _372 <= _78;
        19:
            _372 <= _79;
        20:
            _372 <= _80;
        21:
            _372 <= _81;
        22:
            _372 <= _82;
        23:
            _372 <= _83;
        24:
            _372 <= _84;
        25:
            _372 <= _85;
        26:
            _372 <= _86;
        27:
            _372 <= _87;
        28:
            _372 <= _88;
        29:
            _372 <= _89;
        30:
            _372 <= _90;
        31:
            _372 <= _91;
        32:
            _372 <= _92;
        33:
            _372 <= _93;
        34:
            _372 <= _94;
        35:
            _372 <= _95;
        36:
            _372 <= _96;
        37:
            _372 <= _97;
        38:
            _372 <= _98;
        39:
            _372 <= _99;
        40:
            _372 <= _100;
        41:
            _372 <= _101;
        42:
            _372 <= _102;
        43:
            _372 <= _103;
        44:
            _372 <= _104;
        45:
            _372 <= _105;
        46:
            _372 <= _106;
        47:
            _372 <= _107;
        48:
            _372 <= _108;
        49:
            _372 <= _109;
        50:
            _372 <= _110;
        51:
            _372 <= _111;
        52:
            _372 <= _112;
        53:
            _372 <= _113;
        54:
            _372 <= _114;
        55:
            _372 <= _115;
        56:
            _372 <= _116;
        57:
            _372 <= _117;
        58:
            _372 <= _118;
        59:
            _372 <= _119;
        60:
            _372 <= _120;
        61:
            _372 <= _121;
        62:
            _372 <= _122;
        63:
            _372 <= _123;
        64:
            _372 <= _124;
        65:
            _372 <= _125;
        66:
            _372 <= _126;
        67:
            _372 <= _127;
        68:
            _372 <= _128;
        69:
            _372 <= _129;
        70:
            _372 <= _130;
        71:
            _372 <= _131;
        72:
            _372 <= _132;
        73:
            _372 <= _133;
        74:
            _372 <= _134;
        75:
            _372 <= _135;
        76:
            _372 <= _136;
        77:
            _372 <= _137;
        78:
            _372 <= _138;
        79:
            _372 <= _139;
        80:
            _372 <= _140;
        81:
            _372 <= _141;
        82:
            _372 <= _142;
        83:
            _372 <= _143;
        84:
            _372 <= _144;
        85:
            _372 <= _145;
        86:
            _372 <= _146;
        87:
            _372 <= _147;
        88:
            _372 <= _148;
        89:
            _372 <= _149;
        90:
            _372 <= _150;
        91:
            _372 <= _151;
        92:
            _372 <= _152;
        93:
            _372 <= _153;
        94:
            _372 <= _154;
        95:
            _372 <= _155;
        96:
            _372 <= _156;
        97:
            _372 <= _157;
        98:
            _372 <= _158;
        99:
            _372 <= _159;
        100:
            _372 <= _160;
        101:
            _372 <= _161;
        102:
            _372 <= _162;
        103:
            _372 <= _163;
        104:
            _372 <= _164;
        105:
            _372 <= _165;
        106:
            _372 <= _166;
        107:
            _372 <= _167;
        108:
            _372 <= _168;
        109:
            _372 <= _169;
        110:
            _372 <= _170;
        111:
            _372 <= _171;
        112:
            _372 <= _172;
        113:
            _372 <= _173;
        114:
            _372 <= _174;
        115:
            _372 <= _175;
        116:
            _372 <= _176;
        117:
            _372 <= _177;
        118:
            _372 <= _178;
        119:
            _372 <= _179;
        120:
            _372 <= _180;
        121:
            _372 <= _181;
        122:
            _372 <= _182;
        123:
            _372 <= _183;
        124:
            _372 <= _184;
        125:
            _372 <= _185;
        126:
            _372 <= _186;
        default:
            _372 <= _187;
        endcase
    end
    assign _368 = _203 < _25;
    assign _373 = _368 ? _372 : _50;
    assign _374 = _40 ? _373 : _296;
    assign _376 = _48 ? _375 : _374;
    assign _7 = _376;
    always @(posedge _22) begin
        if (_20)
            _296 <= _50;
        else
            _296 <= _7;
    end
    assign _538 = { _565,
                    _296 };
    assign _535 = _533 * _562;
    assign _536 = _535[63:0];
    assign _539 = _536 + _538;
    assign _284 = _281 ? _278 : _275;
    assign _288 = _284 < _287;
    assign _289 = ~ _288;
    assign _206 = 4'b0110;
    assign _207 = _206 < _194;
    assign _282 = _210 ? _281 : _42;
    assign _283 = _282 & _207;
    assign _290 = _283 & _289;
    assign _385 = _290 ? _284 : _287;
    assign _380 = 8'b00000110;
    assign _381 = _57 + _380;
    always @* begin
        case (_381)
        0:
            _382 <= _60;
        1:
            _382 <= _61;
        2:
            _382 <= _62;
        3:
            _382 <= _63;
        4:
            _382 <= _64;
        5:
            _382 <= _65;
        6:
            _382 <= _66;
        7:
            _382 <= _67;
        8:
            _382 <= _68;
        9:
            _382 <= _69;
        10:
            _382 <= _70;
        11:
            _382 <= _71;
        12:
            _382 <= _72;
        13:
            _382 <= _73;
        14:
            _382 <= _74;
        15:
            _382 <= _75;
        16:
            _382 <= _76;
        17:
            _382 <= _77;
        18:
            _382 <= _78;
        19:
            _382 <= _79;
        20:
            _382 <= _80;
        21:
            _382 <= _81;
        22:
            _382 <= _82;
        23:
            _382 <= _83;
        24:
            _382 <= _84;
        25:
            _382 <= _85;
        26:
            _382 <= _86;
        27:
            _382 <= _87;
        28:
            _382 <= _88;
        29:
            _382 <= _89;
        30:
            _382 <= _90;
        31:
            _382 <= _91;
        32:
            _382 <= _92;
        33:
            _382 <= _93;
        34:
            _382 <= _94;
        35:
            _382 <= _95;
        36:
            _382 <= _96;
        37:
            _382 <= _97;
        38:
            _382 <= _98;
        39:
            _382 <= _99;
        40:
            _382 <= _100;
        41:
            _382 <= _101;
        42:
            _382 <= _102;
        43:
            _382 <= _103;
        44:
            _382 <= _104;
        45:
            _382 <= _105;
        46:
            _382 <= _106;
        47:
            _382 <= _107;
        48:
            _382 <= _108;
        49:
            _382 <= _109;
        50:
            _382 <= _110;
        51:
            _382 <= _111;
        52:
            _382 <= _112;
        53:
            _382 <= _113;
        54:
            _382 <= _114;
        55:
            _382 <= _115;
        56:
            _382 <= _116;
        57:
            _382 <= _117;
        58:
            _382 <= _118;
        59:
            _382 <= _119;
        60:
            _382 <= _120;
        61:
            _382 <= _121;
        62:
            _382 <= _122;
        63:
            _382 <= _123;
        64:
            _382 <= _124;
        65:
            _382 <= _125;
        66:
            _382 <= _126;
        67:
            _382 <= _127;
        68:
            _382 <= _128;
        69:
            _382 <= _129;
        70:
            _382 <= _130;
        71:
            _382 <= _131;
        72:
            _382 <= _132;
        73:
            _382 <= _133;
        74:
            _382 <= _134;
        75:
            _382 <= _135;
        76:
            _382 <= _136;
        77:
            _382 <= _137;
        78:
            _382 <= _138;
        79:
            _382 <= _139;
        80:
            _382 <= _140;
        81:
            _382 <= _141;
        82:
            _382 <= _142;
        83:
            _382 <= _143;
        84:
            _382 <= _144;
        85:
            _382 <= _145;
        86:
            _382 <= _146;
        87:
            _382 <= _147;
        88:
            _382 <= _148;
        89:
            _382 <= _149;
        90:
            _382 <= _150;
        91:
            _382 <= _151;
        92:
            _382 <= _152;
        93:
            _382 <= _153;
        94:
            _382 <= _154;
        95:
            _382 <= _155;
        96:
            _382 <= _156;
        97:
            _382 <= _157;
        98:
            _382 <= _158;
        99:
            _382 <= _159;
        100:
            _382 <= _160;
        101:
            _382 <= _161;
        102:
            _382 <= _162;
        103:
            _382 <= _163;
        104:
            _382 <= _164;
        105:
            _382 <= _165;
        106:
            _382 <= _166;
        107:
            _382 <= _167;
        108:
            _382 <= _168;
        109:
            _382 <= _169;
        110:
            _382 <= _170;
        111:
            _382 <= _171;
        112:
            _382 <= _172;
        113:
            _382 <= _173;
        114:
            _382 <= _174;
        115:
            _382 <= _175;
        116:
            _382 <= _176;
        117:
            _382 <= _177;
        118:
            _382 <= _178;
        119:
            _382 <= _179;
        120:
            _382 <= _180;
        121:
            _382 <= _181;
        122:
            _382 <= _182;
        123:
            _382 <= _183;
        124:
            _382 <= _184;
        125:
            _382 <= _185;
        126:
            _382 <= _186;
        default:
            _382 <= _187;
        endcase
    end
    assign _378 = _206 < _25;
    assign _383 = _378 ? _382 : _50;
    assign _384 = _40 ? _383 : _287;
    assign _386 = _48 ? _385 : _384;
    assign _8 = _386;
    always @(posedge _22) begin
        if (_20)
            _287 <= _50;
        else
            _287 <= _8;
    end
    assign _531 = { _565,
                    _287 };
    assign _528 = _526 * _562;
    assign _529 = _528[63:0];
    assign _532 = _529 + _531;
    assign _275 = _272 ? _269 : _266;
    assign _279 = _275 < _278;
    assign _280 = ~ _279;
    assign _209 = 4'b0101;
    assign _210 = _209 < _194;
    assign _273 = _213 ? _272 : _42;
    assign _274 = _273 & _210;
    assign _281 = _274 & _280;
    assign _395 = _281 ? _275 : _278;
    assign _390 = 8'b00000101;
    assign _391 = _57 + _390;
    always @* begin
        case (_391)
        0:
            _392 <= _60;
        1:
            _392 <= _61;
        2:
            _392 <= _62;
        3:
            _392 <= _63;
        4:
            _392 <= _64;
        5:
            _392 <= _65;
        6:
            _392 <= _66;
        7:
            _392 <= _67;
        8:
            _392 <= _68;
        9:
            _392 <= _69;
        10:
            _392 <= _70;
        11:
            _392 <= _71;
        12:
            _392 <= _72;
        13:
            _392 <= _73;
        14:
            _392 <= _74;
        15:
            _392 <= _75;
        16:
            _392 <= _76;
        17:
            _392 <= _77;
        18:
            _392 <= _78;
        19:
            _392 <= _79;
        20:
            _392 <= _80;
        21:
            _392 <= _81;
        22:
            _392 <= _82;
        23:
            _392 <= _83;
        24:
            _392 <= _84;
        25:
            _392 <= _85;
        26:
            _392 <= _86;
        27:
            _392 <= _87;
        28:
            _392 <= _88;
        29:
            _392 <= _89;
        30:
            _392 <= _90;
        31:
            _392 <= _91;
        32:
            _392 <= _92;
        33:
            _392 <= _93;
        34:
            _392 <= _94;
        35:
            _392 <= _95;
        36:
            _392 <= _96;
        37:
            _392 <= _97;
        38:
            _392 <= _98;
        39:
            _392 <= _99;
        40:
            _392 <= _100;
        41:
            _392 <= _101;
        42:
            _392 <= _102;
        43:
            _392 <= _103;
        44:
            _392 <= _104;
        45:
            _392 <= _105;
        46:
            _392 <= _106;
        47:
            _392 <= _107;
        48:
            _392 <= _108;
        49:
            _392 <= _109;
        50:
            _392 <= _110;
        51:
            _392 <= _111;
        52:
            _392 <= _112;
        53:
            _392 <= _113;
        54:
            _392 <= _114;
        55:
            _392 <= _115;
        56:
            _392 <= _116;
        57:
            _392 <= _117;
        58:
            _392 <= _118;
        59:
            _392 <= _119;
        60:
            _392 <= _120;
        61:
            _392 <= _121;
        62:
            _392 <= _122;
        63:
            _392 <= _123;
        64:
            _392 <= _124;
        65:
            _392 <= _125;
        66:
            _392 <= _126;
        67:
            _392 <= _127;
        68:
            _392 <= _128;
        69:
            _392 <= _129;
        70:
            _392 <= _130;
        71:
            _392 <= _131;
        72:
            _392 <= _132;
        73:
            _392 <= _133;
        74:
            _392 <= _134;
        75:
            _392 <= _135;
        76:
            _392 <= _136;
        77:
            _392 <= _137;
        78:
            _392 <= _138;
        79:
            _392 <= _139;
        80:
            _392 <= _140;
        81:
            _392 <= _141;
        82:
            _392 <= _142;
        83:
            _392 <= _143;
        84:
            _392 <= _144;
        85:
            _392 <= _145;
        86:
            _392 <= _146;
        87:
            _392 <= _147;
        88:
            _392 <= _148;
        89:
            _392 <= _149;
        90:
            _392 <= _150;
        91:
            _392 <= _151;
        92:
            _392 <= _152;
        93:
            _392 <= _153;
        94:
            _392 <= _154;
        95:
            _392 <= _155;
        96:
            _392 <= _156;
        97:
            _392 <= _157;
        98:
            _392 <= _158;
        99:
            _392 <= _159;
        100:
            _392 <= _160;
        101:
            _392 <= _161;
        102:
            _392 <= _162;
        103:
            _392 <= _163;
        104:
            _392 <= _164;
        105:
            _392 <= _165;
        106:
            _392 <= _166;
        107:
            _392 <= _167;
        108:
            _392 <= _168;
        109:
            _392 <= _169;
        110:
            _392 <= _170;
        111:
            _392 <= _171;
        112:
            _392 <= _172;
        113:
            _392 <= _173;
        114:
            _392 <= _174;
        115:
            _392 <= _175;
        116:
            _392 <= _176;
        117:
            _392 <= _177;
        118:
            _392 <= _178;
        119:
            _392 <= _179;
        120:
            _392 <= _180;
        121:
            _392 <= _181;
        122:
            _392 <= _182;
        123:
            _392 <= _183;
        124:
            _392 <= _184;
        125:
            _392 <= _185;
        126:
            _392 <= _186;
        default:
            _392 <= _187;
        endcase
    end
    assign _388 = _209 < _25;
    assign _393 = _388 ? _392 : _50;
    assign _394 = _40 ? _393 : _278;
    assign _396 = _48 ? _395 : _394;
    assign _9 = _396;
    always @(posedge _22) begin
        if (_20)
            _278 <= _50;
        else
            _278 <= _9;
    end
    assign _524 = { _565,
                    _278 };
    assign _521 = _519 * _562;
    assign _522 = _521[63:0];
    assign _525 = _522 + _524;
    assign _266 = _263 ? _260 : _257;
    assign _270 = _266 < _269;
    assign _271 = ~ _270;
    assign _212 = 4'b0100;
    assign _213 = _212 < _194;
    assign _264 = _216 ? _263 : _42;
    assign _265 = _264 & _213;
    assign _272 = _265 & _271;
    assign _405 = _272 ? _266 : _269;
    assign _400 = 8'b00000100;
    assign _401 = _57 + _400;
    always @* begin
        case (_401)
        0:
            _402 <= _60;
        1:
            _402 <= _61;
        2:
            _402 <= _62;
        3:
            _402 <= _63;
        4:
            _402 <= _64;
        5:
            _402 <= _65;
        6:
            _402 <= _66;
        7:
            _402 <= _67;
        8:
            _402 <= _68;
        9:
            _402 <= _69;
        10:
            _402 <= _70;
        11:
            _402 <= _71;
        12:
            _402 <= _72;
        13:
            _402 <= _73;
        14:
            _402 <= _74;
        15:
            _402 <= _75;
        16:
            _402 <= _76;
        17:
            _402 <= _77;
        18:
            _402 <= _78;
        19:
            _402 <= _79;
        20:
            _402 <= _80;
        21:
            _402 <= _81;
        22:
            _402 <= _82;
        23:
            _402 <= _83;
        24:
            _402 <= _84;
        25:
            _402 <= _85;
        26:
            _402 <= _86;
        27:
            _402 <= _87;
        28:
            _402 <= _88;
        29:
            _402 <= _89;
        30:
            _402 <= _90;
        31:
            _402 <= _91;
        32:
            _402 <= _92;
        33:
            _402 <= _93;
        34:
            _402 <= _94;
        35:
            _402 <= _95;
        36:
            _402 <= _96;
        37:
            _402 <= _97;
        38:
            _402 <= _98;
        39:
            _402 <= _99;
        40:
            _402 <= _100;
        41:
            _402 <= _101;
        42:
            _402 <= _102;
        43:
            _402 <= _103;
        44:
            _402 <= _104;
        45:
            _402 <= _105;
        46:
            _402 <= _106;
        47:
            _402 <= _107;
        48:
            _402 <= _108;
        49:
            _402 <= _109;
        50:
            _402 <= _110;
        51:
            _402 <= _111;
        52:
            _402 <= _112;
        53:
            _402 <= _113;
        54:
            _402 <= _114;
        55:
            _402 <= _115;
        56:
            _402 <= _116;
        57:
            _402 <= _117;
        58:
            _402 <= _118;
        59:
            _402 <= _119;
        60:
            _402 <= _120;
        61:
            _402 <= _121;
        62:
            _402 <= _122;
        63:
            _402 <= _123;
        64:
            _402 <= _124;
        65:
            _402 <= _125;
        66:
            _402 <= _126;
        67:
            _402 <= _127;
        68:
            _402 <= _128;
        69:
            _402 <= _129;
        70:
            _402 <= _130;
        71:
            _402 <= _131;
        72:
            _402 <= _132;
        73:
            _402 <= _133;
        74:
            _402 <= _134;
        75:
            _402 <= _135;
        76:
            _402 <= _136;
        77:
            _402 <= _137;
        78:
            _402 <= _138;
        79:
            _402 <= _139;
        80:
            _402 <= _140;
        81:
            _402 <= _141;
        82:
            _402 <= _142;
        83:
            _402 <= _143;
        84:
            _402 <= _144;
        85:
            _402 <= _145;
        86:
            _402 <= _146;
        87:
            _402 <= _147;
        88:
            _402 <= _148;
        89:
            _402 <= _149;
        90:
            _402 <= _150;
        91:
            _402 <= _151;
        92:
            _402 <= _152;
        93:
            _402 <= _153;
        94:
            _402 <= _154;
        95:
            _402 <= _155;
        96:
            _402 <= _156;
        97:
            _402 <= _157;
        98:
            _402 <= _158;
        99:
            _402 <= _159;
        100:
            _402 <= _160;
        101:
            _402 <= _161;
        102:
            _402 <= _162;
        103:
            _402 <= _163;
        104:
            _402 <= _164;
        105:
            _402 <= _165;
        106:
            _402 <= _166;
        107:
            _402 <= _167;
        108:
            _402 <= _168;
        109:
            _402 <= _169;
        110:
            _402 <= _170;
        111:
            _402 <= _171;
        112:
            _402 <= _172;
        113:
            _402 <= _173;
        114:
            _402 <= _174;
        115:
            _402 <= _175;
        116:
            _402 <= _176;
        117:
            _402 <= _177;
        118:
            _402 <= _178;
        119:
            _402 <= _179;
        120:
            _402 <= _180;
        121:
            _402 <= _181;
        122:
            _402 <= _182;
        123:
            _402 <= _183;
        124:
            _402 <= _184;
        125:
            _402 <= _185;
        126:
            _402 <= _186;
        default:
            _402 <= _187;
        endcase
    end
    assign _398 = _212 < _25;
    assign _403 = _398 ? _402 : _50;
    assign _404 = _40 ? _403 : _269;
    assign _406 = _48 ? _405 : _404;
    assign _10 = _406;
    always @(posedge _22) begin
        if (_20)
            _269 <= _50;
        else
            _269 <= _10;
    end
    assign _517 = { _565,
                    _269 };
    assign _514 = _512 * _562;
    assign _515 = _514[63:0];
    assign _518 = _515 + _517;
    assign _257 = _254 ? _251 : _248;
    assign _261 = _257 < _260;
    assign _262 = ~ _261;
    assign _215 = 4'b0011;
    assign _216 = _215 < _194;
    assign _255 = _219 ? _254 : _42;
    assign _256 = _255 & _216;
    assign _263 = _256 & _262;
    assign _415 = _263 ? _257 : _260;
    assign _410 = 8'b00000011;
    assign _411 = _57 + _410;
    always @* begin
        case (_411)
        0:
            _412 <= _60;
        1:
            _412 <= _61;
        2:
            _412 <= _62;
        3:
            _412 <= _63;
        4:
            _412 <= _64;
        5:
            _412 <= _65;
        6:
            _412 <= _66;
        7:
            _412 <= _67;
        8:
            _412 <= _68;
        9:
            _412 <= _69;
        10:
            _412 <= _70;
        11:
            _412 <= _71;
        12:
            _412 <= _72;
        13:
            _412 <= _73;
        14:
            _412 <= _74;
        15:
            _412 <= _75;
        16:
            _412 <= _76;
        17:
            _412 <= _77;
        18:
            _412 <= _78;
        19:
            _412 <= _79;
        20:
            _412 <= _80;
        21:
            _412 <= _81;
        22:
            _412 <= _82;
        23:
            _412 <= _83;
        24:
            _412 <= _84;
        25:
            _412 <= _85;
        26:
            _412 <= _86;
        27:
            _412 <= _87;
        28:
            _412 <= _88;
        29:
            _412 <= _89;
        30:
            _412 <= _90;
        31:
            _412 <= _91;
        32:
            _412 <= _92;
        33:
            _412 <= _93;
        34:
            _412 <= _94;
        35:
            _412 <= _95;
        36:
            _412 <= _96;
        37:
            _412 <= _97;
        38:
            _412 <= _98;
        39:
            _412 <= _99;
        40:
            _412 <= _100;
        41:
            _412 <= _101;
        42:
            _412 <= _102;
        43:
            _412 <= _103;
        44:
            _412 <= _104;
        45:
            _412 <= _105;
        46:
            _412 <= _106;
        47:
            _412 <= _107;
        48:
            _412 <= _108;
        49:
            _412 <= _109;
        50:
            _412 <= _110;
        51:
            _412 <= _111;
        52:
            _412 <= _112;
        53:
            _412 <= _113;
        54:
            _412 <= _114;
        55:
            _412 <= _115;
        56:
            _412 <= _116;
        57:
            _412 <= _117;
        58:
            _412 <= _118;
        59:
            _412 <= _119;
        60:
            _412 <= _120;
        61:
            _412 <= _121;
        62:
            _412 <= _122;
        63:
            _412 <= _123;
        64:
            _412 <= _124;
        65:
            _412 <= _125;
        66:
            _412 <= _126;
        67:
            _412 <= _127;
        68:
            _412 <= _128;
        69:
            _412 <= _129;
        70:
            _412 <= _130;
        71:
            _412 <= _131;
        72:
            _412 <= _132;
        73:
            _412 <= _133;
        74:
            _412 <= _134;
        75:
            _412 <= _135;
        76:
            _412 <= _136;
        77:
            _412 <= _137;
        78:
            _412 <= _138;
        79:
            _412 <= _139;
        80:
            _412 <= _140;
        81:
            _412 <= _141;
        82:
            _412 <= _142;
        83:
            _412 <= _143;
        84:
            _412 <= _144;
        85:
            _412 <= _145;
        86:
            _412 <= _146;
        87:
            _412 <= _147;
        88:
            _412 <= _148;
        89:
            _412 <= _149;
        90:
            _412 <= _150;
        91:
            _412 <= _151;
        92:
            _412 <= _152;
        93:
            _412 <= _153;
        94:
            _412 <= _154;
        95:
            _412 <= _155;
        96:
            _412 <= _156;
        97:
            _412 <= _157;
        98:
            _412 <= _158;
        99:
            _412 <= _159;
        100:
            _412 <= _160;
        101:
            _412 <= _161;
        102:
            _412 <= _162;
        103:
            _412 <= _163;
        104:
            _412 <= _164;
        105:
            _412 <= _165;
        106:
            _412 <= _166;
        107:
            _412 <= _167;
        108:
            _412 <= _168;
        109:
            _412 <= _169;
        110:
            _412 <= _170;
        111:
            _412 <= _171;
        112:
            _412 <= _172;
        113:
            _412 <= _173;
        114:
            _412 <= _174;
        115:
            _412 <= _175;
        116:
            _412 <= _176;
        117:
            _412 <= _177;
        118:
            _412 <= _178;
        119:
            _412 <= _179;
        120:
            _412 <= _180;
        121:
            _412 <= _181;
        122:
            _412 <= _182;
        123:
            _412 <= _183;
        124:
            _412 <= _184;
        125:
            _412 <= _185;
        126:
            _412 <= _186;
        default:
            _412 <= _187;
        endcase
    end
    assign _408 = _215 < _25;
    assign _413 = _408 ? _412 : _50;
    assign _414 = _40 ? _413 : _260;
    assign _416 = _48 ? _415 : _414;
    assign _11 = _416;
    always @(posedge _22) begin
        if (_20)
            _260 <= _50;
        else
            _260 <= _11;
    end
    assign _510 = { _565,
                    _260 };
    assign _507 = _505 * _562;
    assign _508 = _507[63:0];
    assign _511 = _508 + _510;
    assign _248 = _245 ? _242 : _239;
    assign _252 = _248 < _251;
    assign _253 = ~ _252;
    assign _218 = 4'b0010;
    assign _219 = _218 < _194;
    assign _246 = _222 ? _245 : _42;
    assign _247 = _246 & _219;
    assign _254 = _247 & _253;
    assign _425 = _254 ? _248 : _251;
    assign _420 = 8'b00000010;
    assign _421 = _57 + _420;
    always @* begin
        case (_421)
        0:
            _422 <= _60;
        1:
            _422 <= _61;
        2:
            _422 <= _62;
        3:
            _422 <= _63;
        4:
            _422 <= _64;
        5:
            _422 <= _65;
        6:
            _422 <= _66;
        7:
            _422 <= _67;
        8:
            _422 <= _68;
        9:
            _422 <= _69;
        10:
            _422 <= _70;
        11:
            _422 <= _71;
        12:
            _422 <= _72;
        13:
            _422 <= _73;
        14:
            _422 <= _74;
        15:
            _422 <= _75;
        16:
            _422 <= _76;
        17:
            _422 <= _77;
        18:
            _422 <= _78;
        19:
            _422 <= _79;
        20:
            _422 <= _80;
        21:
            _422 <= _81;
        22:
            _422 <= _82;
        23:
            _422 <= _83;
        24:
            _422 <= _84;
        25:
            _422 <= _85;
        26:
            _422 <= _86;
        27:
            _422 <= _87;
        28:
            _422 <= _88;
        29:
            _422 <= _89;
        30:
            _422 <= _90;
        31:
            _422 <= _91;
        32:
            _422 <= _92;
        33:
            _422 <= _93;
        34:
            _422 <= _94;
        35:
            _422 <= _95;
        36:
            _422 <= _96;
        37:
            _422 <= _97;
        38:
            _422 <= _98;
        39:
            _422 <= _99;
        40:
            _422 <= _100;
        41:
            _422 <= _101;
        42:
            _422 <= _102;
        43:
            _422 <= _103;
        44:
            _422 <= _104;
        45:
            _422 <= _105;
        46:
            _422 <= _106;
        47:
            _422 <= _107;
        48:
            _422 <= _108;
        49:
            _422 <= _109;
        50:
            _422 <= _110;
        51:
            _422 <= _111;
        52:
            _422 <= _112;
        53:
            _422 <= _113;
        54:
            _422 <= _114;
        55:
            _422 <= _115;
        56:
            _422 <= _116;
        57:
            _422 <= _117;
        58:
            _422 <= _118;
        59:
            _422 <= _119;
        60:
            _422 <= _120;
        61:
            _422 <= _121;
        62:
            _422 <= _122;
        63:
            _422 <= _123;
        64:
            _422 <= _124;
        65:
            _422 <= _125;
        66:
            _422 <= _126;
        67:
            _422 <= _127;
        68:
            _422 <= _128;
        69:
            _422 <= _129;
        70:
            _422 <= _130;
        71:
            _422 <= _131;
        72:
            _422 <= _132;
        73:
            _422 <= _133;
        74:
            _422 <= _134;
        75:
            _422 <= _135;
        76:
            _422 <= _136;
        77:
            _422 <= _137;
        78:
            _422 <= _138;
        79:
            _422 <= _139;
        80:
            _422 <= _140;
        81:
            _422 <= _141;
        82:
            _422 <= _142;
        83:
            _422 <= _143;
        84:
            _422 <= _144;
        85:
            _422 <= _145;
        86:
            _422 <= _146;
        87:
            _422 <= _147;
        88:
            _422 <= _148;
        89:
            _422 <= _149;
        90:
            _422 <= _150;
        91:
            _422 <= _151;
        92:
            _422 <= _152;
        93:
            _422 <= _153;
        94:
            _422 <= _154;
        95:
            _422 <= _155;
        96:
            _422 <= _156;
        97:
            _422 <= _157;
        98:
            _422 <= _158;
        99:
            _422 <= _159;
        100:
            _422 <= _160;
        101:
            _422 <= _161;
        102:
            _422 <= _162;
        103:
            _422 <= _163;
        104:
            _422 <= _164;
        105:
            _422 <= _165;
        106:
            _422 <= _166;
        107:
            _422 <= _167;
        108:
            _422 <= _168;
        109:
            _422 <= _169;
        110:
            _422 <= _170;
        111:
            _422 <= _171;
        112:
            _422 <= _172;
        113:
            _422 <= _173;
        114:
            _422 <= _174;
        115:
            _422 <= _175;
        116:
            _422 <= _176;
        117:
            _422 <= _177;
        118:
            _422 <= _178;
        119:
            _422 <= _179;
        120:
            _422 <= _180;
        121:
            _422 <= _181;
        122:
            _422 <= _182;
        123:
            _422 <= _183;
        124:
            _422 <= _184;
        125:
            _422 <= _185;
        126:
            _422 <= _186;
        default:
            _422 <= _187;
        endcase
    end
    assign _418 = _218 < _25;
    assign _423 = _418 ? _422 : _50;
    assign _424 = _40 ? _423 : _251;
    assign _426 = _48 ? _425 : _424;
    assign _12 = _426;
    always @(posedge _22) begin
        if (_20)
            _251 <= _50;
        else
            _251 <= _12;
    end
    assign _503 = { _565,
                    _251 };
    assign _500 = _498 * _562;
    assign _501 = _500[63:0];
    assign _504 = _501 + _503;
    assign _239 = _236 ? _233 : _230;
    assign _243 = _239 < _242;
    assign _244 = ~ _243;
    assign _221 = 4'b0001;
    assign _222 = _221 < _194;
    assign _237 = _225 ? _236 : _42;
    assign _238 = _237 & _222;
    assign _245 = _238 & _244;
    assign _435 = _245 ? _239 : _242;
    assign _430 = 8'b00000001;
    assign _431 = _57 + _430;
    always @* begin
        case (_431)
        0:
            _432 <= _60;
        1:
            _432 <= _61;
        2:
            _432 <= _62;
        3:
            _432 <= _63;
        4:
            _432 <= _64;
        5:
            _432 <= _65;
        6:
            _432 <= _66;
        7:
            _432 <= _67;
        8:
            _432 <= _68;
        9:
            _432 <= _69;
        10:
            _432 <= _70;
        11:
            _432 <= _71;
        12:
            _432 <= _72;
        13:
            _432 <= _73;
        14:
            _432 <= _74;
        15:
            _432 <= _75;
        16:
            _432 <= _76;
        17:
            _432 <= _77;
        18:
            _432 <= _78;
        19:
            _432 <= _79;
        20:
            _432 <= _80;
        21:
            _432 <= _81;
        22:
            _432 <= _82;
        23:
            _432 <= _83;
        24:
            _432 <= _84;
        25:
            _432 <= _85;
        26:
            _432 <= _86;
        27:
            _432 <= _87;
        28:
            _432 <= _88;
        29:
            _432 <= _89;
        30:
            _432 <= _90;
        31:
            _432 <= _91;
        32:
            _432 <= _92;
        33:
            _432 <= _93;
        34:
            _432 <= _94;
        35:
            _432 <= _95;
        36:
            _432 <= _96;
        37:
            _432 <= _97;
        38:
            _432 <= _98;
        39:
            _432 <= _99;
        40:
            _432 <= _100;
        41:
            _432 <= _101;
        42:
            _432 <= _102;
        43:
            _432 <= _103;
        44:
            _432 <= _104;
        45:
            _432 <= _105;
        46:
            _432 <= _106;
        47:
            _432 <= _107;
        48:
            _432 <= _108;
        49:
            _432 <= _109;
        50:
            _432 <= _110;
        51:
            _432 <= _111;
        52:
            _432 <= _112;
        53:
            _432 <= _113;
        54:
            _432 <= _114;
        55:
            _432 <= _115;
        56:
            _432 <= _116;
        57:
            _432 <= _117;
        58:
            _432 <= _118;
        59:
            _432 <= _119;
        60:
            _432 <= _120;
        61:
            _432 <= _121;
        62:
            _432 <= _122;
        63:
            _432 <= _123;
        64:
            _432 <= _124;
        65:
            _432 <= _125;
        66:
            _432 <= _126;
        67:
            _432 <= _127;
        68:
            _432 <= _128;
        69:
            _432 <= _129;
        70:
            _432 <= _130;
        71:
            _432 <= _131;
        72:
            _432 <= _132;
        73:
            _432 <= _133;
        74:
            _432 <= _134;
        75:
            _432 <= _135;
        76:
            _432 <= _136;
        77:
            _432 <= _137;
        78:
            _432 <= _138;
        79:
            _432 <= _139;
        80:
            _432 <= _140;
        81:
            _432 <= _141;
        82:
            _432 <= _142;
        83:
            _432 <= _143;
        84:
            _432 <= _144;
        85:
            _432 <= _145;
        86:
            _432 <= _146;
        87:
            _432 <= _147;
        88:
            _432 <= _148;
        89:
            _432 <= _149;
        90:
            _432 <= _150;
        91:
            _432 <= _151;
        92:
            _432 <= _152;
        93:
            _432 <= _153;
        94:
            _432 <= _154;
        95:
            _432 <= _155;
        96:
            _432 <= _156;
        97:
            _432 <= _157;
        98:
            _432 <= _158;
        99:
            _432 <= _159;
        100:
            _432 <= _160;
        101:
            _432 <= _161;
        102:
            _432 <= _162;
        103:
            _432 <= _163;
        104:
            _432 <= _164;
        105:
            _432 <= _165;
        106:
            _432 <= _166;
        107:
            _432 <= _167;
        108:
            _432 <= _168;
        109:
            _432 <= _169;
        110:
            _432 <= _170;
        111:
            _432 <= _171;
        112:
            _432 <= _172;
        113:
            _432 <= _173;
        114:
            _432 <= _174;
        115:
            _432 <= _175;
        116:
            _432 <= _176;
        117:
            _432 <= _177;
        118:
            _432 <= _178;
        119:
            _432 <= _179;
        120:
            _432 <= _180;
        121:
            _432 <= _181;
        122:
            _432 <= _182;
        123:
            _432 <= _183;
        124:
            _432 <= _184;
        125:
            _432 <= _185;
        126:
            _432 <= _186;
        default:
            _432 <= _187;
        endcase
    end
    assign _428 = _221 < _25;
    assign _433 = _428 ? _432 : _50;
    assign _434 = _40 ? _433 : _242;
    assign _436 = _48 ? _435 : _434;
    assign _13 = _436;
    always @(posedge _22) begin
        if (_20)
            _242 <= _50;
        else
            _242 <= _13;
    end
    assign _496 = { _565,
                    _242 };
    assign _493 = _491 * _562;
    assign _494 = _493[63:0];
    assign _497 = _494 + _496;
    always @* begin
        case (_229)
        0:
            _230 <= _60;
        1:
            _230 <= _61;
        2:
            _230 <= _62;
        3:
            _230 <= _63;
        4:
            _230 <= _64;
        5:
            _230 <= _65;
        6:
            _230 <= _66;
        7:
            _230 <= _67;
        8:
            _230 <= _68;
        9:
            _230 <= _69;
        10:
            _230 <= _70;
        11:
            _230 <= _71;
        12:
            _230 <= _72;
        13:
            _230 <= _73;
        14:
            _230 <= _74;
        15:
            _230 <= _75;
        16:
            _230 <= _76;
        17:
            _230 <= _77;
        18:
            _230 <= _78;
        19:
            _230 <= _79;
        20:
            _230 <= _80;
        21:
            _230 <= _81;
        22:
            _230 <= _82;
        23:
            _230 <= _83;
        24:
            _230 <= _84;
        25:
            _230 <= _85;
        26:
            _230 <= _86;
        27:
            _230 <= _87;
        28:
            _230 <= _88;
        29:
            _230 <= _89;
        30:
            _230 <= _90;
        31:
            _230 <= _91;
        32:
            _230 <= _92;
        33:
            _230 <= _93;
        34:
            _230 <= _94;
        35:
            _230 <= _95;
        36:
            _230 <= _96;
        37:
            _230 <= _97;
        38:
            _230 <= _98;
        39:
            _230 <= _99;
        40:
            _230 <= _100;
        41:
            _230 <= _101;
        42:
            _230 <= _102;
        43:
            _230 <= _103;
        44:
            _230 <= _104;
        45:
            _230 <= _105;
        46:
            _230 <= _106;
        47:
            _230 <= _107;
        48:
            _230 <= _108;
        49:
            _230 <= _109;
        50:
            _230 <= _110;
        51:
            _230 <= _111;
        52:
            _230 <= _112;
        53:
            _230 <= _113;
        54:
            _230 <= _114;
        55:
            _230 <= _115;
        56:
            _230 <= _116;
        57:
            _230 <= _117;
        58:
            _230 <= _118;
        59:
            _230 <= _119;
        60:
            _230 <= _120;
        61:
            _230 <= _121;
        62:
            _230 <= _122;
        63:
            _230 <= _123;
        64:
            _230 <= _124;
        65:
            _230 <= _125;
        66:
            _230 <= _126;
        67:
            _230 <= _127;
        68:
            _230 <= _128;
        69:
            _230 <= _129;
        70:
            _230 <= _130;
        71:
            _230 <= _131;
        72:
            _230 <= _132;
        73:
            _230 <= _133;
        74:
            _230 <= _134;
        75:
            _230 <= _135;
        76:
            _230 <= _136;
        77:
            _230 <= _137;
        78:
            _230 <= _138;
        79:
            _230 <= _139;
        80:
            _230 <= _140;
        81:
            _230 <= _141;
        82:
            _230 <= _142;
        83:
            _230 <= _143;
        84:
            _230 <= _144;
        85:
            _230 <= _145;
        86:
            _230 <= _146;
        87:
            _230 <= _147;
        88:
            _230 <= _148;
        89:
            _230 <= _149;
        90:
            _230 <= _150;
        91:
            _230 <= _151;
        92:
            _230 <= _152;
        93:
            _230 <= _153;
        94:
            _230 <= _154;
        95:
            _230 <= _155;
        96:
            _230 <= _156;
        97:
            _230 <= _157;
        98:
            _230 <= _158;
        99:
            _230 <= _159;
        100:
            _230 <= _160;
        101:
            _230 <= _161;
        102:
            _230 <= _162;
        103:
            _230 <= _163;
        104:
            _230 <= _164;
        105:
            _230 <= _165;
        106:
            _230 <= _166;
        107:
            _230 <= _167;
        108:
            _230 <= _168;
        109:
            _230 <= _169;
        110:
            _230 <= _170;
        111:
            _230 <= _171;
        112:
            _230 <= _172;
        113:
            _230 <= _173;
        114:
            _230 <= _174;
        115:
            _230 <= _175;
        116:
            _230 <= _176;
        117:
            _230 <= _177;
        118:
            _230 <= _178;
        119:
            _230 <= _179;
        120:
            _230 <= _180;
        121:
            _230 <= _181;
        122:
            _230 <= _182;
        123:
            _230 <= _183;
        124:
            _230 <= _184;
        125:
            _230 <= _185;
        126:
            _230 <= _186;
        default:
            _230 <= _187;
        endcase
    end
    assign _234 = _230 < _233;
    assign _235 = ~ _234;
    assign _225 = _50 < _194;
    assign _236 = _225 & _235;
    assign _443 = _236 ? _230 : _233;
    assign _187 = _15[511:508];
    assign _186 = _15[507:504];
    assign _185 = _15[503:500];
    assign _184 = _15[499:496];
    assign _183 = _15[495:492];
    assign _182 = _15[491:488];
    assign _181 = _15[487:484];
    assign _180 = _15[483:480];
    assign _179 = _15[479:476];
    assign _178 = _15[475:472];
    assign _177 = _15[471:468];
    assign _176 = _15[467:464];
    assign _175 = _15[463:460];
    assign _174 = _15[459:456];
    assign _173 = _15[455:452];
    assign _172 = _15[451:448];
    assign _171 = _15[447:444];
    assign _170 = _15[443:440];
    assign _169 = _15[439:436];
    assign _168 = _15[435:432];
    assign _167 = _15[431:428];
    assign _166 = _15[427:424];
    assign _165 = _15[423:420];
    assign _164 = _15[419:416];
    assign _163 = _15[415:412];
    assign _162 = _15[411:408];
    assign _161 = _15[407:404];
    assign _160 = _15[403:400];
    assign _159 = _15[399:396];
    assign _158 = _15[395:392];
    assign _157 = _15[391:388];
    assign _156 = _15[387:384];
    assign _155 = _15[383:380];
    assign _154 = _15[379:376];
    assign _153 = _15[375:372];
    assign _152 = _15[371:368];
    assign _151 = _15[367:364];
    assign _150 = _15[363:360];
    assign _149 = _15[359:356];
    assign _148 = _15[355:352];
    assign _147 = _15[351:348];
    assign _146 = _15[347:344];
    assign _145 = _15[343:340];
    assign _144 = _15[339:336];
    assign _143 = _15[335:332];
    assign _142 = _15[331:328];
    assign _141 = _15[327:324];
    assign _140 = _15[323:320];
    assign _139 = _15[319:316];
    assign _138 = _15[315:312];
    assign _137 = _15[311:308];
    assign _136 = _15[307:304];
    assign _135 = _15[303:300];
    assign _134 = _15[299:296];
    assign _133 = _15[295:292];
    assign _132 = _15[291:288];
    assign _131 = _15[287:284];
    assign _130 = _15[283:280];
    assign _129 = _15[279:276];
    assign _128 = _15[275:272];
    assign _127 = _15[271:268];
    assign _126 = _15[267:264];
    assign _125 = _15[263:260];
    assign _124 = _15[259:256];
    assign _123 = _15[255:252];
    assign _122 = _15[251:248];
    assign _121 = _15[247:244];
    assign _120 = _15[243:240];
    assign _119 = _15[239:236];
    assign _118 = _15[235:232];
    assign _117 = _15[231:228];
    assign _116 = _15[227:224];
    assign _115 = _15[223:220];
    assign _114 = _15[219:216];
    assign _113 = _15[215:212];
    assign _112 = _15[211:208];
    assign _111 = _15[207:204];
    assign _110 = _15[203:200];
    assign _109 = _15[199:196];
    assign _108 = _15[195:192];
    assign _107 = _15[191:188];
    assign _106 = _15[187:184];
    assign _105 = _15[183:180];
    assign _104 = _15[179:176];
    assign _103 = _15[175:172];
    assign _102 = _15[171:168];
    assign _101 = _15[167:164];
    assign _100 = _15[163:160];
    assign _99 = _15[159:156];
    assign _98 = _15[155:152];
    assign _97 = _15[151:148];
    assign _96 = _15[147:144];
    assign _95 = _15[143:140];
    assign _94 = _15[139:136];
    assign _93 = _15[135:132];
    assign _92 = _15[131:128];
    assign _91 = _15[127:124];
    assign _90 = _15[123:120];
    assign _89 = _15[119:116];
    assign _88 = _15[115:112];
    assign _87 = _15[111:108];
    assign _86 = _15[107:104];
    assign _85 = _15[103:100];
    assign _84 = _15[99:96];
    assign _83 = _15[95:92];
    assign _82 = _15[91:88];
    assign _81 = _15[87:84];
    assign _80 = _15[83:80];
    assign _79 = _15[79:76];
    assign _78 = _15[75:72];
    assign _77 = _15[71:68];
    assign _76 = _15[67:64];
    assign _75 = _15[63:60];
    assign _74 = _15[59:56];
    assign _73 = _15[55:52];
    assign _72 = _15[51:48];
    assign _71 = _15[47:44];
    assign _70 = _15[43:40];
    assign _69 = _15[39:36];
    assign _68 = _15[35:32];
    assign _67 = _15[31:28];
    assign _66 = _15[27:24];
    assign _65 = _15[23:20];
    assign _64 = _15[19:16];
    assign _63 = _15[15:12];
    assign _62 = _15[11:8];
    assign _61 = _15[7:4];
    assign _15 = data;
    assign _60 = _15[3:0];
    always @* begin
        case (_57)
        0:
            _440 <= _60;
        1:
            _440 <= _61;
        2:
            _440 <= _62;
        3:
            _440 <= _63;
        4:
            _440 <= _64;
        5:
            _440 <= _65;
        6:
            _440 <= _66;
        7:
            _440 <= _67;
        8:
            _440 <= _68;
        9:
            _440 <= _69;
        10:
            _440 <= _70;
        11:
            _440 <= _71;
        12:
            _440 <= _72;
        13:
            _440 <= _73;
        14:
            _440 <= _74;
        15:
            _440 <= _75;
        16:
            _440 <= _76;
        17:
            _440 <= _77;
        18:
            _440 <= _78;
        19:
            _440 <= _79;
        20:
            _440 <= _80;
        21:
            _440 <= _81;
        22:
            _440 <= _82;
        23:
            _440 <= _83;
        24:
            _440 <= _84;
        25:
            _440 <= _85;
        26:
            _440 <= _86;
        27:
            _440 <= _87;
        28:
            _440 <= _88;
        29:
            _440 <= _89;
        30:
            _440 <= _90;
        31:
            _440 <= _91;
        32:
            _440 <= _92;
        33:
            _440 <= _93;
        34:
            _440 <= _94;
        35:
            _440 <= _95;
        36:
            _440 <= _96;
        37:
            _440 <= _97;
        38:
            _440 <= _98;
        39:
            _440 <= _99;
        40:
            _440 <= _100;
        41:
            _440 <= _101;
        42:
            _440 <= _102;
        43:
            _440 <= _103;
        44:
            _440 <= _104;
        45:
            _440 <= _105;
        46:
            _440 <= _106;
        47:
            _440 <= _107;
        48:
            _440 <= _108;
        49:
            _440 <= _109;
        50:
            _440 <= _110;
        51:
            _440 <= _111;
        52:
            _440 <= _112;
        53:
            _440 <= _113;
        54:
            _440 <= _114;
        55:
            _440 <= _115;
        56:
            _440 <= _116;
        57:
            _440 <= _117;
        58:
            _440 <= _118;
        59:
            _440 <= _119;
        60:
            _440 <= _120;
        61:
            _440 <= _121;
        62:
            _440 <= _122;
        63:
            _440 <= _123;
        64:
            _440 <= _124;
        65:
            _440 <= _125;
        66:
            _440 <= _126;
        67:
            _440 <= _127;
        68:
            _440 <= _128;
        69:
            _440 <= _129;
        70:
            _440 <= _130;
        71:
            _440 <= _131;
        72:
            _440 <= _132;
        73:
            _440 <= _133;
        74:
            _440 <= _134;
        75:
            _440 <= _135;
        76:
            _440 <= _136;
        77:
            _440 <= _137;
        78:
            _440 <= _138;
        79:
            _440 <= _139;
        80:
            _440 <= _140;
        81:
            _440 <= _141;
        82:
            _440 <= _142;
        83:
            _440 <= _143;
        84:
            _440 <= _144;
        85:
            _440 <= _145;
        86:
            _440 <= _146;
        87:
            _440 <= _147;
        88:
            _440 <= _148;
        89:
            _440 <= _149;
        90:
            _440 <= _150;
        91:
            _440 <= _151;
        92:
            _440 <= _152;
        93:
            _440 <= _153;
        94:
            _440 <= _154;
        95:
            _440 <= _155;
        96:
            _440 <= _156;
        97:
            _440 <= _157;
        98:
            _440 <= _158;
        99:
            _440 <= _159;
        100:
            _440 <= _160;
        101:
            _440 <= _161;
        102:
            _440 <= _162;
        103:
            _440 <= _163;
        104:
            _440 <= _164;
        105:
            _440 <= _165;
        106:
            _440 <= _166;
        107:
            _440 <= _167;
        108:
            _440 <= _168;
        109:
            _440 <= _169;
        110:
            _440 <= _170;
        111:
            _440 <= _171;
        112:
            _440 <= _172;
        113:
            _440 <= _173;
        114:
            _440 <= _174;
        115:
            _440 <= _175;
        116:
            _440 <= _176;
        117:
            _440 <= _177;
        118:
            _440 <= _178;
        119:
            _440 <= _179;
        120:
            _440 <= _180;
        121:
            _440 <= _181;
        122:
            _440 <= _182;
        123:
            _440 <= _183;
        124:
            _440 <= _184;
        125:
            _440 <= _185;
        126:
            _440 <= _186;
        default:
            _440 <= _187;
        endcase
    end
    assign _438 = _50 < _25;
    assign _441 = _438 ? _440 : _50;
    assign _442 = _40 ? _441 : _233;
    assign _444 = _48 ? _443 : _442;
    assign _16 = _444;
    always @(posedge _22) begin
        if (_20)
            _233 <= _50;
        else
            _233 <= _16;
    end
    assign _490 = { _565,
                    _233 };
    assign _488 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign _487 = _50 < _194;
    assign _491 = _487 ? _490 : _488;
    assign _485 = _221 < _194;
    assign _498 = _485 ? _497 : _491;
    assign _483 = _218 < _194;
    assign _505 = _483 ? _504 : _498;
    assign _481 = _215 < _194;
    assign _512 = _481 ? _511 : _505;
    assign _479 = _212 < _194;
    assign _519 = _479 ? _518 : _512;
    assign _477 = _209 < _194;
    assign _526 = _477 ? _525 : _519;
    assign _475 = _206 < _194;
    assign _533 = _475 ? _532 : _526;
    assign _473 = _203 < _194;
    assign _540 = _473 ? _539 : _533;
    assign _471 = _200 < _194;
    assign _547 = _471 ? _546 : _540;
    assign _469 = _197 < _194;
    assign _554 = _469 ? _553 : _547;
    assign _467 = _191 < _194;
    assign _561 = _467 ? _560 : _554;
    assign _18 = start;
    assign _35 = 2'b10;
    assign _36 = _34 == _35;
    assign _37 = 2'b00;
    assign _459 = 2'b01;
    assign _457 = 8'b00000000;
    assign vdd = 1'b1;
    assign _20 = clear;
    assign _22 = clock;
    assign _449 = _229 - _430;
    assign _446 = _57 - _430;
    assign _447 = _40 ? _446 : _229;
    assign _450 = _48 ? _449 : _447;
    assign _23 = _450;
    always @(posedge _22) begin
        if (_20)
            _229 <= _457;
        else
            _229 <= _23;
    end
    assign _458 = _229 == _457;
    assign _461 = _458 ? _35 : _459;
    assign _25 = k;
    assign _56 = { _50,
                   _25 };
    assign _27 = length;
    assign _57 = _27 - _56;
    assign _452 = _57 == _457;
    assign _455 = _452 ? _35 : _459;
    assign _456 = _40 ? _455 : _34;
    assign _48 = _34 == _459;
    assign _462 = _48 ? _461 : _456;
    assign _28 = _462;
    always @(posedge _22) begin
        if (_20)
            _34 <= _37;
        else
            _34 <= _28;
    end
    assign _38 = _34 == _37;
    assign _39 = _38 | _36;
    assign _40 = _39 & _18;
    assign _463 = _40 ? _25 : _194;
    assign _29 = _463;
    always @(posedge _22) begin
        if (_20)
            _194 <= _50;
        else
            _194 <= _29;
    end
    assign _465 = _328 < _194;
    assign _568 = _465 ? _567 : _561;
    assign result = _568;
    assign done_ = _43;

endmodule
