module day7_opt_a (
    row_bits,
    row_last,
    clear,
    clock,
    width,
    row_valid,
    load,
    ready,
    done_,
    part1_result,
    part2_result,
    state
);

    input [255:0] row_bits;
    input row_last;
    input clear;
    input clock;
    input [7:0] width;
    input row_valid;
    input load;
    output ready;
    output done_;
    output [63:0] part1_result;
    output [63:0] part2_result;
    output [2:0] state;

    wire [63:0] _1099;
    reg [63:0] _1089;
    wire [63:0] _1090;
    wire _317;
    wire [63:0] _1091;
    wire [63:0] _1093;
    wire [63:0] _1095;
    wire [63:0] _2;
    reg [63:0] _320;
    wire [63:0] _1101;
    wire [63:0] _1103;
    wire [63:0] _3;
    reg [63:0] _1100;
    wire [63:0] _6252;
    wire [63:0] _6253;
    wire _1374;
    wire _1373;
    wire _1372;
    wire _1371;
    wire _1370;
    wire _1369;
    wire _1368;
    wire _1367;
    wire _1366;
    wire _1365;
    wire _1364;
    wire _1363;
    wire _1362;
    wire _1361;
    wire _1360;
    wire _1359;
    wire _1358;
    wire _1357;
    wire _1356;
    wire _1355;
    wire _1354;
    wire _1353;
    wire _1352;
    wire _1351;
    wire _1350;
    wire _1349;
    wire _1348;
    wire _1347;
    wire _1346;
    wire _1345;
    wire _1344;
    wire _1343;
    wire _1342;
    wire _1341;
    wire _1340;
    wire _1339;
    wire _1338;
    wire _1337;
    wire _1336;
    wire _1335;
    wire _1334;
    wire _1333;
    wire _1332;
    wire _1331;
    wire _1330;
    wire _1329;
    wire _1328;
    wire _1327;
    wire _1326;
    wire _1325;
    wire _1324;
    wire _1323;
    wire _1322;
    wire _1321;
    wire _1320;
    wire _1319;
    wire _1318;
    wire _1317;
    wire _1316;
    wire _1315;
    wire _1314;
    wire _1313;
    wire _1312;
    wire _1311;
    wire _1310;
    wire _1309;
    wire _1308;
    wire _1307;
    wire _1306;
    wire _1305;
    wire _1304;
    wire _1303;
    wire _1302;
    wire _1301;
    wire _1300;
    wire _1299;
    wire _1298;
    wire _1297;
    wire _1296;
    wire _1295;
    wire _1294;
    wire _1293;
    wire _1292;
    wire _1291;
    wire _1290;
    wire _1289;
    wire _1288;
    wire _1287;
    wire _1286;
    wire _1285;
    wire _1284;
    wire _1283;
    wire _1282;
    wire _1281;
    wire _1280;
    wire _1279;
    wire _1278;
    wire _1277;
    wire _1276;
    wire _1275;
    wire _1274;
    wire _1273;
    wire _1272;
    wire _1271;
    wire _1270;
    wire _1269;
    wire _1268;
    wire _1267;
    wire _1266;
    wire _1265;
    wire _1264;
    wire _1263;
    wire _1262;
    wire _1261;
    wire _1260;
    wire _1259;
    wire _1258;
    wire _1257;
    wire _1256;
    wire _1255;
    wire _1254;
    wire _1253;
    wire _1252;
    wire _1251;
    wire _1250;
    wire _1249;
    wire _1248;
    wire _1247;
    wire _1246;
    wire _1245;
    wire _1244;
    wire _1243;
    wire _1242;
    wire _1241;
    wire _1240;
    wire _1239;
    wire _1238;
    wire _1237;
    wire _1236;
    wire _1235;
    wire _1234;
    wire _1233;
    wire _1232;
    wire _1231;
    wire _1230;
    wire _1229;
    wire _1228;
    wire _1227;
    wire _1226;
    wire _1225;
    wire _1224;
    wire _1223;
    wire _1222;
    wire _1221;
    wire _1220;
    wire _1219;
    wire _1218;
    wire _1217;
    wire _1216;
    wire _1215;
    wire _1214;
    wire _1213;
    wire _1212;
    wire _1211;
    wire _1210;
    wire _1209;
    wire _1208;
    wire _1207;
    wire _1206;
    wire _1205;
    wire _1204;
    wire _1203;
    wire _1202;
    wire _1201;
    wire _1200;
    wire _1199;
    wire _1198;
    wire _1197;
    wire _1196;
    wire _1195;
    wire _1194;
    wire _1193;
    wire _1192;
    wire _1191;
    wire _1190;
    wire _1189;
    wire _1188;
    wire _1187;
    wire _1186;
    wire _1185;
    wire _1184;
    wire _1183;
    wire _1182;
    wire _1181;
    wire _1180;
    wire _1179;
    wire _1178;
    wire _1177;
    wire _1176;
    wire _1175;
    wire _1174;
    wire _1173;
    wire _1172;
    wire _1171;
    wire _1170;
    wire _1169;
    wire _1168;
    wire _1167;
    wire _1166;
    wire _1165;
    wire _1164;
    wire _1163;
    wire _1162;
    wire _1161;
    wire _1160;
    wire _1159;
    wire _1158;
    wire _1157;
    wire _1156;
    wire _1155;
    wire _1154;
    wire _1153;
    wire _1152;
    wire _1151;
    wire _1150;
    wire _1149;
    wire _1148;
    wire _1147;
    wire _1146;
    wire _1145;
    wire _1144;
    wire _1143;
    wire _1142;
    wire _1141;
    wire _1140;
    wire _1139;
    wire _1138;
    wire _1137;
    wire _1136;
    wire _1135;
    wire _1134;
    wire _1133;
    wire _1132;
    wire _1131;
    wire _1130;
    wire _1129;
    wire _1128;
    wire _1127;
    wire _1126;
    wire _1125;
    wire _1124;
    wire _1123;
    wire _1122;
    wire _1121;
    wire _1120;
    wire [255:0] _1108;
    wire [255:0] _6;
    wire [255:0] _1110;
    wire [255:0] _1112;
    wire [255:0] _7;
    reg [255:0] _1109;
    wire _1119;
    reg _1375;
    wire [7:0] _6243;
    wire _6244;
    wire [63:0] _6247;
    wire [7:0] _6224;
    wire _6225;
    wire [63:0] _6228;
    wire [7:0] _1398;
    wire _1399;
    wire [63:0] _1402;
    wire _1388;
    wire _1389;
    wire [63:0] _1392;
    wire _1383;
    wire _1384;
    wire [63:0] _1395;
    wire _1378;
    wire _1379;
    wire [63:0] _1397;
    wire [63:0] _1403;
    wire [63:0] _8;
    reg [63:0] _1088;
    wire [7:0] _1417;
    wire _1418;
    wire [63:0] _1421;
    wire _1411;
    wire _1412;
    wire [63:0] _1413;
    wire _1408;
    wire _1409;
    wire [63:0] _1414;
    wire _1405;
    wire _1406;
    wire [63:0] _1416;
    wire [63:0] _1422;
    wire [63:0] _9;
    reg [63:0] _1085;
    wire [7:0] _1436;
    wire _1437;
    wire [63:0] _1440;
    wire _1430;
    wire _1431;
    wire [63:0] _1432;
    wire _1427;
    wire _1428;
    wire [63:0] _1433;
    wire _1424;
    wire _1425;
    wire [63:0] _1435;
    wire [63:0] _1441;
    wire [63:0] _10;
    reg [63:0] _1082;
    wire [7:0] _1455;
    wire _1456;
    wire [63:0] _1459;
    wire _1449;
    wire _1450;
    wire [63:0] _1451;
    wire _1446;
    wire _1447;
    wire [63:0] _1452;
    wire _1443;
    wire _1444;
    wire [63:0] _1454;
    wire [63:0] _1460;
    wire [63:0] _11;
    reg [63:0] _1079;
    wire [7:0] _1474;
    wire _1475;
    wire [63:0] _1478;
    wire _1468;
    wire _1469;
    wire [63:0] _1470;
    wire _1465;
    wire _1466;
    wire [63:0] _1471;
    wire _1462;
    wire _1463;
    wire [63:0] _1473;
    wire [63:0] _1479;
    wire [63:0] _12;
    reg [63:0] _1076;
    wire [7:0] _1493;
    wire _1494;
    wire [63:0] _1497;
    wire _1487;
    wire _1488;
    wire [63:0] _1489;
    wire _1484;
    wire _1485;
    wire [63:0] _1490;
    wire _1481;
    wire _1482;
    wire [63:0] _1492;
    wire [63:0] _1498;
    wire [63:0] _13;
    reg [63:0] _1073;
    wire [7:0] _1512;
    wire _1513;
    wire [63:0] _1516;
    wire _1506;
    wire _1507;
    wire [63:0] _1508;
    wire _1503;
    wire _1504;
    wire [63:0] _1509;
    wire _1500;
    wire _1501;
    wire [63:0] _1511;
    wire [63:0] _1517;
    wire [63:0] _14;
    reg [63:0] _1070;
    wire [7:0] _1531;
    wire _1532;
    wire [63:0] _1535;
    wire _1525;
    wire _1526;
    wire [63:0] _1527;
    wire _1522;
    wire _1523;
    wire [63:0] _1528;
    wire _1519;
    wire _1520;
    wire [63:0] _1530;
    wire [63:0] _1536;
    wire [63:0] _15;
    reg [63:0] _1067;
    wire [7:0] _1550;
    wire _1551;
    wire [63:0] _1554;
    wire _1544;
    wire _1545;
    wire [63:0] _1546;
    wire _1541;
    wire _1542;
    wire [63:0] _1547;
    wire _1538;
    wire _1539;
    wire [63:0] _1549;
    wire [63:0] _1555;
    wire [63:0] _16;
    reg [63:0] _1064;
    wire [7:0] _1569;
    wire _1570;
    wire [63:0] _1573;
    wire _1563;
    wire _1564;
    wire [63:0] _1565;
    wire _1560;
    wire _1561;
    wire [63:0] _1566;
    wire _1557;
    wire _1558;
    wire [63:0] _1568;
    wire [63:0] _1574;
    wire [63:0] _17;
    reg [63:0] _1061;
    wire [7:0] _1588;
    wire _1589;
    wire [63:0] _1592;
    wire _1582;
    wire _1583;
    wire [63:0] _1584;
    wire _1579;
    wire _1580;
    wire [63:0] _1585;
    wire _1576;
    wire _1577;
    wire [63:0] _1587;
    wire [63:0] _1593;
    wire [63:0] _18;
    reg [63:0] _1058;
    wire [7:0] _1607;
    wire _1608;
    wire [63:0] _1611;
    wire _1601;
    wire _1602;
    wire [63:0] _1603;
    wire _1598;
    wire _1599;
    wire [63:0] _1604;
    wire _1595;
    wire _1596;
    wire [63:0] _1606;
    wire [63:0] _1612;
    wire [63:0] _19;
    reg [63:0] _1055;
    wire [7:0] _1626;
    wire _1627;
    wire [63:0] _1630;
    wire _1620;
    wire _1621;
    wire [63:0] _1622;
    wire _1617;
    wire _1618;
    wire [63:0] _1623;
    wire _1614;
    wire _1615;
    wire [63:0] _1625;
    wire [63:0] _1631;
    wire [63:0] _20;
    reg [63:0] _1052;
    wire [7:0] _1645;
    wire _1646;
    wire [63:0] _1649;
    wire _1639;
    wire _1640;
    wire [63:0] _1641;
    wire _1636;
    wire _1637;
    wire [63:0] _1642;
    wire _1633;
    wire _1634;
    wire [63:0] _1644;
    wire [63:0] _1650;
    wire [63:0] _21;
    reg [63:0] _1049;
    wire [7:0] _1664;
    wire _1665;
    wire [63:0] _1668;
    wire _1658;
    wire _1659;
    wire [63:0] _1660;
    wire _1655;
    wire _1656;
    wire [63:0] _1661;
    wire _1652;
    wire _1653;
    wire [63:0] _1663;
    wire [63:0] _1669;
    wire [63:0] _22;
    reg [63:0] _1046;
    wire [7:0] _1683;
    wire _1684;
    wire [63:0] _1687;
    wire _1677;
    wire _1678;
    wire [63:0] _1679;
    wire _1674;
    wire _1675;
    wire [63:0] _1680;
    wire _1671;
    wire _1672;
    wire [63:0] _1682;
    wire [63:0] _1688;
    wire [63:0] _23;
    reg [63:0] _1043;
    wire [7:0] _1702;
    wire _1703;
    wire [63:0] _1706;
    wire _1696;
    wire _1697;
    wire [63:0] _1698;
    wire _1693;
    wire _1694;
    wire [63:0] _1699;
    wire _1690;
    wire _1691;
    wire [63:0] _1701;
    wire [63:0] _1707;
    wire [63:0] _24;
    reg [63:0] _1040;
    wire [7:0] _1721;
    wire _1722;
    wire [63:0] _1725;
    wire _1715;
    wire _1716;
    wire [63:0] _1717;
    wire _1712;
    wire _1713;
    wire [63:0] _1718;
    wire _1709;
    wire _1710;
    wire [63:0] _1720;
    wire [63:0] _1726;
    wire [63:0] _25;
    reg [63:0] _1037;
    wire [7:0] _1740;
    wire _1741;
    wire [63:0] _1744;
    wire _1734;
    wire _1735;
    wire [63:0] _1736;
    wire _1731;
    wire _1732;
    wire [63:0] _1737;
    wire _1728;
    wire _1729;
    wire [63:0] _1739;
    wire [63:0] _1745;
    wire [63:0] _26;
    reg [63:0] _1034;
    wire [7:0] _1759;
    wire _1760;
    wire [63:0] _1763;
    wire _1753;
    wire _1754;
    wire [63:0] _1755;
    wire _1750;
    wire _1751;
    wire [63:0] _1756;
    wire _1747;
    wire _1748;
    wire [63:0] _1758;
    wire [63:0] _1764;
    wire [63:0] _27;
    reg [63:0] _1031;
    wire [7:0] _1778;
    wire _1779;
    wire [63:0] _1782;
    wire _1772;
    wire _1773;
    wire [63:0] _1774;
    wire _1769;
    wire _1770;
    wire [63:0] _1775;
    wire _1766;
    wire _1767;
    wire [63:0] _1777;
    wire [63:0] _1783;
    wire [63:0] _28;
    reg [63:0] _1028;
    wire [7:0] _1797;
    wire _1798;
    wire [63:0] _1801;
    wire _1791;
    wire _1792;
    wire [63:0] _1793;
    wire _1788;
    wire _1789;
    wire [63:0] _1794;
    wire _1785;
    wire _1786;
    wire [63:0] _1796;
    wire [63:0] _1802;
    wire [63:0] _29;
    reg [63:0] _1025;
    wire [7:0] _1816;
    wire _1817;
    wire [63:0] _1820;
    wire _1810;
    wire _1811;
    wire [63:0] _1812;
    wire _1807;
    wire _1808;
    wire [63:0] _1813;
    wire _1804;
    wire _1805;
    wire [63:0] _1815;
    wire [63:0] _1821;
    wire [63:0] _30;
    reg [63:0] _1022;
    wire [7:0] _1835;
    wire _1836;
    wire [63:0] _1839;
    wire _1829;
    wire _1830;
    wire [63:0] _1831;
    wire _1826;
    wire _1827;
    wire [63:0] _1832;
    wire _1823;
    wire _1824;
    wire [63:0] _1834;
    wire [63:0] _1840;
    wire [63:0] _31;
    reg [63:0] _1019;
    wire [7:0] _1854;
    wire _1855;
    wire [63:0] _1858;
    wire _1848;
    wire _1849;
    wire [63:0] _1850;
    wire _1845;
    wire _1846;
    wire [63:0] _1851;
    wire _1842;
    wire _1843;
    wire [63:0] _1853;
    wire [63:0] _1859;
    wire [63:0] _32;
    reg [63:0] _1016;
    wire [7:0] _1873;
    wire _1874;
    wire [63:0] _1877;
    wire _1867;
    wire _1868;
    wire [63:0] _1869;
    wire _1864;
    wire _1865;
    wire [63:0] _1870;
    wire _1861;
    wire _1862;
    wire [63:0] _1872;
    wire [63:0] _1878;
    wire [63:0] _33;
    reg [63:0] _1013;
    wire [7:0] _1892;
    wire _1893;
    wire [63:0] _1896;
    wire _1886;
    wire _1887;
    wire [63:0] _1888;
    wire _1883;
    wire _1884;
    wire [63:0] _1889;
    wire _1880;
    wire _1881;
    wire [63:0] _1891;
    wire [63:0] _1897;
    wire [63:0] _34;
    reg [63:0] _1010;
    wire [7:0] _1911;
    wire _1912;
    wire [63:0] _1915;
    wire _1905;
    wire _1906;
    wire [63:0] _1907;
    wire _1902;
    wire _1903;
    wire [63:0] _1908;
    wire _1899;
    wire _1900;
    wire [63:0] _1910;
    wire [63:0] _1916;
    wire [63:0] _35;
    reg [63:0] _1007;
    wire [7:0] _1930;
    wire _1931;
    wire [63:0] _1934;
    wire _1924;
    wire _1925;
    wire [63:0] _1926;
    wire _1921;
    wire _1922;
    wire [63:0] _1927;
    wire _1918;
    wire _1919;
    wire [63:0] _1929;
    wire [63:0] _1935;
    wire [63:0] _36;
    reg [63:0] _1004;
    wire [7:0] _1949;
    wire _1950;
    wire [63:0] _1953;
    wire _1943;
    wire _1944;
    wire [63:0] _1945;
    wire _1940;
    wire _1941;
    wire [63:0] _1946;
    wire _1937;
    wire _1938;
    wire [63:0] _1948;
    wire [63:0] _1954;
    wire [63:0] _37;
    reg [63:0] _1001;
    wire [7:0] _1968;
    wire _1969;
    wire [63:0] _1972;
    wire _1962;
    wire _1963;
    wire [63:0] _1964;
    wire _1959;
    wire _1960;
    wire [63:0] _1965;
    wire _1956;
    wire _1957;
    wire [63:0] _1967;
    wire [63:0] _1973;
    wire [63:0] _38;
    reg [63:0] _998;
    wire [7:0] _1987;
    wire _1988;
    wire [63:0] _1991;
    wire _1981;
    wire _1982;
    wire [63:0] _1983;
    wire _1978;
    wire _1979;
    wire [63:0] _1984;
    wire _1975;
    wire _1976;
    wire [63:0] _1986;
    wire [63:0] _1992;
    wire [63:0] _39;
    reg [63:0] _995;
    wire [7:0] _2006;
    wire _2007;
    wire [63:0] _2010;
    wire _2000;
    wire _2001;
    wire [63:0] _2002;
    wire _1997;
    wire _1998;
    wire [63:0] _2003;
    wire _1994;
    wire _1995;
    wire [63:0] _2005;
    wire [63:0] _2011;
    wire [63:0] _40;
    reg [63:0] _992;
    wire [7:0] _2025;
    wire _2026;
    wire [63:0] _2029;
    wire _2019;
    wire _2020;
    wire [63:0] _2021;
    wire _2016;
    wire _2017;
    wire [63:0] _2022;
    wire _2013;
    wire _2014;
    wire [63:0] _2024;
    wire [63:0] _2030;
    wire [63:0] _41;
    reg [63:0] _989;
    wire [7:0] _2044;
    wire _2045;
    wire [63:0] _2048;
    wire _2038;
    wire _2039;
    wire [63:0] _2040;
    wire _2035;
    wire _2036;
    wire [63:0] _2041;
    wire _2032;
    wire _2033;
    wire [63:0] _2043;
    wire [63:0] _2049;
    wire [63:0] _42;
    reg [63:0] _986;
    wire [7:0] _2063;
    wire _2064;
    wire [63:0] _2067;
    wire _2057;
    wire _2058;
    wire [63:0] _2059;
    wire _2054;
    wire _2055;
    wire [63:0] _2060;
    wire _2051;
    wire _2052;
    wire [63:0] _2062;
    wire [63:0] _2068;
    wire [63:0] _43;
    reg [63:0] _983;
    wire [7:0] _2082;
    wire _2083;
    wire [63:0] _2086;
    wire _2076;
    wire _2077;
    wire [63:0] _2078;
    wire _2073;
    wire _2074;
    wire [63:0] _2079;
    wire _2070;
    wire _2071;
    wire [63:0] _2081;
    wire [63:0] _2087;
    wire [63:0] _44;
    reg [63:0] _980;
    wire [7:0] _2101;
    wire _2102;
    wire [63:0] _2105;
    wire _2095;
    wire _2096;
    wire [63:0] _2097;
    wire _2092;
    wire _2093;
    wire [63:0] _2098;
    wire _2089;
    wire _2090;
    wire [63:0] _2100;
    wire [63:0] _2106;
    wire [63:0] _45;
    reg [63:0] _977;
    wire [7:0] _2120;
    wire _2121;
    wire [63:0] _2124;
    wire _2114;
    wire _2115;
    wire [63:0] _2116;
    wire _2111;
    wire _2112;
    wire [63:0] _2117;
    wire _2108;
    wire _2109;
    wire [63:0] _2119;
    wire [63:0] _2125;
    wire [63:0] _46;
    reg [63:0] _974;
    wire [7:0] _2139;
    wire _2140;
    wire [63:0] _2143;
    wire _2133;
    wire _2134;
    wire [63:0] _2135;
    wire _2130;
    wire _2131;
    wire [63:0] _2136;
    wire _2127;
    wire _2128;
    wire [63:0] _2138;
    wire [63:0] _2144;
    wire [63:0] _47;
    reg [63:0] _971;
    wire [7:0] _2158;
    wire _2159;
    wire [63:0] _2162;
    wire _2152;
    wire _2153;
    wire [63:0] _2154;
    wire _2149;
    wire _2150;
    wire [63:0] _2155;
    wire _2146;
    wire _2147;
    wire [63:0] _2157;
    wire [63:0] _2163;
    wire [63:0] _48;
    reg [63:0] _968;
    wire [7:0] _2177;
    wire _2178;
    wire [63:0] _2181;
    wire _2171;
    wire _2172;
    wire [63:0] _2173;
    wire _2168;
    wire _2169;
    wire [63:0] _2174;
    wire _2165;
    wire _2166;
    wire [63:0] _2176;
    wire [63:0] _2182;
    wire [63:0] _49;
    reg [63:0] _965;
    wire [7:0] _2196;
    wire _2197;
    wire [63:0] _2200;
    wire _2190;
    wire _2191;
    wire [63:0] _2192;
    wire _2187;
    wire _2188;
    wire [63:0] _2193;
    wire _2184;
    wire _2185;
    wire [63:0] _2195;
    wire [63:0] _2201;
    wire [63:0] _50;
    reg [63:0] _962;
    wire [7:0] _2215;
    wire _2216;
    wire [63:0] _2219;
    wire _2209;
    wire _2210;
    wire [63:0] _2211;
    wire _2206;
    wire _2207;
    wire [63:0] _2212;
    wire _2203;
    wire _2204;
    wire [63:0] _2214;
    wire [63:0] _2220;
    wire [63:0] _51;
    reg [63:0] _959;
    wire [7:0] _2234;
    wire _2235;
    wire [63:0] _2238;
    wire _2228;
    wire _2229;
    wire [63:0] _2230;
    wire _2225;
    wire _2226;
    wire [63:0] _2231;
    wire _2222;
    wire _2223;
    wire [63:0] _2233;
    wire [63:0] _2239;
    wire [63:0] _52;
    reg [63:0] _956;
    wire [7:0] _2253;
    wire _2254;
    wire [63:0] _2257;
    wire _2247;
    wire _2248;
    wire [63:0] _2249;
    wire _2244;
    wire _2245;
    wire [63:0] _2250;
    wire _2241;
    wire _2242;
    wire [63:0] _2252;
    wire [63:0] _2258;
    wire [63:0] _53;
    reg [63:0] _953;
    wire [7:0] _2272;
    wire _2273;
    wire [63:0] _2276;
    wire _2266;
    wire _2267;
    wire [63:0] _2268;
    wire _2263;
    wire _2264;
    wire [63:0] _2269;
    wire _2260;
    wire _2261;
    wire [63:0] _2271;
    wire [63:0] _2277;
    wire [63:0] _54;
    reg [63:0] _950;
    wire [7:0] _2291;
    wire _2292;
    wire [63:0] _2295;
    wire _2285;
    wire _2286;
    wire [63:0] _2287;
    wire _2282;
    wire _2283;
    wire [63:0] _2288;
    wire _2279;
    wire _2280;
    wire [63:0] _2290;
    wire [63:0] _2296;
    wire [63:0] _55;
    reg [63:0] _947;
    wire [7:0] _2310;
    wire _2311;
    wire [63:0] _2314;
    wire _2304;
    wire _2305;
    wire [63:0] _2306;
    wire _2301;
    wire _2302;
    wire [63:0] _2307;
    wire _2298;
    wire _2299;
    wire [63:0] _2309;
    wire [63:0] _2315;
    wire [63:0] _56;
    reg [63:0] _944;
    wire [7:0] _2329;
    wire _2330;
    wire [63:0] _2333;
    wire _2323;
    wire _2324;
    wire [63:0] _2325;
    wire _2320;
    wire _2321;
    wire [63:0] _2326;
    wire _2317;
    wire _2318;
    wire [63:0] _2328;
    wire [63:0] _2334;
    wire [63:0] _57;
    reg [63:0] _941;
    wire [7:0] _2348;
    wire _2349;
    wire [63:0] _2352;
    wire _2342;
    wire _2343;
    wire [63:0] _2344;
    wire _2339;
    wire _2340;
    wire [63:0] _2345;
    wire _2336;
    wire _2337;
    wire [63:0] _2347;
    wire [63:0] _2353;
    wire [63:0] _58;
    reg [63:0] _938;
    wire [7:0] _2367;
    wire _2368;
    wire [63:0] _2371;
    wire _2361;
    wire _2362;
    wire [63:0] _2363;
    wire _2358;
    wire _2359;
    wire [63:0] _2364;
    wire _2355;
    wire _2356;
    wire [63:0] _2366;
    wire [63:0] _2372;
    wire [63:0] _59;
    reg [63:0] _935;
    wire [7:0] _2386;
    wire _2387;
    wire [63:0] _2390;
    wire _2380;
    wire _2381;
    wire [63:0] _2382;
    wire _2377;
    wire _2378;
    wire [63:0] _2383;
    wire _2374;
    wire _2375;
    wire [63:0] _2385;
    wire [63:0] _2391;
    wire [63:0] _60;
    reg [63:0] _932;
    wire [7:0] _2405;
    wire _2406;
    wire [63:0] _2409;
    wire _2399;
    wire _2400;
    wire [63:0] _2401;
    wire _2396;
    wire _2397;
    wire [63:0] _2402;
    wire _2393;
    wire _2394;
    wire [63:0] _2404;
    wire [63:0] _2410;
    wire [63:0] _61;
    reg [63:0] _929;
    wire [7:0] _2424;
    wire _2425;
    wire [63:0] _2428;
    wire _2418;
    wire _2419;
    wire [63:0] _2420;
    wire _2415;
    wire _2416;
    wire [63:0] _2421;
    wire _2412;
    wire _2413;
    wire [63:0] _2423;
    wire [63:0] _2429;
    wire [63:0] _62;
    reg [63:0] _926;
    wire [7:0] _2443;
    wire _2444;
    wire [63:0] _2447;
    wire _2437;
    wire _2438;
    wire [63:0] _2439;
    wire _2434;
    wire _2435;
    wire [63:0] _2440;
    wire _2431;
    wire _2432;
    wire [63:0] _2442;
    wire [63:0] _2448;
    wire [63:0] _63;
    reg [63:0] _923;
    wire [7:0] _2462;
    wire _2463;
    wire [63:0] _2466;
    wire _2456;
    wire _2457;
    wire [63:0] _2458;
    wire _2453;
    wire _2454;
    wire [63:0] _2459;
    wire _2450;
    wire _2451;
    wire [63:0] _2461;
    wire [63:0] _2467;
    wire [63:0] _64;
    reg [63:0] _920;
    wire [7:0] _2481;
    wire _2482;
    wire [63:0] _2485;
    wire _2475;
    wire _2476;
    wire [63:0] _2477;
    wire _2472;
    wire _2473;
    wire [63:0] _2478;
    wire _2469;
    wire _2470;
    wire [63:0] _2480;
    wire [63:0] _2486;
    wire [63:0] _65;
    reg [63:0] _917;
    wire [7:0] _2500;
    wire _2501;
    wire [63:0] _2504;
    wire _2494;
    wire _2495;
    wire [63:0] _2496;
    wire _2491;
    wire _2492;
    wire [63:0] _2497;
    wire _2488;
    wire _2489;
    wire [63:0] _2499;
    wire [63:0] _2505;
    wire [63:0] _66;
    reg [63:0] _914;
    wire [7:0] _2519;
    wire _2520;
    wire [63:0] _2523;
    wire _2513;
    wire _2514;
    wire [63:0] _2515;
    wire _2510;
    wire _2511;
    wire [63:0] _2516;
    wire _2507;
    wire _2508;
    wire [63:0] _2518;
    wire [63:0] _2524;
    wire [63:0] _67;
    reg [63:0] _911;
    wire [7:0] _2538;
    wire _2539;
    wire [63:0] _2542;
    wire _2532;
    wire _2533;
    wire [63:0] _2534;
    wire _2529;
    wire _2530;
    wire [63:0] _2535;
    wire _2526;
    wire _2527;
    wire [63:0] _2537;
    wire [63:0] _2543;
    wire [63:0] _68;
    reg [63:0] _908;
    wire [7:0] _2557;
    wire _2558;
    wire [63:0] _2561;
    wire _2551;
    wire _2552;
    wire [63:0] _2553;
    wire _2548;
    wire _2549;
    wire [63:0] _2554;
    wire _2545;
    wire _2546;
    wire [63:0] _2556;
    wire [63:0] _2562;
    wire [63:0] _69;
    reg [63:0] _905;
    wire [7:0] _2576;
    wire _2577;
    wire [63:0] _2580;
    wire _2570;
    wire _2571;
    wire [63:0] _2572;
    wire _2567;
    wire _2568;
    wire [63:0] _2573;
    wire _2564;
    wire _2565;
    wire [63:0] _2575;
    wire [63:0] _2581;
    wire [63:0] _70;
    reg [63:0] _902;
    wire [7:0] _2595;
    wire _2596;
    wire [63:0] _2599;
    wire _2589;
    wire _2590;
    wire [63:0] _2591;
    wire _2586;
    wire _2587;
    wire [63:0] _2592;
    wire _2583;
    wire _2584;
    wire [63:0] _2594;
    wire [63:0] _2600;
    wire [63:0] _71;
    reg [63:0] _899;
    wire [7:0] _2614;
    wire _2615;
    wire [63:0] _2618;
    wire _2608;
    wire _2609;
    wire [63:0] _2610;
    wire _2605;
    wire _2606;
    wire [63:0] _2611;
    wire _2602;
    wire _2603;
    wire [63:0] _2613;
    wire [63:0] _2619;
    wire [63:0] _72;
    reg [63:0] _896;
    wire [7:0] _2633;
    wire _2634;
    wire [63:0] _2637;
    wire _2627;
    wire _2628;
    wire [63:0] _2629;
    wire _2624;
    wire _2625;
    wire [63:0] _2630;
    wire _2621;
    wire _2622;
    wire [63:0] _2632;
    wire [63:0] _2638;
    wire [63:0] _73;
    reg [63:0] _893;
    wire [7:0] _2652;
    wire _2653;
    wire [63:0] _2656;
    wire _2646;
    wire _2647;
    wire [63:0] _2648;
    wire _2643;
    wire _2644;
    wire [63:0] _2649;
    wire _2640;
    wire _2641;
    wire [63:0] _2651;
    wire [63:0] _2657;
    wire [63:0] _74;
    reg [63:0] _890;
    wire [7:0] _2671;
    wire _2672;
    wire [63:0] _2675;
    wire _2665;
    wire _2666;
    wire [63:0] _2667;
    wire _2662;
    wire _2663;
    wire [63:0] _2668;
    wire _2659;
    wire _2660;
    wire [63:0] _2670;
    wire [63:0] _2676;
    wire [63:0] _75;
    reg [63:0] _887;
    wire [7:0] _2690;
    wire _2691;
    wire [63:0] _2694;
    wire _2684;
    wire _2685;
    wire [63:0] _2686;
    wire _2681;
    wire _2682;
    wire [63:0] _2687;
    wire _2678;
    wire _2679;
    wire [63:0] _2689;
    wire [63:0] _2695;
    wire [63:0] _76;
    reg [63:0] _884;
    wire [7:0] _2709;
    wire _2710;
    wire [63:0] _2713;
    wire _2703;
    wire _2704;
    wire [63:0] _2705;
    wire _2700;
    wire _2701;
    wire [63:0] _2706;
    wire _2697;
    wire _2698;
    wire [63:0] _2708;
    wire [63:0] _2714;
    wire [63:0] _77;
    reg [63:0] _881;
    wire [7:0] _2728;
    wire _2729;
    wire [63:0] _2732;
    wire _2722;
    wire _2723;
    wire [63:0] _2724;
    wire _2719;
    wire _2720;
    wire [63:0] _2725;
    wire _2716;
    wire _2717;
    wire [63:0] _2727;
    wire [63:0] _2733;
    wire [63:0] _78;
    reg [63:0] _878;
    wire [7:0] _2747;
    wire _2748;
    wire [63:0] _2751;
    wire _2741;
    wire _2742;
    wire [63:0] _2743;
    wire _2738;
    wire _2739;
    wire [63:0] _2744;
    wire _2735;
    wire _2736;
    wire [63:0] _2746;
    wire [63:0] _2752;
    wire [63:0] _79;
    reg [63:0] _875;
    wire [7:0] _2766;
    wire _2767;
    wire [63:0] _2770;
    wire _2760;
    wire _2761;
    wire [63:0] _2762;
    wire _2757;
    wire _2758;
    wire [63:0] _2763;
    wire _2754;
    wire _2755;
    wire [63:0] _2765;
    wire [63:0] _2771;
    wire [63:0] _80;
    reg [63:0] _872;
    wire [7:0] _2785;
    wire _2786;
    wire [63:0] _2789;
    wire _2779;
    wire _2780;
    wire [63:0] _2781;
    wire _2776;
    wire _2777;
    wire [63:0] _2782;
    wire _2773;
    wire _2774;
    wire [63:0] _2784;
    wire [63:0] _2790;
    wire [63:0] _81;
    reg [63:0] _869;
    wire [7:0] _2804;
    wire _2805;
    wire [63:0] _2808;
    wire _2798;
    wire _2799;
    wire [63:0] _2800;
    wire _2795;
    wire _2796;
    wire [63:0] _2801;
    wire _2792;
    wire _2793;
    wire [63:0] _2803;
    wire [63:0] _2809;
    wire [63:0] _82;
    reg [63:0] _866;
    wire [7:0] _2823;
    wire _2824;
    wire [63:0] _2827;
    wire _2817;
    wire _2818;
    wire [63:0] _2819;
    wire _2814;
    wire _2815;
    wire [63:0] _2820;
    wire _2811;
    wire _2812;
    wire [63:0] _2822;
    wire [63:0] _2828;
    wire [63:0] _83;
    reg [63:0] _863;
    wire [7:0] _2842;
    wire _2843;
    wire [63:0] _2846;
    wire _2836;
    wire _2837;
    wire [63:0] _2838;
    wire _2833;
    wire _2834;
    wire [63:0] _2839;
    wire _2830;
    wire _2831;
    wire [63:0] _2841;
    wire [63:0] _2847;
    wire [63:0] _84;
    reg [63:0] _860;
    wire [7:0] _2861;
    wire _2862;
    wire [63:0] _2865;
    wire _2855;
    wire _2856;
    wire [63:0] _2857;
    wire _2852;
    wire _2853;
    wire [63:0] _2858;
    wire _2849;
    wire _2850;
    wire [63:0] _2860;
    wire [63:0] _2866;
    wire [63:0] _85;
    reg [63:0] _857;
    wire [7:0] _2880;
    wire _2881;
    wire [63:0] _2884;
    wire _2874;
    wire _2875;
    wire [63:0] _2876;
    wire _2871;
    wire _2872;
    wire [63:0] _2877;
    wire _2868;
    wire _2869;
    wire [63:0] _2879;
    wire [63:0] _2885;
    wire [63:0] _86;
    reg [63:0] _854;
    wire [7:0] _2899;
    wire _2900;
    wire [63:0] _2903;
    wire _2893;
    wire _2894;
    wire [63:0] _2895;
    wire _2890;
    wire _2891;
    wire [63:0] _2896;
    wire _2887;
    wire _2888;
    wire [63:0] _2898;
    wire [63:0] _2904;
    wire [63:0] _87;
    reg [63:0] _851;
    wire [7:0] _2918;
    wire _2919;
    wire [63:0] _2922;
    wire _2912;
    wire _2913;
    wire [63:0] _2914;
    wire _2909;
    wire _2910;
    wire [63:0] _2915;
    wire _2906;
    wire _2907;
    wire [63:0] _2917;
    wire [63:0] _2923;
    wire [63:0] _88;
    reg [63:0] _848;
    wire [7:0] _2937;
    wire _2938;
    wire [63:0] _2941;
    wire _2931;
    wire _2932;
    wire [63:0] _2933;
    wire _2928;
    wire _2929;
    wire [63:0] _2934;
    wire _2925;
    wire _2926;
    wire [63:0] _2936;
    wire [63:0] _2942;
    wire [63:0] _89;
    reg [63:0] _845;
    wire [7:0] _2956;
    wire _2957;
    wire [63:0] _2960;
    wire _2950;
    wire _2951;
    wire [63:0] _2952;
    wire _2947;
    wire _2948;
    wire [63:0] _2953;
    wire _2944;
    wire _2945;
    wire [63:0] _2955;
    wire [63:0] _2961;
    wire [63:0] _90;
    reg [63:0] _842;
    wire [7:0] _2975;
    wire _2976;
    wire [63:0] _2979;
    wire _2969;
    wire _2970;
    wire [63:0] _2971;
    wire _2966;
    wire _2967;
    wire [63:0] _2972;
    wire _2963;
    wire _2964;
    wire [63:0] _2974;
    wire [63:0] _2980;
    wire [63:0] _91;
    reg [63:0] _839;
    wire [7:0] _2994;
    wire _2995;
    wire [63:0] _2998;
    wire _2988;
    wire _2989;
    wire [63:0] _2990;
    wire _2985;
    wire _2986;
    wire [63:0] _2991;
    wire _2982;
    wire _2983;
    wire [63:0] _2993;
    wire [63:0] _2999;
    wire [63:0] _92;
    reg [63:0] _836;
    wire [7:0] _3013;
    wire _3014;
    wire [63:0] _3017;
    wire _3007;
    wire _3008;
    wire [63:0] _3009;
    wire _3004;
    wire _3005;
    wire [63:0] _3010;
    wire _3001;
    wire _3002;
    wire [63:0] _3012;
    wire [63:0] _3018;
    wire [63:0] _93;
    reg [63:0] _833;
    wire [7:0] _3032;
    wire _3033;
    wire [63:0] _3036;
    wire _3026;
    wire _3027;
    wire [63:0] _3028;
    wire _3023;
    wire _3024;
    wire [63:0] _3029;
    wire _3020;
    wire _3021;
    wire [63:0] _3031;
    wire [63:0] _3037;
    wire [63:0] _94;
    reg [63:0] _830;
    wire [7:0] _3051;
    wire _3052;
    wire [63:0] _3055;
    wire _3045;
    wire _3046;
    wire [63:0] _3047;
    wire _3042;
    wire _3043;
    wire [63:0] _3048;
    wire _3039;
    wire _3040;
    wire [63:0] _3050;
    wire [63:0] _3056;
    wire [63:0] _95;
    reg [63:0] _827;
    wire [7:0] _3070;
    wire _3071;
    wire [63:0] _3074;
    wire _3064;
    wire _3065;
    wire [63:0] _3066;
    wire _3061;
    wire _3062;
    wire [63:0] _3067;
    wire _3058;
    wire _3059;
    wire [63:0] _3069;
    wire [63:0] _3075;
    wire [63:0] _96;
    reg [63:0] _824;
    wire [7:0] _3089;
    wire _3090;
    wire [63:0] _3093;
    wire _3083;
    wire _3084;
    wire [63:0] _3085;
    wire _3080;
    wire _3081;
    wire [63:0] _3086;
    wire _3077;
    wire _3078;
    wire [63:0] _3088;
    wire [63:0] _3094;
    wire [63:0] _97;
    reg [63:0] _821;
    wire [7:0] _3108;
    wire _3109;
    wire [63:0] _3112;
    wire _3102;
    wire _3103;
    wire [63:0] _3104;
    wire _3099;
    wire _3100;
    wire [63:0] _3105;
    wire _3096;
    wire _3097;
    wire [63:0] _3107;
    wire [63:0] _3113;
    wire [63:0] _98;
    reg [63:0] _818;
    wire [7:0] _3127;
    wire _3128;
    wire [63:0] _3131;
    wire _3121;
    wire _3122;
    wire [63:0] _3123;
    wire _3118;
    wire _3119;
    wire [63:0] _3124;
    wire _3115;
    wire _3116;
    wire [63:0] _3126;
    wire [63:0] _3132;
    wire [63:0] _99;
    reg [63:0] _815;
    wire [7:0] _3146;
    wire _3147;
    wire [63:0] _3150;
    wire _3140;
    wire _3141;
    wire [63:0] _3142;
    wire _3137;
    wire _3138;
    wire [63:0] _3143;
    wire _3134;
    wire _3135;
    wire [63:0] _3145;
    wire [63:0] _3151;
    wire [63:0] _100;
    reg [63:0] _812;
    wire [7:0] _3165;
    wire _3166;
    wire [63:0] _3169;
    wire _3159;
    wire _3160;
    wire [63:0] _3161;
    wire _3156;
    wire _3157;
    wire [63:0] _3162;
    wire _3153;
    wire _3154;
    wire [63:0] _3164;
    wire [63:0] _3170;
    wire [63:0] _101;
    reg [63:0] _809;
    wire [7:0] _3184;
    wire _3185;
    wire [63:0] _3188;
    wire _3178;
    wire _3179;
    wire [63:0] _3180;
    wire _3175;
    wire _3176;
    wire [63:0] _3181;
    wire _3172;
    wire _3173;
    wire [63:0] _3183;
    wire [63:0] _3189;
    wire [63:0] _102;
    reg [63:0] _806;
    wire [7:0] _3203;
    wire _3204;
    wire [63:0] _3207;
    wire _3197;
    wire _3198;
    wire [63:0] _3199;
    wire _3194;
    wire _3195;
    wire [63:0] _3200;
    wire _3191;
    wire _3192;
    wire [63:0] _3202;
    wire [63:0] _3208;
    wire [63:0] _103;
    reg [63:0] _803;
    wire [7:0] _3222;
    wire _3223;
    wire [63:0] _3226;
    wire _3216;
    wire _3217;
    wire [63:0] _3218;
    wire _3213;
    wire _3214;
    wire [63:0] _3219;
    wire _3210;
    wire _3211;
    wire [63:0] _3221;
    wire [63:0] _3227;
    wire [63:0] _104;
    reg [63:0] _800;
    wire [7:0] _3241;
    wire _3242;
    wire [63:0] _3245;
    wire _3235;
    wire _3236;
    wire [63:0] _3237;
    wire _3232;
    wire _3233;
    wire [63:0] _3238;
    wire _3229;
    wire _3230;
    wire [63:0] _3240;
    wire [63:0] _3246;
    wire [63:0] _105;
    reg [63:0] _797;
    wire [7:0] _3260;
    wire _3261;
    wire [63:0] _3264;
    wire _3254;
    wire _3255;
    wire [63:0] _3256;
    wire _3251;
    wire _3252;
    wire [63:0] _3257;
    wire _3248;
    wire _3249;
    wire [63:0] _3259;
    wire [63:0] _3265;
    wire [63:0] _106;
    reg [63:0] _794;
    wire [7:0] _3279;
    wire _3280;
    wire [63:0] _3283;
    wire _3273;
    wire _3274;
    wire [63:0] _3275;
    wire _3270;
    wire _3271;
    wire [63:0] _3276;
    wire _3267;
    wire _3268;
    wire [63:0] _3278;
    wire [63:0] _3284;
    wire [63:0] _107;
    reg [63:0] _791;
    wire [7:0] _3298;
    wire _3299;
    wire [63:0] _3302;
    wire _3292;
    wire _3293;
    wire [63:0] _3294;
    wire _3289;
    wire _3290;
    wire [63:0] _3295;
    wire _3286;
    wire _3287;
    wire [63:0] _3297;
    wire [63:0] _3303;
    wire [63:0] _108;
    reg [63:0] _788;
    wire [7:0] _3317;
    wire _3318;
    wire [63:0] _3321;
    wire _3311;
    wire _3312;
    wire [63:0] _3313;
    wire _3308;
    wire _3309;
    wire [63:0] _3314;
    wire _3305;
    wire _3306;
    wire [63:0] _3316;
    wire [63:0] _3322;
    wire [63:0] _109;
    reg [63:0] _785;
    wire [7:0] _3336;
    wire _3337;
    wire [63:0] _3340;
    wire _3330;
    wire _3331;
    wire [63:0] _3332;
    wire _3327;
    wire _3328;
    wire [63:0] _3333;
    wire _3324;
    wire _3325;
    wire [63:0] _3335;
    wire [63:0] _3341;
    wire [63:0] _110;
    reg [63:0] _782;
    wire [7:0] _3355;
    wire _3356;
    wire [63:0] _3359;
    wire _3349;
    wire _3350;
    wire [63:0] _3351;
    wire _3346;
    wire _3347;
    wire [63:0] _3352;
    wire _3343;
    wire _3344;
    wire [63:0] _3354;
    wire [63:0] _3360;
    wire [63:0] _111;
    reg [63:0] _779;
    wire [7:0] _3374;
    wire _3375;
    wire [63:0] _3378;
    wire _3368;
    wire _3369;
    wire [63:0] _3370;
    wire _3365;
    wire _3366;
    wire [63:0] _3371;
    wire _3362;
    wire _3363;
    wire [63:0] _3373;
    wire [63:0] _3379;
    wire [63:0] _112;
    reg [63:0] _776;
    wire [7:0] _3393;
    wire _3394;
    wire [63:0] _3397;
    wire _3387;
    wire _3388;
    wire [63:0] _3389;
    wire _3384;
    wire _3385;
    wire [63:0] _3390;
    wire _3381;
    wire _3382;
    wire [63:0] _3392;
    wire [63:0] _3398;
    wire [63:0] _113;
    reg [63:0] _773;
    wire [7:0] _3412;
    wire _3413;
    wire [63:0] _3416;
    wire _3406;
    wire _3407;
    wire [63:0] _3408;
    wire _3403;
    wire _3404;
    wire [63:0] _3409;
    wire _3400;
    wire _3401;
    wire [63:0] _3411;
    wire [63:0] _3417;
    wire [63:0] _114;
    reg [63:0] _770;
    wire [7:0] _3431;
    wire _3432;
    wire [63:0] _3435;
    wire _3425;
    wire _3426;
    wire [63:0] _3427;
    wire _3422;
    wire _3423;
    wire [63:0] _3428;
    wire _3419;
    wire _3420;
    wire [63:0] _3430;
    wire [63:0] _3436;
    wire [63:0] _115;
    reg [63:0] _767;
    wire [7:0] _3450;
    wire _3451;
    wire [63:0] _3454;
    wire _3444;
    wire _3445;
    wire [63:0] _3446;
    wire _3441;
    wire _3442;
    wire [63:0] _3447;
    wire _3438;
    wire _3439;
    wire [63:0] _3449;
    wire [63:0] _3455;
    wire [63:0] _116;
    reg [63:0] _764;
    wire [7:0] _3469;
    wire _3470;
    wire [63:0] _3473;
    wire _3463;
    wire _3464;
    wire [63:0] _3465;
    wire _3460;
    wire _3461;
    wire [63:0] _3466;
    wire _3457;
    wire _3458;
    wire [63:0] _3468;
    wire [63:0] _3474;
    wire [63:0] _117;
    reg [63:0] _761;
    wire [7:0] _3488;
    wire _3489;
    wire [63:0] _3492;
    wire _3482;
    wire _3483;
    wire [63:0] _3484;
    wire _3479;
    wire _3480;
    wire [63:0] _3485;
    wire _3476;
    wire _3477;
    wire [63:0] _3487;
    wire [63:0] _3493;
    wire [63:0] _118;
    reg [63:0] _758;
    wire [7:0] _3507;
    wire _3508;
    wire [63:0] _3511;
    wire _3501;
    wire _3502;
    wire [63:0] _3503;
    wire _3498;
    wire _3499;
    wire [63:0] _3504;
    wire _3495;
    wire _3496;
    wire [63:0] _3506;
    wire [63:0] _3512;
    wire [63:0] _119;
    reg [63:0] _755;
    wire [7:0] _3526;
    wire _3527;
    wire [63:0] _3530;
    wire _3520;
    wire _3521;
    wire [63:0] _3522;
    wire _3517;
    wire _3518;
    wire [63:0] _3523;
    wire _3514;
    wire _3515;
    wire [63:0] _3525;
    wire [63:0] _3531;
    wire [63:0] _120;
    reg [63:0] _752;
    wire [7:0] _3545;
    wire _3546;
    wire [63:0] _3549;
    wire _3539;
    wire _3540;
    wire [63:0] _3541;
    wire _3536;
    wire _3537;
    wire [63:0] _3542;
    wire _3533;
    wire _3534;
    wire [63:0] _3544;
    wire [63:0] _3550;
    wire [63:0] _121;
    reg [63:0] _749;
    wire [7:0] _3564;
    wire _3565;
    wire [63:0] _3568;
    wire _3558;
    wire _3559;
    wire [63:0] _3560;
    wire _3555;
    wire _3556;
    wire [63:0] _3561;
    wire _3552;
    wire _3553;
    wire [63:0] _3563;
    wire [63:0] _3569;
    wire [63:0] _122;
    reg [63:0] _746;
    wire [7:0] _3583;
    wire _3584;
    wire [63:0] _3587;
    wire _3577;
    wire _3578;
    wire [63:0] _3579;
    wire _3574;
    wire _3575;
    wire [63:0] _3580;
    wire _3571;
    wire _3572;
    wire [63:0] _3582;
    wire [63:0] _3588;
    wire [63:0] _123;
    reg [63:0] _743;
    wire [7:0] _3602;
    wire _3603;
    wire [63:0] _3606;
    wire _3596;
    wire _3597;
    wire [63:0] _3598;
    wire _3593;
    wire _3594;
    wire [63:0] _3599;
    wire _3590;
    wire _3591;
    wire [63:0] _3601;
    wire [63:0] _3607;
    wire [63:0] _124;
    reg [63:0] _740;
    wire [7:0] _3621;
    wire _3622;
    wire [63:0] _3625;
    wire _3615;
    wire _3616;
    wire [63:0] _3617;
    wire _3612;
    wire _3613;
    wire [63:0] _3618;
    wire _3609;
    wire _3610;
    wire [63:0] _3620;
    wire [63:0] _3626;
    wire [63:0] _125;
    reg [63:0] _737;
    wire [7:0] _3640;
    wire _3641;
    wire [63:0] _3644;
    wire _3634;
    wire _3635;
    wire [63:0] _3636;
    wire _3631;
    wire _3632;
    wire [63:0] _3637;
    wire _3628;
    wire _3629;
    wire [63:0] _3639;
    wire [63:0] _3645;
    wire [63:0] _126;
    reg [63:0] _734;
    wire [7:0] _3659;
    wire _3660;
    wire [63:0] _3663;
    wire _3653;
    wire _3654;
    wire [63:0] _3655;
    wire _3650;
    wire _3651;
    wire [63:0] _3656;
    wire _3647;
    wire _3648;
    wire [63:0] _3658;
    wire [63:0] _3664;
    wire [63:0] _127;
    reg [63:0] _731;
    wire [7:0] _3678;
    wire _3679;
    wire [63:0] _3682;
    wire _3672;
    wire _3673;
    wire [63:0] _3674;
    wire _3669;
    wire _3670;
    wire [63:0] _3675;
    wire _3666;
    wire _3667;
    wire [63:0] _3677;
    wire [63:0] _3683;
    wire [63:0] _128;
    reg [63:0] _728;
    wire [7:0] _3697;
    wire _3698;
    wire [63:0] _3701;
    wire _3691;
    wire _3692;
    wire [63:0] _3693;
    wire _3688;
    wire _3689;
    wire [63:0] _3694;
    wire _3685;
    wire _3686;
    wire [63:0] _3696;
    wire [63:0] _3702;
    wire [63:0] _129;
    reg [63:0] _725;
    wire [7:0] _3716;
    wire _3717;
    wire [63:0] _3720;
    wire _3710;
    wire _3711;
    wire [63:0] _3712;
    wire _3707;
    wire _3708;
    wire [63:0] _3713;
    wire _3704;
    wire _3705;
    wire [63:0] _3715;
    wire [63:0] _3721;
    wire [63:0] _130;
    reg [63:0] _722;
    wire [7:0] _3735;
    wire _3736;
    wire [63:0] _3739;
    wire _3729;
    wire _3730;
    wire [63:0] _3731;
    wire _3726;
    wire _3727;
    wire [63:0] _3732;
    wire _3723;
    wire _3724;
    wire [63:0] _3734;
    wire [63:0] _3740;
    wire [63:0] _131;
    reg [63:0] _719;
    wire [7:0] _3754;
    wire _3755;
    wire [63:0] _3758;
    wire _3748;
    wire _3749;
    wire [63:0] _3750;
    wire _3745;
    wire _3746;
    wire [63:0] _3751;
    wire _3742;
    wire _3743;
    wire [63:0] _3753;
    wire [63:0] _3759;
    wire [63:0] _132;
    reg [63:0] _716;
    wire [7:0] _3773;
    wire _3774;
    wire [63:0] _3777;
    wire _3767;
    wire _3768;
    wire [63:0] _3769;
    wire _3764;
    wire _3765;
    wire [63:0] _3770;
    wire _3761;
    wire _3762;
    wire [63:0] _3772;
    wire [63:0] _3778;
    wire [63:0] _133;
    reg [63:0] _713;
    wire [7:0] _3792;
    wire _3793;
    wire [63:0] _3796;
    wire _3786;
    wire _3787;
    wire [63:0] _3788;
    wire _3783;
    wire _3784;
    wire [63:0] _3789;
    wire _3780;
    wire _3781;
    wire [63:0] _3791;
    wire [63:0] _3797;
    wire [63:0] _134;
    reg [63:0] _710;
    wire [7:0] _3811;
    wire _3812;
    wire [63:0] _3815;
    wire _3805;
    wire _3806;
    wire [63:0] _3807;
    wire _3802;
    wire _3803;
    wire [63:0] _3808;
    wire _3799;
    wire _3800;
    wire [63:0] _3810;
    wire [63:0] _3816;
    wire [63:0] _135;
    reg [63:0] _707;
    wire [7:0] _3830;
    wire _3831;
    wire [63:0] _3834;
    wire _3824;
    wire _3825;
    wire [63:0] _3826;
    wire _3821;
    wire _3822;
    wire [63:0] _3827;
    wire _3818;
    wire _3819;
    wire [63:0] _3829;
    wire [63:0] _3835;
    wire [63:0] _136;
    reg [63:0] _704;
    wire [7:0] _3849;
    wire _3850;
    wire [63:0] _3853;
    wire _3843;
    wire _3844;
    wire [63:0] _3845;
    wire _3840;
    wire _3841;
    wire [63:0] _3846;
    wire _3837;
    wire _3838;
    wire [63:0] _3848;
    wire [63:0] _3854;
    wire [63:0] _137;
    reg [63:0] _701;
    wire [7:0] _3868;
    wire _3869;
    wire [63:0] _3872;
    wire _3862;
    wire _3863;
    wire [63:0] _3864;
    wire _3859;
    wire _3860;
    wire [63:0] _3865;
    wire _3856;
    wire _3857;
    wire [63:0] _3867;
    wire [63:0] _3873;
    wire [63:0] _138;
    reg [63:0] _698;
    wire [7:0] _3887;
    wire _3888;
    wire [63:0] _3891;
    wire _3881;
    wire _3882;
    wire [63:0] _3883;
    wire _3878;
    wire _3879;
    wire [63:0] _3884;
    wire _3875;
    wire _3876;
    wire [63:0] _3886;
    wire [63:0] _3892;
    wire [63:0] _139;
    reg [63:0] _695;
    wire [7:0] _3906;
    wire _3907;
    wire [63:0] _3910;
    wire _3900;
    wire _3901;
    wire [63:0] _3902;
    wire _3897;
    wire _3898;
    wire [63:0] _3903;
    wire _3894;
    wire _3895;
    wire [63:0] _3905;
    wire [63:0] _3911;
    wire [63:0] _140;
    reg [63:0] _692;
    wire [7:0] _3925;
    wire _3926;
    wire [63:0] _3929;
    wire _3919;
    wire _3920;
    wire [63:0] _3921;
    wire _3916;
    wire _3917;
    wire [63:0] _3922;
    wire _3913;
    wire _3914;
    wire [63:0] _3924;
    wire [63:0] _3930;
    wire [63:0] _141;
    reg [63:0] _689;
    wire [7:0] _3944;
    wire _3945;
    wire [63:0] _3948;
    wire _3938;
    wire _3939;
    wire [63:0] _3940;
    wire _3935;
    wire _3936;
    wire [63:0] _3941;
    wire _3932;
    wire _3933;
    wire [63:0] _3943;
    wire [63:0] _3949;
    wire [63:0] _142;
    reg [63:0] _686;
    wire [7:0] _3963;
    wire _3964;
    wire [63:0] _3967;
    wire _3957;
    wire _3958;
    wire [63:0] _3959;
    wire _3954;
    wire _3955;
    wire [63:0] _3960;
    wire _3951;
    wire _3952;
    wire [63:0] _3962;
    wire [63:0] _3968;
    wire [63:0] _143;
    reg [63:0] _683;
    wire [7:0] _3982;
    wire _3983;
    wire [63:0] _3986;
    wire _3976;
    wire _3977;
    wire [63:0] _3978;
    wire _3973;
    wire _3974;
    wire [63:0] _3979;
    wire _3970;
    wire _3971;
    wire [63:0] _3981;
    wire [63:0] _3987;
    wire [63:0] _144;
    reg [63:0] _680;
    wire [7:0] _4001;
    wire _4002;
    wire [63:0] _4005;
    wire _3995;
    wire _3996;
    wire [63:0] _3997;
    wire _3992;
    wire _3993;
    wire [63:0] _3998;
    wire _3989;
    wire _3990;
    wire [63:0] _4000;
    wire [63:0] _4006;
    wire [63:0] _145;
    reg [63:0] _677;
    wire [7:0] _4020;
    wire _4021;
    wire [63:0] _4024;
    wire _4014;
    wire _4015;
    wire [63:0] _4016;
    wire _4011;
    wire _4012;
    wire [63:0] _4017;
    wire _4008;
    wire _4009;
    wire [63:0] _4019;
    wire [63:0] _4025;
    wire [63:0] _146;
    reg [63:0] _674;
    wire [7:0] _4039;
    wire _4040;
    wire [63:0] _4043;
    wire _4033;
    wire _4034;
    wire [63:0] _4035;
    wire _4030;
    wire _4031;
    wire [63:0] _4036;
    wire _4027;
    wire _4028;
    wire [63:0] _4038;
    wire [63:0] _4044;
    wire [63:0] _147;
    reg [63:0] _671;
    wire [7:0] _4058;
    wire _4059;
    wire [63:0] _4062;
    wire _4052;
    wire _4053;
    wire [63:0] _4054;
    wire _4049;
    wire _4050;
    wire [63:0] _4055;
    wire _4046;
    wire _4047;
    wire [63:0] _4057;
    wire [63:0] _4063;
    wire [63:0] _148;
    reg [63:0] _668;
    wire [7:0] _4077;
    wire _4078;
    wire [63:0] _4081;
    wire _4071;
    wire _4072;
    wire [63:0] _4073;
    wire _4068;
    wire _4069;
    wire [63:0] _4074;
    wire _4065;
    wire _4066;
    wire [63:0] _4076;
    wire [63:0] _4082;
    wire [63:0] _149;
    reg [63:0] _665;
    wire [7:0] _4096;
    wire _4097;
    wire [63:0] _4100;
    wire _4090;
    wire _4091;
    wire [63:0] _4092;
    wire _4087;
    wire _4088;
    wire [63:0] _4093;
    wire _4084;
    wire _4085;
    wire [63:0] _4095;
    wire [63:0] _4101;
    wire [63:0] _150;
    reg [63:0] _662;
    wire [7:0] _4115;
    wire _4116;
    wire [63:0] _4119;
    wire _4109;
    wire _4110;
    wire [63:0] _4111;
    wire _4106;
    wire _4107;
    wire [63:0] _4112;
    wire _4103;
    wire _4104;
    wire [63:0] _4114;
    wire [63:0] _4120;
    wire [63:0] _151;
    reg [63:0] _659;
    wire [7:0] _4134;
    wire _4135;
    wire [63:0] _4138;
    wire _4128;
    wire _4129;
    wire [63:0] _4130;
    wire _4125;
    wire _4126;
    wire [63:0] _4131;
    wire _4122;
    wire _4123;
    wire [63:0] _4133;
    wire [63:0] _4139;
    wire [63:0] _152;
    reg [63:0] _656;
    wire [7:0] _4153;
    wire _4154;
    wire [63:0] _4157;
    wire _4147;
    wire _4148;
    wire [63:0] _4149;
    wire _4144;
    wire _4145;
    wire [63:0] _4150;
    wire _4141;
    wire _4142;
    wire [63:0] _4152;
    wire [63:0] _4158;
    wire [63:0] _153;
    reg [63:0] _653;
    wire [7:0] _4172;
    wire _4173;
    wire [63:0] _4176;
    wire _4166;
    wire _4167;
    wire [63:0] _4168;
    wire _4163;
    wire _4164;
    wire [63:0] _4169;
    wire _4160;
    wire _4161;
    wire [63:0] _4171;
    wire [63:0] _4177;
    wire [63:0] _154;
    reg [63:0] _650;
    wire [7:0] _4191;
    wire _4192;
    wire [63:0] _4195;
    wire _4185;
    wire _4186;
    wire [63:0] _4187;
    wire _4182;
    wire _4183;
    wire [63:0] _4188;
    wire _4179;
    wire _4180;
    wire [63:0] _4190;
    wire [63:0] _4196;
    wire [63:0] _155;
    reg [63:0] _647;
    wire [7:0] _4210;
    wire _4211;
    wire [63:0] _4214;
    wire _4204;
    wire _4205;
    wire [63:0] _4206;
    wire _4201;
    wire _4202;
    wire [63:0] _4207;
    wire _4198;
    wire _4199;
    wire [63:0] _4209;
    wire [63:0] _4215;
    wire [63:0] _156;
    reg [63:0] _644;
    wire [7:0] _4229;
    wire _4230;
    wire [63:0] _4233;
    wire _4223;
    wire _4224;
    wire [63:0] _4225;
    wire _4220;
    wire _4221;
    wire [63:0] _4226;
    wire _4217;
    wire _4218;
    wire [63:0] _4228;
    wire [63:0] _4234;
    wire [63:0] _157;
    reg [63:0] _641;
    wire [7:0] _4248;
    wire _4249;
    wire [63:0] _4252;
    wire _4242;
    wire _4243;
    wire [63:0] _4244;
    wire _4239;
    wire _4240;
    wire [63:0] _4245;
    wire _4236;
    wire _4237;
    wire [63:0] _4247;
    wire [63:0] _4253;
    wire [63:0] _158;
    reg [63:0] _638;
    wire [7:0] _4267;
    wire _4268;
    wire [63:0] _4271;
    wire _4261;
    wire _4262;
    wire [63:0] _4263;
    wire _4258;
    wire _4259;
    wire [63:0] _4264;
    wire _4255;
    wire _4256;
    wire [63:0] _4266;
    wire [63:0] _4272;
    wire [63:0] _159;
    reg [63:0] _635;
    wire [7:0] _4286;
    wire _4287;
    wire [63:0] _4290;
    wire _4280;
    wire _4281;
    wire [63:0] _4282;
    wire _4277;
    wire _4278;
    wire [63:0] _4283;
    wire _4274;
    wire _4275;
    wire [63:0] _4285;
    wire [63:0] _4291;
    wire [63:0] _160;
    reg [63:0] _632;
    wire [7:0] _4305;
    wire _4306;
    wire [63:0] _4309;
    wire _4299;
    wire _4300;
    wire [63:0] _4301;
    wire _4296;
    wire _4297;
    wire [63:0] _4302;
    wire _4293;
    wire _4294;
    wire [63:0] _4304;
    wire [63:0] _4310;
    wire [63:0] _161;
    reg [63:0] _629;
    wire [7:0] _4324;
    wire _4325;
    wire [63:0] _4328;
    wire _4318;
    wire _4319;
    wire [63:0] _4320;
    wire _4315;
    wire _4316;
    wire [63:0] _4321;
    wire _4312;
    wire _4313;
    wire [63:0] _4323;
    wire [63:0] _4329;
    wire [63:0] _162;
    reg [63:0] _626;
    wire [7:0] _4343;
    wire _4344;
    wire [63:0] _4347;
    wire _4337;
    wire _4338;
    wire [63:0] _4339;
    wire _4334;
    wire _4335;
    wire [63:0] _4340;
    wire _4331;
    wire _4332;
    wire [63:0] _4342;
    wire [63:0] _4348;
    wire [63:0] _163;
    reg [63:0] _623;
    wire [7:0] _4362;
    wire _4363;
    wire [63:0] _4366;
    wire _4356;
    wire _4357;
    wire [63:0] _4358;
    wire _4353;
    wire _4354;
    wire [63:0] _4359;
    wire _4350;
    wire _4351;
    wire [63:0] _4361;
    wire [63:0] _4367;
    wire [63:0] _164;
    reg [63:0] _620;
    wire [7:0] _4381;
    wire _4382;
    wire [63:0] _4385;
    wire _4375;
    wire _4376;
    wire [63:0] _4377;
    wire _4372;
    wire _4373;
    wire [63:0] _4378;
    wire _4369;
    wire _4370;
    wire [63:0] _4380;
    wire [63:0] _4386;
    wire [63:0] _165;
    reg [63:0] _617;
    wire [7:0] _4400;
    wire _4401;
    wire [63:0] _4404;
    wire _4394;
    wire _4395;
    wire [63:0] _4396;
    wire _4391;
    wire _4392;
    wire [63:0] _4397;
    wire _4388;
    wire _4389;
    wire [63:0] _4399;
    wire [63:0] _4405;
    wire [63:0] _166;
    reg [63:0] _614;
    wire [7:0] _4419;
    wire _4420;
    wire [63:0] _4423;
    wire _4413;
    wire _4414;
    wire [63:0] _4415;
    wire _4410;
    wire _4411;
    wire [63:0] _4416;
    wire _4407;
    wire _4408;
    wire [63:0] _4418;
    wire [63:0] _4424;
    wire [63:0] _167;
    reg [63:0] _611;
    wire [7:0] _4438;
    wire _4439;
    wire [63:0] _4442;
    wire _4432;
    wire _4433;
    wire [63:0] _4434;
    wire _4429;
    wire _4430;
    wire [63:0] _4435;
    wire _4426;
    wire _4427;
    wire [63:0] _4437;
    wire [63:0] _4443;
    wire [63:0] _168;
    reg [63:0] _608;
    wire [7:0] _4457;
    wire _4458;
    wire [63:0] _4461;
    wire _4451;
    wire _4452;
    wire [63:0] _4453;
    wire _4448;
    wire _4449;
    wire [63:0] _4454;
    wire _4445;
    wire _4446;
    wire [63:0] _4456;
    wire [63:0] _4462;
    wire [63:0] _169;
    reg [63:0] _605;
    wire [7:0] _4476;
    wire _4477;
    wire [63:0] _4480;
    wire _4470;
    wire _4471;
    wire [63:0] _4472;
    wire _4467;
    wire _4468;
    wire [63:0] _4473;
    wire _4464;
    wire _4465;
    wire [63:0] _4475;
    wire [63:0] _4481;
    wire [63:0] _170;
    reg [63:0] _602;
    wire [7:0] _4495;
    wire _4496;
    wire [63:0] _4499;
    wire _4489;
    wire _4490;
    wire [63:0] _4491;
    wire _4486;
    wire _4487;
    wire [63:0] _4492;
    wire _4483;
    wire _4484;
    wire [63:0] _4494;
    wire [63:0] _4500;
    wire [63:0] _171;
    reg [63:0] _599;
    wire [7:0] _4514;
    wire _4515;
    wire [63:0] _4518;
    wire _4508;
    wire _4509;
    wire [63:0] _4510;
    wire _4505;
    wire _4506;
    wire [63:0] _4511;
    wire _4502;
    wire _4503;
    wire [63:0] _4513;
    wire [63:0] _4519;
    wire [63:0] _172;
    reg [63:0] _596;
    wire [7:0] _4533;
    wire _4534;
    wire [63:0] _4537;
    wire _4527;
    wire _4528;
    wire [63:0] _4529;
    wire _4524;
    wire _4525;
    wire [63:0] _4530;
    wire _4521;
    wire _4522;
    wire [63:0] _4532;
    wire [63:0] _4538;
    wire [63:0] _173;
    reg [63:0] _593;
    wire [7:0] _4552;
    wire _4553;
    wire [63:0] _4556;
    wire _4546;
    wire _4547;
    wire [63:0] _4548;
    wire _4543;
    wire _4544;
    wire [63:0] _4549;
    wire _4540;
    wire _4541;
    wire [63:0] _4551;
    wire [63:0] _4557;
    wire [63:0] _174;
    reg [63:0] _590;
    wire [7:0] _4571;
    wire _4572;
    wire [63:0] _4575;
    wire _4565;
    wire _4566;
    wire [63:0] _4567;
    wire _4562;
    wire _4563;
    wire [63:0] _4568;
    wire _4559;
    wire _4560;
    wire [63:0] _4570;
    wire [63:0] _4576;
    wire [63:0] _175;
    reg [63:0] _587;
    wire [7:0] _4590;
    wire _4591;
    wire [63:0] _4594;
    wire _4584;
    wire _4585;
    wire [63:0] _4586;
    wire _4581;
    wire _4582;
    wire [63:0] _4587;
    wire _4578;
    wire _4579;
    wire [63:0] _4589;
    wire [63:0] _4595;
    wire [63:0] _176;
    reg [63:0] _584;
    wire [7:0] _4609;
    wire _4610;
    wire [63:0] _4613;
    wire _4603;
    wire _4604;
    wire [63:0] _4605;
    wire _4600;
    wire _4601;
    wire [63:0] _4606;
    wire _4597;
    wire _4598;
    wire [63:0] _4608;
    wire [63:0] _4614;
    wire [63:0] _177;
    reg [63:0] _581;
    wire [7:0] _4628;
    wire _4629;
    wire [63:0] _4632;
    wire _4622;
    wire _4623;
    wire [63:0] _4624;
    wire _4619;
    wire _4620;
    wire [63:0] _4625;
    wire _4616;
    wire _4617;
    wire [63:0] _4627;
    wire [63:0] _4633;
    wire [63:0] _178;
    reg [63:0] _578;
    wire [7:0] _4647;
    wire _4648;
    wire [63:0] _4651;
    wire _4641;
    wire _4642;
    wire [63:0] _4643;
    wire _4638;
    wire _4639;
    wire [63:0] _4644;
    wire _4635;
    wire _4636;
    wire [63:0] _4646;
    wire [63:0] _4652;
    wire [63:0] _179;
    reg [63:0] _575;
    wire [7:0] _4666;
    wire _4667;
    wire [63:0] _4670;
    wire _4660;
    wire _4661;
    wire [63:0] _4662;
    wire _4657;
    wire _4658;
    wire [63:0] _4663;
    wire _4654;
    wire _4655;
    wire [63:0] _4665;
    wire [63:0] _4671;
    wire [63:0] _180;
    reg [63:0] _572;
    wire [7:0] _4685;
    wire _4686;
    wire [63:0] _4689;
    wire _4679;
    wire _4680;
    wire [63:0] _4681;
    wire _4676;
    wire _4677;
    wire [63:0] _4682;
    wire _4673;
    wire _4674;
    wire [63:0] _4684;
    wire [63:0] _4690;
    wire [63:0] _181;
    reg [63:0] _569;
    wire [7:0] _4704;
    wire _4705;
    wire [63:0] _4708;
    wire _4698;
    wire _4699;
    wire [63:0] _4700;
    wire _4695;
    wire _4696;
    wire [63:0] _4701;
    wire _4692;
    wire _4693;
    wire [63:0] _4703;
    wire [63:0] _4709;
    wire [63:0] _182;
    reg [63:0] _566;
    wire [7:0] _4723;
    wire _4724;
    wire [63:0] _4727;
    wire _4717;
    wire _4718;
    wire [63:0] _4719;
    wire _4714;
    wire _4715;
    wire [63:0] _4720;
    wire _4711;
    wire _4712;
    wire [63:0] _4722;
    wire [63:0] _4728;
    wire [63:0] _183;
    reg [63:0] _563;
    wire [7:0] _4742;
    wire _4743;
    wire [63:0] _4746;
    wire _4736;
    wire _4737;
    wire [63:0] _4738;
    wire _4733;
    wire _4734;
    wire [63:0] _4739;
    wire _4730;
    wire _4731;
    wire [63:0] _4741;
    wire [63:0] _4747;
    wire [63:0] _184;
    reg [63:0] _560;
    wire [7:0] _4761;
    wire _4762;
    wire [63:0] _4765;
    wire _4755;
    wire _4756;
    wire [63:0] _4757;
    wire _4752;
    wire _4753;
    wire [63:0] _4758;
    wire _4749;
    wire _4750;
    wire [63:0] _4760;
    wire [63:0] _4766;
    wire [63:0] _185;
    reg [63:0] _557;
    wire [7:0] _4780;
    wire _4781;
    wire [63:0] _4784;
    wire _4774;
    wire _4775;
    wire [63:0] _4776;
    wire _4771;
    wire _4772;
    wire [63:0] _4777;
    wire _4768;
    wire _4769;
    wire [63:0] _4779;
    wire [63:0] _4785;
    wire [63:0] _186;
    reg [63:0] _554;
    wire [7:0] _4799;
    wire _4800;
    wire [63:0] _4803;
    wire _4793;
    wire _4794;
    wire [63:0] _4795;
    wire _4790;
    wire _4791;
    wire [63:0] _4796;
    wire _4787;
    wire _4788;
    wire [63:0] _4798;
    wire [63:0] _4804;
    wire [63:0] _187;
    reg [63:0] _551;
    wire [7:0] _4818;
    wire _4819;
    wire [63:0] _4822;
    wire _4812;
    wire _4813;
    wire [63:0] _4814;
    wire _4809;
    wire _4810;
    wire [63:0] _4815;
    wire _4806;
    wire _4807;
    wire [63:0] _4817;
    wire [63:0] _4823;
    wire [63:0] _188;
    reg [63:0] _548;
    wire [7:0] _4837;
    wire _4838;
    wire [63:0] _4841;
    wire _4831;
    wire _4832;
    wire [63:0] _4833;
    wire _4828;
    wire _4829;
    wire [63:0] _4834;
    wire _4825;
    wire _4826;
    wire [63:0] _4836;
    wire [63:0] _4842;
    wire [63:0] _189;
    reg [63:0] _545;
    wire [7:0] _4856;
    wire _4857;
    wire [63:0] _4860;
    wire _4850;
    wire _4851;
    wire [63:0] _4852;
    wire _4847;
    wire _4848;
    wire [63:0] _4853;
    wire _4844;
    wire _4845;
    wire [63:0] _4855;
    wire [63:0] _4861;
    wire [63:0] _190;
    reg [63:0] _542;
    wire [7:0] _4875;
    wire _4876;
    wire [63:0] _4879;
    wire _4869;
    wire _4870;
    wire [63:0] _4871;
    wire _4866;
    wire _4867;
    wire [63:0] _4872;
    wire _4863;
    wire _4864;
    wire [63:0] _4874;
    wire [63:0] _4880;
    wire [63:0] _191;
    reg [63:0] _539;
    wire [7:0] _4894;
    wire _4895;
    wire [63:0] _4898;
    wire _4888;
    wire _4889;
    wire [63:0] _4890;
    wire _4885;
    wire _4886;
    wire [63:0] _4891;
    wire _4882;
    wire _4883;
    wire [63:0] _4893;
    wire [63:0] _4899;
    wire [63:0] _192;
    reg [63:0] _536;
    wire [7:0] _4913;
    wire _4914;
    wire [63:0] _4917;
    wire _4907;
    wire _4908;
    wire [63:0] _4909;
    wire _4904;
    wire _4905;
    wire [63:0] _4910;
    wire _4901;
    wire _4902;
    wire [63:0] _4912;
    wire [63:0] _4918;
    wire [63:0] _193;
    reg [63:0] _533;
    wire [7:0] _4932;
    wire _4933;
    wire [63:0] _4936;
    wire _4926;
    wire _4927;
    wire [63:0] _4928;
    wire _4923;
    wire _4924;
    wire [63:0] _4929;
    wire _4920;
    wire _4921;
    wire [63:0] _4931;
    wire [63:0] _4937;
    wire [63:0] _194;
    reg [63:0] _530;
    wire [7:0] _4951;
    wire _4952;
    wire [63:0] _4955;
    wire _4945;
    wire _4946;
    wire [63:0] _4947;
    wire _4942;
    wire _4943;
    wire [63:0] _4948;
    wire _4939;
    wire _4940;
    wire [63:0] _4950;
    wire [63:0] _4956;
    wire [63:0] _195;
    reg [63:0] _527;
    wire [7:0] _4970;
    wire _4971;
    wire [63:0] _4974;
    wire _4964;
    wire _4965;
    wire [63:0] _4966;
    wire _4961;
    wire _4962;
    wire [63:0] _4967;
    wire _4958;
    wire _4959;
    wire [63:0] _4969;
    wire [63:0] _4975;
    wire [63:0] _196;
    reg [63:0] _524;
    wire [7:0] _4989;
    wire _4990;
    wire [63:0] _4993;
    wire _4983;
    wire _4984;
    wire [63:0] _4985;
    wire _4980;
    wire _4981;
    wire [63:0] _4986;
    wire _4977;
    wire _4978;
    wire [63:0] _4988;
    wire [63:0] _4994;
    wire [63:0] _197;
    reg [63:0] _521;
    wire [7:0] _5008;
    wire _5009;
    wire [63:0] _5012;
    wire _5002;
    wire _5003;
    wire [63:0] _5004;
    wire _4999;
    wire _5000;
    wire [63:0] _5005;
    wire _4996;
    wire _4997;
    wire [63:0] _5007;
    wire [63:0] _5013;
    wire [63:0] _198;
    reg [63:0] _518;
    wire [7:0] _5027;
    wire _5028;
    wire [63:0] _5031;
    wire _5021;
    wire _5022;
    wire [63:0] _5023;
    wire _5018;
    wire _5019;
    wire [63:0] _5024;
    wire _5015;
    wire _5016;
    wire [63:0] _5026;
    wire [63:0] _5032;
    wire [63:0] _199;
    reg [63:0] _515;
    wire [7:0] _5046;
    wire _5047;
    wire [63:0] _5050;
    wire _5040;
    wire _5041;
    wire [63:0] _5042;
    wire _5037;
    wire _5038;
    wire [63:0] _5043;
    wire _5034;
    wire _5035;
    wire [63:0] _5045;
    wire [63:0] _5051;
    wire [63:0] _200;
    reg [63:0] _512;
    wire [7:0] _5065;
    wire _5066;
    wire [63:0] _5069;
    wire _5059;
    wire _5060;
    wire [63:0] _5061;
    wire _5056;
    wire _5057;
    wire [63:0] _5062;
    wire _5053;
    wire _5054;
    wire [63:0] _5064;
    wire [63:0] _5070;
    wire [63:0] _201;
    reg [63:0] _509;
    wire [7:0] _5084;
    wire _5085;
    wire [63:0] _5088;
    wire _5078;
    wire _5079;
    wire [63:0] _5080;
    wire _5075;
    wire _5076;
    wire [63:0] _5081;
    wire _5072;
    wire _5073;
    wire [63:0] _5083;
    wire [63:0] _5089;
    wire [63:0] _202;
    reg [63:0] _506;
    wire [7:0] _5103;
    wire _5104;
    wire [63:0] _5107;
    wire _5097;
    wire _5098;
    wire [63:0] _5099;
    wire _5094;
    wire _5095;
    wire [63:0] _5100;
    wire _5091;
    wire _5092;
    wire [63:0] _5102;
    wire [63:0] _5108;
    wire [63:0] _203;
    reg [63:0] _503;
    wire [7:0] _5122;
    wire _5123;
    wire [63:0] _5126;
    wire _5116;
    wire _5117;
    wire [63:0] _5118;
    wire _5113;
    wire _5114;
    wire [63:0] _5119;
    wire _5110;
    wire _5111;
    wire [63:0] _5121;
    wire [63:0] _5127;
    wire [63:0] _204;
    reg [63:0] _500;
    wire [7:0] _5141;
    wire _5142;
    wire [63:0] _5145;
    wire _5135;
    wire _5136;
    wire [63:0] _5137;
    wire _5132;
    wire _5133;
    wire [63:0] _5138;
    wire _5129;
    wire _5130;
    wire [63:0] _5140;
    wire [63:0] _5146;
    wire [63:0] _205;
    reg [63:0] _497;
    wire [7:0] _5160;
    wire _5161;
    wire [63:0] _5164;
    wire _5154;
    wire _5155;
    wire [63:0] _5156;
    wire _5151;
    wire _5152;
    wire [63:0] _5157;
    wire _5148;
    wire _5149;
    wire [63:0] _5159;
    wire [63:0] _5165;
    wire [63:0] _206;
    reg [63:0] _494;
    wire [7:0] _5179;
    wire _5180;
    wire [63:0] _5183;
    wire _5173;
    wire _5174;
    wire [63:0] _5175;
    wire _5170;
    wire _5171;
    wire [63:0] _5176;
    wire _5167;
    wire _5168;
    wire [63:0] _5178;
    wire [63:0] _5184;
    wire [63:0] _207;
    reg [63:0] _491;
    wire [7:0] _5198;
    wire _5199;
    wire [63:0] _5202;
    wire _5192;
    wire _5193;
    wire [63:0] _5194;
    wire _5189;
    wire _5190;
    wire [63:0] _5195;
    wire _5186;
    wire _5187;
    wire [63:0] _5197;
    wire [63:0] _5203;
    wire [63:0] _208;
    reg [63:0] _488;
    wire [7:0] _5217;
    wire _5218;
    wire [63:0] _5221;
    wire _5211;
    wire _5212;
    wire [63:0] _5213;
    wire _5208;
    wire _5209;
    wire [63:0] _5214;
    wire _5205;
    wire _5206;
    wire [63:0] _5216;
    wire [63:0] _5222;
    wire [63:0] _209;
    reg [63:0] _485;
    wire [7:0] _5236;
    wire _5237;
    wire [63:0] _5240;
    wire _5230;
    wire _5231;
    wire [63:0] _5232;
    wire _5227;
    wire _5228;
    wire [63:0] _5233;
    wire _5224;
    wire _5225;
    wire [63:0] _5235;
    wire [63:0] _5241;
    wire [63:0] _210;
    reg [63:0] _482;
    wire [7:0] _5255;
    wire _5256;
    wire [63:0] _5259;
    wire _5249;
    wire _5250;
    wire [63:0] _5251;
    wire _5246;
    wire _5247;
    wire [63:0] _5252;
    wire _5243;
    wire _5244;
    wire [63:0] _5254;
    wire [63:0] _5260;
    wire [63:0] _211;
    reg [63:0] _479;
    wire [7:0] _5274;
    wire _5275;
    wire [63:0] _5278;
    wire _5268;
    wire _5269;
    wire [63:0] _5270;
    wire _5265;
    wire _5266;
    wire [63:0] _5271;
    wire _5262;
    wire _5263;
    wire [63:0] _5273;
    wire [63:0] _5279;
    wire [63:0] _212;
    reg [63:0] _476;
    wire [7:0] _5293;
    wire _5294;
    wire [63:0] _5297;
    wire _5287;
    wire _5288;
    wire [63:0] _5289;
    wire _5284;
    wire _5285;
    wire [63:0] _5290;
    wire _5281;
    wire _5282;
    wire [63:0] _5292;
    wire [63:0] _5298;
    wire [63:0] _213;
    reg [63:0] _473;
    wire [7:0] _5312;
    wire _5313;
    wire [63:0] _5316;
    wire _5306;
    wire _5307;
    wire [63:0] _5308;
    wire _5303;
    wire _5304;
    wire [63:0] _5309;
    wire _5300;
    wire _5301;
    wire [63:0] _5311;
    wire [63:0] _5317;
    wire [63:0] _214;
    reg [63:0] _470;
    wire [7:0] _5331;
    wire _5332;
    wire [63:0] _5335;
    wire _5325;
    wire _5326;
    wire [63:0] _5327;
    wire _5322;
    wire _5323;
    wire [63:0] _5328;
    wire _5319;
    wire _5320;
    wire [63:0] _5330;
    wire [63:0] _5336;
    wire [63:0] _215;
    reg [63:0] _467;
    wire [7:0] _5350;
    wire _5351;
    wire [63:0] _5354;
    wire _5344;
    wire _5345;
    wire [63:0] _5346;
    wire _5341;
    wire _5342;
    wire [63:0] _5347;
    wire _5338;
    wire _5339;
    wire [63:0] _5349;
    wire [63:0] _5355;
    wire [63:0] _216;
    reg [63:0] _464;
    wire [7:0] _5369;
    wire _5370;
    wire [63:0] _5373;
    wire _5363;
    wire _5364;
    wire [63:0] _5365;
    wire _5360;
    wire _5361;
    wire [63:0] _5366;
    wire _5357;
    wire _5358;
    wire [63:0] _5368;
    wire [63:0] _5374;
    wire [63:0] _217;
    reg [63:0] _461;
    wire [7:0] _5388;
    wire _5389;
    wire [63:0] _5392;
    wire _5382;
    wire _5383;
    wire [63:0] _5384;
    wire _5379;
    wire _5380;
    wire [63:0] _5385;
    wire _5376;
    wire _5377;
    wire [63:0] _5387;
    wire [63:0] _5393;
    wire [63:0] _218;
    reg [63:0] _458;
    wire [7:0] _5407;
    wire _5408;
    wire [63:0] _5411;
    wire _5401;
    wire _5402;
    wire [63:0] _5403;
    wire _5398;
    wire _5399;
    wire [63:0] _5404;
    wire _5395;
    wire _5396;
    wire [63:0] _5406;
    wire [63:0] _5412;
    wire [63:0] _219;
    reg [63:0] _455;
    wire [7:0] _5426;
    wire _5427;
    wire [63:0] _5430;
    wire _5420;
    wire _5421;
    wire [63:0] _5422;
    wire _5417;
    wire _5418;
    wire [63:0] _5423;
    wire _5414;
    wire _5415;
    wire [63:0] _5425;
    wire [63:0] _5431;
    wire [63:0] _220;
    reg [63:0] _452;
    wire [7:0] _5445;
    wire _5446;
    wire [63:0] _5449;
    wire _5439;
    wire _5440;
    wire [63:0] _5441;
    wire _5436;
    wire _5437;
    wire [63:0] _5442;
    wire _5433;
    wire _5434;
    wire [63:0] _5444;
    wire [63:0] _5450;
    wire [63:0] _221;
    reg [63:0] _449;
    wire [7:0] _5464;
    wire _5465;
    wire [63:0] _5468;
    wire _5458;
    wire _5459;
    wire [63:0] _5460;
    wire _5455;
    wire _5456;
    wire [63:0] _5461;
    wire _5452;
    wire _5453;
    wire [63:0] _5463;
    wire [63:0] _5469;
    wire [63:0] _222;
    reg [63:0] _446;
    wire [7:0] _5483;
    wire _5484;
    wire [63:0] _5487;
    wire _5477;
    wire _5478;
    wire [63:0] _5479;
    wire _5474;
    wire _5475;
    wire [63:0] _5480;
    wire _5471;
    wire _5472;
    wire [63:0] _5482;
    wire [63:0] _5488;
    wire [63:0] _223;
    reg [63:0] _443;
    wire [7:0] _5502;
    wire _5503;
    wire [63:0] _5506;
    wire _5496;
    wire _5497;
    wire [63:0] _5498;
    wire _5493;
    wire _5494;
    wire [63:0] _5499;
    wire _5490;
    wire _5491;
    wire [63:0] _5501;
    wire [63:0] _5507;
    wire [63:0] _224;
    reg [63:0] _440;
    wire [7:0] _5521;
    wire _5522;
    wire [63:0] _5525;
    wire _5515;
    wire _5516;
    wire [63:0] _5517;
    wire _5512;
    wire _5513;
    wire [63:0] _5518;
    wire _5509;
    wire _5510;
    wire [63:0] _5520;
    wire [63:0] _5526;
    wire [63:0] _225;
    reg [63:0] _437;
    wire [7:0] _5540;
    wire _5541;
    wire [63:0] _5544;
    wire _5534;
    wire _5535;
    wire [63:0] _5536;
    wire _5531;
    wire _5532;
    wire [63:0] _5537;
    wire _5528;
    wire _5529;
    wire [63:0] _5539;
    wire [63:0] _5545;
    wire [63:0] _226;
    reg [63:0] _434;
    wire [7:0] _5559;
    wire _5560;
    wire [63:0] _5563;
    wire _5553;
    wire _5554;
    wire [63:0] _5555;
    wire _5550;
    wire _5551;
    wire [63:0] _5556;
    wire _5547;
    wire _5548;
    wire [63:0] _5558;
    wire [63:0] _5564;
    wire [63:0] _227;
    reg [63:0] _431;
    wire [7:0] _5578;
    wire _5579;
    wire [63:0] _5582;
    wire _5572;
    wire _5573;
    wire [63:0] _5574;
    wire _5569;
    wire _5570;
    wire [63:0] _5575;
    wire _5566;
    wire _5567;
    wire [63:0] _5577;
    wire [63:0] _5583;
    wire [63:0] _228;
    reg [63:0] _428;
    wire [7:0] _5597;
    wire _5598;
    wire [63:0] _5601;
    wire _5591;
    wire _5592;
    wire [63:0] _5593;
    wire _5588;
    wire _5589;
    wire [63:0] _5594;
    wire _5585;
    wire _5586;
    wire [63:0] _5596;
    wire [63:0] _5602;
    wire [63:0] _229;
    reg [63:0] _425;
    wire [7:0] _5616;
    wire _5617;
    wire [63:0] _5620;
    wire _5610;
    wire _5611;
    wire [63:0] _5612;
    wire _5607;
    wire _5608;
    wire [63:0] _5613;
    wire _5604;
    wire _5605;
    wire [63:0] _5615;
    wire [63:0] _5621;
    wire [63:0] _230;
    reg [63:0] _422;
    wire [7:0] _5635;
    wire _5636;
    wire [63:0] _5639;
    wire _5629;
    wire _5630;
    wire [63:0] _5631;
    wire _5626;
    wire _5627;
    wire [63:0] _5632;
    wire _5623;
    wire _5624;
    wire [63:0] _5634;
    wire [63:0] _5640;
    wire [63:0] _231;
    reg [63:0] _419;
    wire [7:0] _5654;
    wire _5655;
    wire [63:0] _5658;
    wire _5648;
    wire _5649;
    wire [63:0] _5650;
    wire _5645;
    wire _5646;
    wire [63:0] _5651;
    wire _5642;
    wire _5643;
    wire [63:0] _5653;
    wire [63:0] _5659;
    wire [63:0] _232;
    reg [63:0] _416;
    wire [7:0] _5673;
    wire _5674;
    wire [63:0] _5677;
    wire _5667;
    wire _5668;
    wire [63:0] _5669;
    wire _5664;
    wire _5665;
    wire [63:0] _5670;
    wire _5661;
    wire _5662;
    wire [63:0] _5672;
    wire [63:0] _5678;
    wire [63:0] _233;
    reg [63:0] _413;
    wire [7:0] _5692;
    wire _5693;
    wire [63:0] _5696;
    wire _5686;
    wire _5687;
    wire [63:0] _5688;
    wire _5683;
    wire _5684;
    wire [63:0] _5689;
    wire _5680;
    wire _5681;
    wire [63:0] _5691;
    wire [63:0] _5697;
    wire [63:0] _234;
    reg [63:0] _410;
    wire [7:0] _5711;
    wire _5712;
    wire [63:0] _5715;
    wire _5705;
    wire _5706;
    wire [63:0] _5707;
    wire _5702;
    wire _5703;
    wire [63:0] _5708;
    wire _5699;
    wire _5700;
    wire [63:0] _5710;
    wire [63:0] _5716;
    wire [63:0] _235;
    reg [63:0] _407;
    wire [7:0] _5730;
    wire _5731;
    wire [63:0] _5734;
    wire _5724;
    wire _5725;
    wire [63:0] _5726;
    wire _5721;
    wire _5722;
    wire [63:0] _5727;
    wire _5718;
    wire _5719;
    wire [63:0] _5729;
    wire [63:0] _5735;
    wire [63:0] _236;
    reg [63:0] _404;
    wire [7:0] _5749;
    wire _5750;
    wire [63:0] _5753;
    wire _5743;
    wire _5744;
    wire [63:0] _5745;
    wire _5740;
    wire _5741;
    wire [63:0] _5746;
    wire _5737;
    wire _5738;
    wire [63:0] _5748;
    wire [63:0] _5754;
    wire [63:0] _237;
    reg [63:0] _401;
    wire [7:0] _5768;
    wire _5769;
    wire [63:0] _5772;
    wire _5762;
    wire _5763;
    wire [63:0] _5764;
    wire _5759;
    wire _5760;
    wire [63:0] _5765;
    wire _5756;
    wire _5757;
    wire [63:0] _5767;
    wire [63:0] _5773;
    wire [63:0] _238;
    reg [63:0] _398;
    wire [7:0] _5787;
    wire _5788;
    wire [63:0] _5791;
    wire _5781;
    wire _5782;
    wire [63:0] _5783;
    wire _5778;
    wire _5779;
    wire [63:0] _5784;
    wire _5775;
    wire _5776;
    wire [63:0] _5786;
    wire [63:0] _5792;
    wire [63:0] _239;
    reg [63:0] _395;
    wire [7:0] _5806;
    wire _5807;
    wire [63:0] _5810;
    wire _5800;
    wire _5801;
    wire [63:0] _5802;
    wire _5797;
    wire _5798;
    wire [63:0] _5803;
    wire _5794;
    wire _5795;
    wire [63:0] _5805;
    wire [63:0] _5811;
    wire [63:0] _240;
    reg [63:0] _392;
    wire [7:0] _5825;
    wire _5826;
    wire [63:0] _5829;
    wire _5819;
    wire _5820;
    wire [63:0] _5821;
    wire _5816;
    wire _5817;
    wire [63:0] _5822;
    wire _5813;
    wire _5814;
    wire [63:0] _5824;
    wire [63:0] _5830;
    wire [63:0] _241;
    reg [63:0] _389;
    wire [7:0] _5844;
    wire _5845;
    wire [63:0] _5848;
    wire _5838;
    wire _5839;
    wire [63:0] _5840;
    wire _5835;
    wire _5836;
    wire [63:0] _5841;
    wire _5832;
    wire _5833;
    wire [63:0] _5843;
    wire [63:0] _5849;
    wire [63:0] _242;
    reg [63:0] _386;
    wire [7:0] _5863;
    wire _5864;
    wire [63:0] _5867;
    wire _5857;
    wire _5858;
    wire [63:0] _5859;
    wire _5854;
    wire _5855;
    wire [63:0] _5860;
    wire _5851;
    wire _5852;
    wire [63:0] _5862;
    wire [63:0] _5868;
    wire [63:0] _243;
    reg [63:0] _383;
    wire [7:0] _5882;
    wire _5883;
    wire [63:0] _5886;
    wire _5876;
    wire _5877;
    wire [63:0] _5878;
    wire _5873;
    wire _5874;
    wire [63:0] _5879;
    wire _5870;
    wire _5871;
    wire [63:0] _5881;
    wire [63:0] _5887;
    wire [63:0] _244;
    reg [63:0] _380;
    wire [7:0] _5901;
    wire _5902;
    wire [63:0] _5905;
    wire _5895;
    wire _5896;
    wire [63:0] _5897;
    wire _5892;
    wire _5893;
    wire [63:0] _5898;
    wire _5889;
    wire _5890;
    wire [63:0] _5900;
    wire [63:0] _5906;
    wire [63:0] _245;
    reg [63:0] _377;
    wire [7:0] _5920;
    wire _5921;
    wire [63:0] _5924;
    wire _5914;
    wire _5915;
    wire [63:0] _5916;
    wire _5911;
    wire _5912;
    wire [63:0] _5917;
    wire _5908;
    wire _5909;
    wire [63:0] _5919;
    wire [63:0] _5925;
    wire [63:0] _246;
    reg [63:0] _374;
    wire [7:0] _5939;
    wire _5940;
    wire [63:0] _5943;
    wire _5933;
    wire _5934;
    wire [63:0] _5935;
    wire _5930;
    wire _5931;
    wire [63:0] _5936;
    wire _5927;
    wire _5928;
    wire [63:0] _5938;
    wire [63:0] _5944;
    wire [63:0] _247;
    reg [63:0] _371;
    wire [7:0] _5958;
    wire _5959;
    wire [63:0] _5962;
    wire _5952;
    wire _5953;
    wire [63:0] _5954;
    wire _5949;
    wire _5950;
    wire [63:0] _5955;
    wire _5946;
    wire _5947;
    wire [63:0] _5957;
    wire [63:0] _5963;
    wire [63:0] _248;
    reg [63:0] _368;
    wire [7:0] _5977;
    wire _5978;
    wire [63:0] _5981;
    wire _5971;
    wire _5972;
    wire [63:0] _5973;
    wire _5968;
    wire _5969;
    wire [63:0] _5974;
    wire _5965;
    wire _5966;
    wire [63:0] _5976;
    wire [63:0] _5982;
    wire [63:0] _249;
    reg [63:0] _365;
    wire [7:0] _5996;
    wire _5997;
    wire [63:0] _6000;
    wire _5990;
    wire _5991;
    wire [63:0] _5992;
    wire _5987;
    wire _5988;
    wire [63:0] _5993;
    wire _5984;
    wire _5985;
    wire [63:0] _5995;
    wire [63:0] _6001;
    wire [63:0] _250;
    reg [63:0] _362;
    wire [7:0] _6015;
    wire _6016;
    wire [63:0] _6019;
    wire _6009;
    wire _6010;
    wire [63:0] _6011;
    wire _6006;
    wire _6007;
    wire [63:0] _6012;
    wire _6003;
    wire _6004;
    wire [63:0] _6014;
    wire [63:0] _6020;
    wire [63:0] _251;
    reg [63:0] _359;
    wire [7:0] _6034;
    wire _6035;
    wire [63:0] _6038;
    wire _6028;
    wire _6029;
    wire [63:0] _6030;
    wire _6025;
    wire _6026;
    wire [63:0] _6031;
    wire _6022;
    wire _6023;
    wire [63:0] _6033;
    wire [63:0] _6039;
    wire [63:0] _252;
    reg [63:0] _356;
    wire [7:0] _6053;
    wire _6054;
    wire [63:0] _6057;
    wire _6047;
    wire _6048;
    wire [63:0] _6049;
    wire _6044;
    wire _6045;
    wire [63:0] _6050;
    wire _6041;
    wire _6042;
    wire [63:0] _6052;
    wire [63:0] _6058;
    wire [63:0] _253;
    reg [63:0] _353;
    wire [7:0] _6072;
    wire _6073;
    wire [63:0] _6076;
    wire _6066;
    wire _6067;
    wire [63:0] _6068;
    wire _6063;
    wire _6064;
    wire [63:0] _6069;
    wire _6060;
    wire _6061;
    wire [63:0] _6071;
    wire [63:0] _6077;
    wire [63:0] _254;
    reg [63:0] _350;
    wire [7:0] _6091;
    wire _6092;
    wire [63:0] _6095;
    wire _6085;
    wire _6086;
    wire [63:0] _6087;
    wire _6082;
    wire _6083;
    wire [63:0] _6088;
    wire _6079;
    wire _6080;
    wire [63:0] _6090;
    wire [63:0] _6096;
    wire [63:0] _255;
    reg [63:0] _347;
    wire [7:0] _6110;
    wire _6111;
    wire [63:0] _6114;
    wire _6104;
    wire _6105;
    wire [63:0] _6106;
    wire _6101;
    wire _6102;
    wire [63:0] _6107;
    wire _6098;
    wire _6099;
    wire [63:0] _6109;
    wire [63:0] _6115;
    wire [63:0] _256;
    reg [63:0] _344;
    wire [7:0] _6129;
    wire _6130;
    wire [63:0] _6133;
    wire _6123;
    wire _6124;
    wire [63:0] _6125;
    wire _6120;
    wire _6121;
    wire [63:0] _6126;
    wire _6117;
    wire _6118;
    wire [63:0] _6128;
    wire [63:0] _6134;
    wire [63:0] _257;
    reg [63:0] _341;
    wire [7:0] _6148;
    wire _6149;
    wire [63:0] _6152;
    wire _6142;
    wire _6143;
    wire [63:0] _6144;
    wire _6139;
    wire _6140;
    wire [63:0] _6145;
    wire _6136;
    wire _6137;
    wire [63:0] _6147;
    wire [63:0] _6153;
    wire [63:0] _258;
    reg [63:0] _338;
    wire [7:0] _6167;
    wire _6168;
    wire [63:0] _6171;
    wire _6161;
    wire _6162;
    wire [63:0] _6163;
    wire _6158;
    wire _6159;
    wire [63:0] _6164;
    wire _6155;
    wire _6156;
    wire [63:0] _6166;
    wire [63:0] _6172;
    wire [63:0] _259;
    reg [63:0] _335;
    wire [7:0] _6186;
    wire _6187;
    wire [63:0] _6190;
    wire _6180;
    wire _6181;
    wire [63:0] _6182;
    wire _6177;
    wire _6178;
    wire [63:0] _6183;
    wire _6174;
    wire _6175;
    wire [63:0] _6185;
    wire [63:0] _6191;
    wire [63:0] _260;
    reg [63:0] _332;
    wire [7:0] _6205;
    wire _6206;
    wire [63:0] _6209;
    wire _6199;
    wire _6200;
    wire [63:0] _6201;
    wire _6196;
    wire _6197;
    wire [63:0] _6202;
    wire _6193;
    wire _6194;
    wire [63:0] _6204;
    wire [63:0] _6210;
    wire [63:0] _261;
    reg [63:0] _329;
    reg [63:0] _1393;
    wire [63:0] _1394;
    wire _6218;
    wire _6219;
    wire [63:0] _6220;
    wire _6215;
    wire _6216;
    wire [63:0] _6221;
    wire _6212;
    wire _6213;
    wire [63:0] _6223;
    wire [63:0] _6229;
    wire [63:0] _262;
    reg [63:0] _326;
    reg [63:0] _1390;
    wire [63:0] _1391;
    wire [7:0] _1386;
    wire _6237;
    wire _6238;
    wire [63:0] _6239;
    wire [7:0] _1381;
    wire _6234;
    wire _6235;
    wire [63:0] _6240;
    wire _6231;
    wire _6232;
    wire [63:0] _6242;
    wire [63:0] _6248;
    wire [63:0] _263;
    reg [63:0] _323;
    reg [63:0] _1114;
    wire _1116;
    wire _1117;
    wire _1113;
    wire _1118;
    wire _1376;
    wire [63:0] _6254;
    wire [63:0] _6256;
    wire [63:0] _264;
    reg [63:0] _6251;
    wire _6258;
    wire [2:0] _289;
    wire [2:0] _1104;
    wire [2:0] _6298;
    wire [2:0] _6257;
    wire [7:0] _6259;
    wire [7:0] _267;
    reg [7:0] _315;
    wire [7:0] _6264;
    wire [7:0] _6265;
    wire _305;
    wire _269;
    wire _6260;
    wire _6262;
    wire _270;
    reg _306;
    wire _307;
    wire [7:0] _6267;
    wire [7:0] _6269;
    wire [7:0] _271;
    reg [7:0] _312;
    wire _316;
    wire _1096;
    wire [2:0] _308;
    wire _309;
    wire _1097;
    wire [2:0] _6297;
    wire [7:0] _6280;
    wire [7:0] _6272;
    wire _6270;
    wire [7:0] _6273;
    wire [7:0] _6281;
    wire [7:0] _6283;
    wire [7:0] _272;
    reg [7:0] _299;
    wire [7:0] _6285;
    wire [7:0] _6286;
    wire [7:0] _6288;
    wire [7:0] _273;
    reg [7:0] _6279;
    wire vdd;
    wire _275;
    wire _277;
    wire [7:0] _279;
    wire [6:0] _6290;
    wire [7:0] _6291;
    wire [7:0] _6292;
    wire [7:0] _280;
    reg [7:0] _6276;
    wire [7:0] _6293;
    wire [7:0] _6294;
    wire [7:0] _6296;
    wire [7:0] _281;
    reg [7:0] _296;
    wire _300;
    wire _301;
    wire _302;
    wire [2:0] _292;
    wire _293;
    wire _303;
    wire [2:0] _6299;
    wire _283;
    wire _1106;
    wire [2:0] _6300;
    wire _285;
    wire [2:0] _6301;
    wire [2:0] _286;
    reg [2:0] _291;
    wire _1105;
    assign _1099 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    always @* begin
        case (_312)
        0:
            _1089 <= _323;
        1:
            _1089 <= _326;
        2:
            _1089 <= _329;
        3:
            _1089 <= _332;
        4:
            _1089 <= _335;
        5:
            _1089 <= _338;
        6:
            _1089 <= _341;
        7:
            _1089 <= _344;
        8:
            _1089 <= _347;
        9:
            _1089 <= _350;
        10:
            _1089 <= _353;
        11:
            _1089 <= _356;
        12:
            _1089 <= _359;
        13:
            _1089 <= _362;
        14:
            _1089 <= _365;
        15:
            _1089 <= _368;
        16:
            _1089 <= _371;
        17:
            _1089 <= _374;
        18:
            _1089 <= _377;
        19:
            _1089 <= _380;
        20:
            _1089 <= _383;
        21:
            _1089 <= _386;
        22:
            _1089 <= _389;
        23:
            _1089 <= _392;
        24:
            _1089 <= _395;
        25:
            _1089 <= _398;
        26:
            _1089 <= _401;
        27:
            _1089 <= _404;
        28:
            _1089 <= _407;
        29:
            _1089 <= _410;
        30:
            _1089 <= _413;
        31:
            _1089 <= _416;
        32:
            _1089 <= _419;
        33:
            _1089 <= _422;
        34:
            _1089 <= _425;
        35:
            _1089 <= _428;
        36:
            _1089 <= _431;
        37:
            _1089 <= _434;
        38:
            _1089 <= _437;
        39:
            _1089 <= _440;
        40:
            _1089 <= _443;
        41:
            _1089 <= _446;
        42:
            _1089 <= _449;
        43:
            _1089 <= _452;
        44:
            _1089 <= _455;
        45:
            _1089 <= _458;
        46:
            _1089 <= _461;
        47:
            _1089 <= _464;
        48:
            _1089 <= _467;
        49:
            _1089 <= _470;
        50:
            _1089 <= _473;
        51:
            _1089 <= _476;
        52:
            _1089 <= _479;
        53:
            _1089 <= _482;
        54:
            _1089 <= _485;
        55:
            _1089 <= _488;
        56:
            _1089 <= _491;
        57:
            _1089 <= _494;
        58:
            _1089 <= _497;
        59:
            _1089 <= _500;
        60:
            _1089 <= _503;
        61:
            _1089 <= _506;
        62:
            _1089 <= _509;
        63:
            _1089 <= _512;
        64:
            _1089 <= _515;
        65:
            _1089 <= _518;
        66:
            _1089 <= _521;
        67:
            _1089 <= _524;
        68:
            _1089 <= _527;
        69:
            _1089 <= _530;
        70:
            _1089 <= _533;
        71:
            _1089 <= _536;
        72:
            _1089 <= _539;
        73:
            _1089 <= _542;
        74:
            _1089 <= _545;
        75:
            _1089 <= _548;
        76:
            _1089 <= _551;
        77:
            _1089 <= _554;
        78:
            _1089 <= _557;
        79:
            _1089 <= _560;
        80:
            _1089 <= _563;
        81:
            _1089 <= _566;
        82:
            _1089 <= _569;
        83:
            _1089 <= _572;
        84:
            _1089 <= _575;
        85:
            _1089 <= _578;
        86:
            _1089 <= _581;
        87:
            _1089 <= _584;
        88:
            _1089 <= _587;
        89:
            _1089 <= _590;
        90:
            _1089 <= _593;
        91:
            _1089 <= _596;
        92:
            _1089 <= _599;
        93:
            _1089 <= _602;
        94:
            _1089 <= _605;
        95:
            _1089 <= _608;
        96:
            _1089 <= _611;
        97:
            _1089 <= _614;
        98:
            _1089 <= _617;
        99:
            _1089 <= _620;
        100:
            _1089 <= _623;
        101:
            _1089 <= _626;
        102:
            _1089 <= _629;
        103:
            _1089 <= _632;
        104:
            _1089 <= _635;
        105:
            _1089 <= _638;
        106:
            _1089 <= _641;
        107:
            _1089 <= _644;
        108:
            _1089 <= _647;
        109:
            _1089 <= _650;
        110:
            _1089 <= _653;
        111:
            _1089 <= _656;
        112:
            _1089 <= _659;
        113:
            _1089 <= _662;
        114:
            _1089 <= _665;
        115:
            _1089 <= _668;
        116:
            _1089 <= _671;
        117:
            _1089 <= _674;
        118:
            _1089 <= _677;
        119:
            _1089 <= _680;
        120:
            _1089 <= _683;
        121:
            _1089 <= _686;
        122:
            _1089 <= _689;
        123:
            _1089 <= _692;
        124:
            _1089 <= _695;
        125:
            _1089 <= _698;
        126:
            _1089 <= _701;
        127:
            _1089 <= _704;
        128:
            _1089 <= _707;
        129:
            _1089 <= _710;
        130:
            _1089 <= _713;
        131:
            _1089 <= _716;
        132:
            _1089 <= _719;
        133:
            _1089 <= _722;
        134:
            _1089 <= _725;
        135:
            _1089 <= _728;
        136:
            _1089 <= _731;
        137:
            _1089 <= _734;
        138:
            _1089 <= _737;
        139:
            _1089 <= _740;
        140:
            _1089 <= _743;
        141:
            _1089 <= _746;
        142:
            _1089 <= _749;
        143:
            _1089 <= _752;
        144:
            _1089 <= _755;
        145:
            _1089 <= _758;
        146:
            _1089 <= _761;
        147:
            _1089 <= _764;
        148:
            _1089 <= _767;
        149:
            _1089 <= _770;
        150:
            _1089 <= _773;
        151:
            _1089 <= _776;
        152:
            _1089 <= _779;
        153:
            _1089 <= _782;
        154:
            _1089 <= _785;
        155:
            _1089 <= _788;
        156:
            _1089 <= _791;
        157:
            _1089 <= _794;
        158:
            _1089 <= _797;
        159:
            _1089 <= _800;
        160:
            _1089 <= _803;
        161:
            _1089 <= _806;
        162:
            _1089 <= _809;
        163:
            _1089 <= _812;
        164:
            _1089 <= _815;
        165:
            _1089 <= _818;
        166:
            _1089 <= _821;
        167:
            _1089 <= _824;
        168:
            _1089 <= _827;
        169:
            _1089 <= _830;
        170:
            _1089 <= _833;
        171:
            _1089 <= _836;
        172:
            _1089 <= _839;
        173:
            _1089 <= _842;
        174:
            _1089 <= _845;
        175:
            _1089 <= _848;
        176:
            _1089 <= _851;
        177:
            _1089 <= _854;
        178:
            _1089 <= _857;
        179:
            _1089 <= _860;
        180:
            _1089 <= _863;
        181:
            _1089 <= _866;
        182:
            _1089 <= _869;
        183:
            _1089 <= _872;
        184:
            _1089 <= _875;
        185:
            _1089 <= _878;
        186:
            _1089 <= _881;
        187:
            _1089 <= _884;
        188:
            _1089 <= _887;
        189:
            _1089 <= _890;
        190:
            _1089 <= _893;
        191:
            _1089 <= _896;
        192:
            _1089 <= _899;
        193:
            _1089 <= _902;
        194:
            _1089 <= _905;
        195:
            _1089 <= _908;
        196:
            _1089 <= _911;
        197:
            _1089 <= _914;
        198:
            _1089 <= _917;
        199:
            _1089 <= _920;
        200:
            _1089 <= _923;
        201:
            _1089 <= _926;
        202:
            _1089 <= _929;
        203:
            _1089 <= _932;
        204:
            _1089 <= _935;
        205:
            _1089 <= _938;
        206:
            _1089 <= _941;
        207:
            _1089 <= _944;
        208:
            _1089 <= _947;
        209:
            _1089 <= _950;
        210:
            _1089 <= _953;
        211:
            _1089 <= _956;
        212:
            _1089 <= _959;
        213:
            _1089 <= _962;
        214:
            _1089 <= _965;
        215:
            _1089 <= _968;
        216:
            _1089 <= _971;
        217:
            _1089 <= _974;
        218:
            _1089 <= _977;
        219:
            _1089 <= _980;
        220:
            _1089 <= _983;
        221:
            _1089 <= _986;
        222:
            _1089 <= _989;
        223:
            _1089 <= _992;
        224:
            _1089 <= _995;
        225:
            _1089 <= _998;
        226:
            _1089 <= _1001;
        227:
            _1089 <= _1004;
        228:
            _1089 <= _1007;
        229:
            _1089 <= _1010;
        230:
            _1089 <= _1013;
        231:
            _1089 <= _1016;
        232:
            _1089 <= _1019;
        233:
            _1089 <= _1022;
        234:
            _1089 <= _1025;
        235:
            _1089 <= _1028;
        236:
            _1089 <= _1031;
        237:
            _1089 <= _1034;
        238:
            _1089 <= _1037;
        239:
            _1089 <= _1040;
        240:
            _1089 <= _1043;
        241:
            _1089 <= _1046;
        242:
            _1089 <= _1049;
        243:
            _1089 <= _1052;
        244:
            _1089 <= _1055;
        245:
            _1089 <= _1058;
        246:
            _1089 <= _1061;
        247:
            _1089 <= _1064;
        248:
            _1089 <= _1067;
        249:
            _1089 <= _1070;
        250:
            _1089 <= _1073;
        251:
            _1089 <= _1076;
        252:
            _1089 <= _1079;
        253:
            _1089 <= _1082;
        254:
            _1089 <= _1085;
        default:
            _1089 <= _1088;
        endcase
    end
    assign _1090 = _320 + _1089;
    assign _317 = _309 & _316;
    assign _1091 = _317 ? _1090 : _320;
    assign _1093 = _307 ? _1099 : _1091;
    assign _1095 = _285 ? _1099 : _1093;
    assign _2 = _1095;
    always @(posedge _277) begin
        if (_275)
            _320 <= _1099;
        else
            _320 <= _2;
    end
    assign _1101 = _1097 ? _320 : _1100;
    assign _1103 = _285 ? _1099 : _1101;
    assign _3 = _1103;
    always @(posedge _277) begin
        if (_275)
            _1100 <= _1099;
        else
            _1100 <= _3;
    end
    assign _6252 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    assign _6253 = _6251 + _6252;
    assign _1374 = _1109[255:255];
    assign _1373 = _1109[254:254];
    assign _1372 = _1109[253:253];
    assign _1371 = _1109[252:252];
    assign _1370 = _1109[251:251];
    assign _1369 = _1109[250:250];
    assign _1368 = _1109[249:249];
    assign _1367 = _1109[248:248];
    assign _1366 = _1109[247:247];
    assign _1365 = _1109[246:246];
    assign _1364 = _1109[245:245];
    assign _1363 = _1109[244:244];
    assign _1362 = _1109[243:243];
    assign _1361 = _1109[242:242];
    assign _1360 = _1109[241:241];
    assign _1359 = _1109[240:240];
    assign _1358 = _1109[239:239];
    assign _1357 = _1109[238:238];
    assign _1356 = _1109[237:237];
    assign _1355 = _1109[236:236];
    assign _1354 = _1109[235:235];
    assign _1353 = _1109[234:234];
    assign _1352 = _1109[233:233];
    assign _1351 = _1109[232:232];
    assign _1350 = _1109[231:231];
    assign _1349 = _1109[230:230];
    assign _1348 = _1109[229:229];
    assign _1347 = _1109[228:228];
    assign _1346 = _1109[227:227];
    assign _1345 = _1109[226:226];
    assign _1344 = _1109[225:225];
    assign _1343 = _1109[224:224];
    assign _1342 = _1109[223:223];
    assign _1341 = _1109[222:222];
    assign _1340 = _1109[221:221];
    assign _1339 = _1109[220:220];
    assign _1338 = _1109[219:219];
    assign _1337 = _1109[218:218];
    assign _1336 = _1109[217:217];
    assign _1335 = _1109[216:216];
    assign _1334 = _1109[215:215];
    assign _1333 = _1109[214:214];
    assign _1332 = _1109[213:213];
    assign _1331 = _1109[212:212];
    assign _1330 = _1109[211:211];
    assign _1329 = _1109[210:210];
    assign _1328 = _1109[209:209];
    assign _1327 = _1109[208:208];
    assign _1326 = _1109[207:207];
    assign _1325 = _1109[206:206];
    assign _1324 = _1109[205:205];
    assign _1323 = _1109[204:204];
    assign _1322 = _1109[203:203];
    assign _1321 = _1109[202:202];
    assign _1320 = _1109[201:201];
    assign _1319 = _1109[200:200];
    assign _1318 = _1109[199:199];
    assign _1317 = _1109[198:198];
    assign _1316 = _1109[197:197];
    assign _1315 = _1109[196:196];
    assign _1314 = _1109[195:195];
    assign _1313 = _1109[194:194];
    assign _1312 = _1109[193:193];
    assign _1311 = _1109[192:192];
    assign _1310 = _1109[191:191];
    assign _1309 = _1109[190:190];
    assign _1308 = _1109[189:189];
    assign _1307 = _1109[188:188];
    assign _1306 = _1109[187:187];
    assign _1305 = _1109[186:186];
    assign _1304 = _1109[185:185];
    assign _1303 = _1109[184:184];
    assign _1302 = _1109[183:183];
    assign _1301 = _1109[182:182];
    assign _1300 = _1109[181:181];
    assign _1299 = _1109[180:180];
    assign _1298 = _1109[179:179];
    assign _1297 = _1109[178:178];
    assign _1296 = _1109[177:177];
    assign _1295 = _1109[176:176];
    assign _1294 = _1109[175:175];
    assign _1293 = _1109[174:174];
    assign _1292 = _1109[173:173];
    assign _1291 = _1109[172:172];
    assign _1290 = _1109[171:171];
    assign _1289 = _1109[170:170];
    assign _1288 = _1109[169:169];
    assign _1287 = _1109[168:168];
    assign _1286 = _1109[167:167];
    assign _1285 = _1109[166:166];
    assign _1284 = _1109[165:165];
    assign _1283 = _1109[164:164];
    assign _1282 = _1109[163:163];
    assign _1281 = _1109[162:162];
    assign _1280 = _1109[161:161];
    assign _1279 = _1109[160:160];
    assign _1278 = _1109[159:159];
    assign _1277 = _1109[158:158];
    assign _1276 = _1109[157:157];
    assign _1275 = _1109[156:156];
    assign _1274 = _1109[155:155];
    assign _1273 = _1109[154:154];
    assign _1272 = _1109[153:153];
    assign _1271 = _1109[152:152];
    assign _1270 = _1109[151:151];
    assign _1269 = _1109[150:150];
    assign _1268 = _1109[149:149];
    assign _1267 = _1109[148:148];
    assign _1266 = _1109[147:147];
    assign _1265 = _1109[146:146];
    assign _1264 = _1109[145:145];
    assign _1263 = _1109[144:144];
    assign _1262 = _1109[143:143];
    assign _1261 = _1109[142:142];
    assign _1260 = _1109[141:141];
    assign _1259 = _1109[140:140];
    assign _1258 = _1109[139:139];
    assign _1257 = _1109[138:138];
    assign _1256 = _1109[137:137];
    assign _1255 = _1109[136:136];
    assign _1254 = _1109[135:135];
    assign _1253 = _1109[134:134];
    assign _1252 = _1109[133:133];
    assign _1251 = _1109[132:132];
    assign _1250 = _1109[131:131];
    assign _1249 = _1109[130:130];
    assign _1248 = _1109[129:129];
    assign _1247 = _1109[128:128];
    assign _1246 = _1109[127:127];
    assign _1245 = _1109[126:126];
    assign _1244 = _1109[125:125];
    assign _1243 = _1109[124:124];
    assign _1242 = _1109[123:123];
    assign _1241 = _1109[122:122];
    assign _1240 = _1109[121:121];
    assign _1239 = _1109[120:120];
    assign _1238 = _1109[119:119];
    assign _1237 = _1109[118:118];
    assign _1236 = _1109[117:117];
    assign _1235 = _1109[116:116];
    assign _1234 = _1109[115:115];
    assign _1233 = _1109[114:114];
    assign _1232 = _1109[113:113];
    assign _1231 = _1109[112:112];
    assign _1230 = _1109[111:111];
    assign _1229 = _1109[110:110];
    assign _1228 = _1109[109:109];
    assign _1227 = _1109[108:108];
    assign _1226 = _1109[107:107];
    assign _1225 = _1109[106:106];
    assign _1224 = _1109[105:105];
    assign _1223 = _1109[104:104];
    assign _1222 = _1109[103:103];
    assign _1221 = _1109[102:102];
    assign _1220 = _1109[101:101];
    assign _1219 = _1109[100:100];
    assign _1218 = _1109[99:99];
    assign _1217 = _1109[98:98];
    assign _1216 = _1109[97:97];
    assign _1215 = _1109[96:96];
    assign _1214 = _1109[95:95];
    assign _1213 = _1109[94:94];
    assign _1212 = _1109[93:93];
    assign _1211 = _1109[92:92];
    assign _1210 = _1109[91:91];
    assign _1209 = _1109[90:90];
    assign _1208 = _1109[89:89];
    assign _1207 = _1109[88:88];
    assign _1206 = _1109[87:87];
    assign _1205 = _1109[86:86];
    assign _1204 = _1109[85:85];
    assign _1203 = _1109[84:84];
    assign _1202 = _1109[83:83];
    assign _1201 = _1109[82:82];
    assign _1200 = _1109[81:81];
    assign _1199 = _1109[80:80];
    assign _1198 = _1109[79:79];
    assign _1197 = _1109[78:78];
    assign _1196 = _1109[77:77];
    assign _1195 = _1109[76:76];
    assign _1194 = _1109[75:75];
    assign _1193 = _1109[74:74];
    assign _1192 = _1109[73:73];
    assign _1191 = _1109[72:72];
    assign _1190 = _1109[71:71];
    assign _1189 = _1109[70:70];
    assign _1188 = _1109[69:69];
    assign _1187 = _1109[68:68];
    assign _1186 = _1109[67:67];
    assign _1185 = _1109[66:66];
    assign _1184 = _1109[65:65];
    assign _1183 = _1109[64:64];
    assign _1182 = _1109[63:63];
    assign _1181 = _1109[62:62];
    assign _1180 = _1109[61:61];
    assign _1179 = _1109[60:60];
    assign _1178 = _1109[59:59];
    assign _1177 = _1109[58:58];
    assign _1176 = _1109[57:57];
    assign _1175 = _1109[56:56];
    assign _1174 = _1109[55:55];
    assign _1173 = _1109[54:54];
    assign _1172 = _1109[53:53];
    assign _1171 = _1109[52:52];
    assign _1170 = _1109[51:51];
    assign _1169 = _1109[50:50];
    assign _1168 = _1109[49:49];
    assign _1167 = _1109[48:48];
    assign _1166 = _1109[47:47];
    assign _1165 = _1109[46:46];
    assign _1164 = _1109[45:45];
    assign _1163 = _1109[44:44];
    assign _1162 = _1109[43:43];
    assign _1161 = _1109[42:42];
    assign _1160 = _1109[41:41];
    assign _1159 = _1109[40:40];
    assign _1158 = _1109[39:39];
    assign _1157 = _1109[38:38];
    assign _1156 = _1109[37:37];
    assign _1155 = _1109[36:36];
    assign _1154 = _1109[35:35];
    assign _1153 = _1109[34:34];
    assign _1152 = _1109[33:33];
    assign _1151 = _1109[32:32];
    assign _1150 = _1109[31:31];
    assign _1149 = _1109[30:30];
    assign _1148 = _1109[29:29];
    assign _1147 = _1109[28:28];
    assign _1146 = _1109[27:27];
    assign _1145 = _1109[26:26];
    assign _1144 = _1109[25:25];
    assign _1143 = _1109[24:24];
    assign _1142 = _1109[23:23];
    assign _1141 = _1109[22:22];
    assign _1140 = _1109[21:21];
    assign _1139 = _1109[20:20];
    assign _1138 = _1109[19:19];
    assign _1137 = _1109[18:18];
    assign _1136 = _1109[17:17];
    assign _1135 = _1109[16:16];
    assign _1134 = _1109[15:15];
    assign _1133 = _1109[14:14];
    assign _1132 = _1109[13:13];
    assign _1131 = _1109[12:12];
    assign _1130 = _1109[11:11];
    assign _1129 = _1109[10:10];
    assign _1128 = _1109[9:9];
    assign _1127 = _1109[8:8];
    assign _1126 = _1109[7:7];
    assign _1125 = _1109[6:6];
    assign _1124 = _1109[5:5];
    assign _1123 = _1109[4:4];
    assign _1122 = _1109[3:3];
    assign _1121 = _1109[2:2];
    assign _1120 = _1109[1:1];
    assign _1108 = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign _6 = row_bits;
    assign _1110 = _1106 ? _6 : _1109;
    assign _1112 = _285 ? _1108 : _1110;
    assign _7 = _1112;
    always @(posedge _277) begin
        if (_275)
            _1109 <= _1108;
        else
            _1109 <= _7;
    end
    assign _1119 = _1109[0:0];
    always @* begin
        case (_299)
        0:
            _1375 <= _1119;
        1:
            _1375 <= _1120;
        2:
            _1375 <= _1121;
        3:
            _1375 <= _1122;
        4:
            _1375 <= _1123;
        5:
            _1375 <= _1124;
        6:
            _1375 <= _1125;
        7:
            _1375 <= _1126;
        8:
            _1375 <= _1127;
        9:
            _1375 <= _1128;
        10:
            _1375 <= _1129;
        11:
            _1375 <= _1130;
        12:
            _1375 <= _1131;
        13:
            _1375 <= _1132;
        14:
            _1375 <= _1133;
        15:
            _1375 <= _1134;
        16:
            _1375 <= _1135;
        17:
            _1375 <= _1136;
        18:
            _1375 <= _1137;
        19:
            _1375 <= _1138;
        20:
            _1375 <= _1139;
        21:
            _1375 <= _1140;
        22:
            _1375 <= _1141;
        23:
            _1375 <= _1142;
        24:
            _1375 <= _1143;
        25:
            _1375 <= _1144;
        26:
            _1375 <= _1145;
        27:
            _1375 <= _1146;
        28:
            _1375 <= _1147;
        29:
            _1375 <= _1148;
        30:
            _1375 <= _1149;
        31:
            _1375 <= _1150;
        32:
            _1375 <= _1151;
        33:
            _1375 <= _1152;
        34:
            _1375 <= _1153;
        35:
            _1375 <= _1154;
        36:
            _1375 <= _1155;
        37:
            _1375 <= _1156;
        38:
            _1375 <= _1157;
        39:
            _1375 <= _1158;
        40:
            _1375 <= _1159;
        41:
            _1375 <= _1160;
        42:
            _1375 <= _1161;
        43:
            _1375 <= _1162;
        44:
            _1375 <= _1163;
        45:
            _1375 <= _1164;
        46:
            _1375 <= _1165;
        47:
            _1375 <= _1166;
        48:
            _1375 <= _1167;
        49:
            _1375 <= _1168;
        50:
            _1375 <= _1169;
        51:
            _1375 <= _1170;
        52:
            _1375 <= _1171;
        53:
            _1375 <= _1172;
        54:
            _1375 <= _1173;
        55:
            _1375 <= _1174;
        56:
            _1375 <= _1175;
        57:
            _1375 <= _1176;
        58:
            _1375 <= _1177;
        59:
            _1375 <= _1178;
        60:
            _1375 <= _1179;
        61:
            _1375 <= _1180;
        62:
            _1375 <= _1181;
        63:
            _1375 <= _1182;
        64:
            _1375 <= _1183;
        65:
            _1375 <= _1184;
        66:
            _1375 <= _1185;
        67:
            _1375 <= _1186;
        68:
            _1375 <= _1187;
        69:
            _1375 <= _1188;
        70:
            _1375 <= _1189;
        71:
            _1375 <= _1190;
        72:
            _1375 <= _1191;
        73:
            _1375 <= _1192;
        74:
            _1375 <= _1193;
        75:
            _1375 <= _1194;
        76:
            _1375 <= _1195;
        77:
            _1375 <= _1196;
        78:
            _1375 <= _1197;
        79:
            _1375 <= _1198;
        80:
            _1375 <= _1199;
        81:
            _1375 <= _1200;
        82:
            _1375 <= _1201;
        83:
            _1375 <= _1202;
        84:
            _1375 <= _1203;
        85:
            _1375 <= _1204;
        86:
            _1375 <= _1205;
        87:
            _1375 <= _1206;
        88:
            _1375 <= _1207;
        89:
            _1375 <= _1208;
        90:
            _1375 <= _1209;
        91:
            _1375 <= _1210;
        92:
            _1375 <= _1211;
        93:
            _1375 <= _1212;
        94:
            _1375 <= _1213;
        95:
            _1375 <= _1214;
        96:
            _1375 <= _1215;
        97:
            _1375 <= _1216;
        98:
            _1375 <= _1217;
        99:
            _1375 <= _1218;
        100:
            _1375 <= _1219;
        101:
            _1375 <= _1220;
        102:
            _1375 <= _1221;
        103:
            _1375 <= _1222;
        104:
            _1375 <= _1223;
        105:
            _1375 <= _1224;
        106:
            _1375 <= _1225;
        107:
            _1375 <= _1226;
        108:
            _1375 <= _1227;
        109:
            _1375 <= _1228;
        110:
            _1375 <= _1229;
        111:
            _1375 <= _1230;
        112:
            _1375 <= _1231;
        113:
            _1375 <= _1232;
        114:
            _1375 <= _1233;
        115:
            _1375 <= _1234;
        116:
            _1375 <= _1235;
        117:
            _1375 <= _1236;
        118:
            _1375 <= _1237;
        119:
            _1375 <= _1238;
        120:
            _1375 <= _1239;
        121:
            _1375 <= _1240;
        122:
            _1375 <= _1241;
        123:
            _1375 <= _1242;
        124:
            _1375 <= _1243;
        125:
            _1375 <= _1244;
        126:
            _1375 <= _1245;
        127:
            _1375 <= _1246;
        128:
            _1375 <= _1247;
        129:
            _1375 <= _1248;
        130:
            _1375 <= _1249;
        131:
            _1375 <= _1250;
        132:
            _1375 <= _1251;
        133:
            _1375 <= _1252;
        134:
            _1375 <= _1253;
        135:
            _1375 <= _1254;
        136:
            _1375 <= _1255;
        137:
            _1375 <= _1256;
        138:
            _1375 <= _1257;
        139:
            _1375 <= _1258;
        140:
            _1375 <= _1259;
        141:
            _1375 <= _1260;
        142:
            _1375 <= _1261;
        143:
            _1375 <= _1262;
        144:
            _1375 <= _1263;
        145:
            _1375 <= _1264;
        146:
            _1375 <= _1265;
        147:
            _1375 <= _1266;
        148:
            _1375 <= _1267;
        149:
            _1375 <= _1268;
        150:
            _1375 <= _1269;
        151:
            _1375 <= _1270;
        152:
            _1375 <= _1271;
        153:
            _1375 <= _1272;
        154:
            _1375 <= _1273;
        155:
            _1375 <= _1274;
        156:
            _1375 <= _1275;
        157:
            _1375 <= _1276;
        158:
            _1375 <= _1277;
        159:
            _1375 <= _1278;
        160:
            _1375 <= _1279;
        161:
            _1375 <= _1280;
        162:
            _1375 <= _1281;
        163:
            _1375 <= _1282;
        164:
            _1375 <= _1283;
        165:
            _1375 <= _1284;
        166:
            _1375 <= _1285;
        167:
            _1375 <= _1286;
        168:
            _1375 <= _1287;
        169:
            _1375 <= _1288;
        170:
            _1375 <= _1289;
        171:
            _1375 <= _1290;
        172:
            _1375 <= _1291;
        173:
            _1375 <= _1292;
        174:
            _1375 <= _1293;
        175:
            _1375 <= _1294;
        176:
            _1375 <= _1295;
        177:
            _1375 <= _1296;
        178:
            _1375 <= _1297;
        179:
            _1375 <= _1298;
        180:
            _1375 <= _1299;
        181:
            _1375 <= _1300;
        182:
            _1375 <= _1301;
        183:
            _1375 <= _1302;
        184:
            _1375 <= _1303;
        185:
            _1375 <= _1304;
        186:
            _1375 <= _1305;
        187:
            _1375 <= _1306;
        188:
            _1375 <= _1307;
        189:
            _1375 <= _1308;
        190:
            _1375 <= _1309;
        191:
            _1375 <= _1310;
        192:
            _1375 <= _1311;
        193:
            _1375 <= _1312;
        194:
            _1375 <= _1313;
        195:
            _1375 <= _1314;
        196:
            _1375 <= _1315;
        197:
            _1375 <= _1316;
        198:
            _1375 <= _1317;
        199:
            _1375 <= _1318;
        200:
            _1375 <= _1319;
        201:
            _1375 <= _1320;
        202:
            _1375 <= _1321;
        203:
            _1375 <= _1322;
        204:
            _1375 <= _1323;
        205:
            _1375 <= _1324;
        206:
            _1375 <= _1325;
        207:
            _1375 <= _1326;
        208:
            _1375 <= _1327;
        209:
            _1375 <= _1328;
        210:
            _1375 <= _1329;
        211:
            _1375 <= _1330;
        212:
            _1375 <= _1331;
        213:
            _1375 <= _1332;
        214:
            _1375 <= _1333;
        215:
            _1375 <= _1334;
        216:
            _1375 <= _1335;
        217:
            _1375 <= _1336;
        218:
            _1375 <= _1337;
        219:
            _1375 <= _1338;
        220:
            _1375 <= _1339;
        221:
            _1375 <= _1340;
        222:
            _1375 <= _1341;
        223:
            _1375 <= _1342;
        224:
            _1375 <= _1343;
        225:
            _1375 <= _1344;
        226:
            _1375 <= _1345;
        227:
            _1375 <= _1346;
        228:
            _1375 <= _1347;
        229:
            _1375 <= _1348;
        230:
            _1375 <= _1349;
        231:
            _1375 <= _1350;
        232:
            _1375 <= _1351;
        233:
            _1375 <= _1352;
        234:
            _1375 <= _1353;
        235:
            _1375 <= _1354;
        236:
            _1375 <= _1355;
        237:
            _1375 <= _1356;
        238:
            _1375 <= _1357;
        239:
            _1375 <= _1358;
        240:
            _1375 <= _1359;
        241:
            _1375 <= _1360;
        242:
            _1375 <= _1361;
        243:
            _1375 <= _1362;
        244:
            _1375 <= _1363;
        245:
            _1375 <= _1364;
        246:
            _1375 <= _1365;
        247:
            _1375 <= _1366;
        248:
            _1375 <= _1367;
        249:
            _1375 <= _1368;
        250:
            _1375 <= _1369;
        251:
            _1375 <= _1370;
        252:
            _1375 <= _1371;
        253:
            _1375 <= _1372;
        254:
            _1375 <= _1373;
        default:
            _1375 <= _1374;
        endcase
    end
    assign _6243 = 8'b00000000;
    assign _6244 = _280 == _6243;
    assign _6247 = _6244 ? _6252 : _1099;
    assign _6224 = 8'b00000001;
    assign _6225 = _280 == _6224;
    assign _6228 = _6225 ? _6252 : _1099;
    assign _1398 = 8'b11111111;
    assign _1399 = _280 == _1398;
    assign _1402 = _1399 ? _6252 : _1099;
    assign _1388 = _1386 == _1398;
    assign _1389 = _1376 & _1388;
    assign _1392 = _1389 ? _1391 : _1088;
    assign _1383 = _1381 == _1398;
    assign _1384 = _1376 & _1383;
    assign _1395 = _1384 ? _1394 : _1392;
    assign _1378 = _299 == _1398;
    assign _1379 = _1376 & _1378;
    assign _1397 = _1379 ? _1099 : _1395;
    assign _1403 = _285 ? _1402 : _1397;
    assign _8 = _1403;
    always @(posedge _277) begin
        if (_275)
            _1088 <= _1099;
        else
            _1088 <= _8;
    end
    assign _1417 = 8'b11111110;
    assign _1418 = _280 == _1417;
    assign _1421 = _1418 ? _6252 : _1099;
    assign _1411 = _1386 == _1417;
    assign _1412 = _1376 & _1411;
    assign _1413 = _1412 ? _1391 : _1085;
    assign _1408 = _1381 == _1417;
    assign _1409 = _1376 & _1408;
    assign _1414 = _1409 ? _1394 : _1413;
    assign _1405 = _299 == _1417;
    assign _1406 = _1376 & _1405;
    assign _1416 = _1406 ? _1099 : _1414;
    assign _1422 = _285 ? _1421 : _1416;
    assign _9 = _1422;
    always @(posedge _277) begin
        if (_275)
            _1085 <= _1099;
        else
            _1085 <= _9;
    end
    assign _1436 = 8'b11111101;
    assign _1437 = _280 == _1436;
    assign _1440 = _1437 ? _6252 : _1099;
    assign _1430 = _1386 == _1436;
    assign _1431 = _1376 & _1430;
    assign _1432 = _1431 ? _1391 : _1082;
    assign _1427 = _1381 == _1436;
    assign _1428 = _1376 & _1427;
    assign _1433 = _1428 ? _1394 : _1432;
    assign _1424 = _299 == _1436;
    assign _1425 = _1376 & _1424;
    assign _1435 = _1425 ? _1099 : _1433;
    assign _1441 = _285 ? _1440 : _1435;
    assign _10 = _1441;
    always @(posedge _277) begin
        if (_275)
            _1082 <= _1099;
        else
            _1082 <= _10;
    end
    assign _1455 = 8'b11111100;
    assign _1456 = _280 == _1455;
    assign _1459 = _1456 ? _6252 : _1099;
    assign _1449 = _1386 == _1455;
    assign _1450 = _1376 & _1449;
    assign _1451 = _1450 ? _1391 : _1079;
    assign _1446 = _1381 == _1455;
    assign _1447 = _1376 & _1446;
    assign _1452 = _1447 ? _1394 : _1451;
    assign _1443 = _299 == _1455;
    assign _1444 = _1376 & _1443;
    assign _1454 = _1444 ? _1099 : _1452;
    assign _1460 = _285 ? _1459 : _1454;
    assign _11 = _1460;
    always @(posedge _277) begin
        if (_275)
            _1079 <= _1099;
        else
            _1079 <= _11;
    end
    assign _1474 = 8'b11111011;
    assign _1475 = _280 == _1474;
    assign _1478 = _1475 ? _6252 : _1099;
    assign _1468 = _1386 == _1474;
    assign _1469 = _1376 & _1468;
    assign _1470 = _1469 ? _1391 : _1076;
    assign _1465 = _1381 == _1474;
    assign _1466 = _1376 & _1465;
    assign _1471 = _1466 ? _1394 : _1470;
    assign _1462 = _299 == _1474;
    assign _1463 = _1376 & _1462;
    assign _1473 = _1463 ? _1099 : _1471;
    assign _1479 = _285 ? _1478 : _1473;
    assign _12 = _1479;
    always @(posedge _277) begin
        if (_275)
            _1076 <= _1099;
        else
            _1076 <= _12;
    end
    assign _1493 = 8'b11111010;
    assign _1494 = _280 == _1493;
    assign _1497 = _1494 ? _6252 : _1099;
    assign _1487 = _1386 == _1493;
    assign _1488 = _1376 & _1487;
    assign _1489 = _1488 ? _1391 : _1073;
    assign _1484 = _1381 == _1493;
    assign _1485 = _1376 & _1484;
    assign _1490 = _1485 ? _1394 : _1489;
    assign _1481 = _299 == _1493;
    assign _1482 = _1376 & _1481;
    assign _1492 = _1482 ? _1099 : _1490;
    assign _1498 = _285 ? _1497 : _1492;
    assign _13 = _1498;
    always @(posedge _277) begin
        if (_275)
            _1073 <= _1099;
        else
            _1073 <= _13;
    end
    assign _1512 = 8'b11111001;
    assign _1513 = _280 == _1512;
    assign _1516 = _1513 ? _6252 : _1099;
    assign _1506 = _1386 == _1512;
    assign _1507 = _1376 & _1506;
    assign _1508 = _1507 ? _1391 : _1070;
    assign _1503 = _1381 == _1512;
    assign _1504 = _1376 & _1503;
    assign _1509 = _1504 ? _1394 : _1508;
    assign _1500 = _299 == _1512;
    assign _1501 = _1376 & _1500;
    assign _1511 = _1501 ? _1099 : _1509;
    assign _1517 = _285 ? _1516 : _1511;
    assign _14 = _1517;
    always @(posedge _277) begin
        if (_275)
            _1070 <= _1099;
        else
            _1070 <= _14;
    end
    assign _1531 = 8'b11111000;
    assign _1532 = _280 == _1531;
    assign _1535 = _1532 ? _6252 : _1099;
    assign _1525 = _1386 == _1531;
    assign _1526 = _1376 & _1525;
    assign _1527 = _1526 ? _1391 : _1067;
    assign _1522 = _1381 == _1531;
    assign _1523 = _1376 & _1522;
    assign _1528 = _1523 ? _1394 : _1527;
    assign _1519 = _299 == _1531;
    assign _1520 = _1376 & _1519;
    assign _1530 = _1520 ? _1099 : _1528;
    assign _1536 = _285 ? _1535 : _1530;
    assign _15 = _1536;
    always @(posedge _277) begin
        if (_275)
            _1067 <= _1099;
        else
            _1067 <= _15;
    end
    assign _1550 = 8'b11110111;
    assign _1551 = _280 == _1550;
    assign _1554 = _1551 ? _6252 : _1099;
    assign _1544 = _1386 == _1550;
    assign _1545 = _1376 & _1544;
    assign _1546 = _1545 ? _1391 : _1064;
    assign _1541 = _1381 == _1550;
    assign _1542 = _1376 & _1541;
    assign _1547 = _1542 ? _1394 : _1546;
    assign _1538 = _299 == _1550;
    assign _1539 = _1376 & _1538;
    assign _1549 = _1539 ? _1099 : _1547;
    assign _1555 = _285 ? _1554 : _1549;
    assign _16 = _1555;
    always @(posedge _277) begin
        if (_275)
            _1064 <= _1099;
        else
            _1064 <= _16;
    end
    assign _1569 = 8'b11110110;
    assign _1570 = _280 == _1569;
    assign _1573 = _1570 ? _6252 : _1099;
    assign _1563 = _1386 == _1569;
    assign _1564 = _1376 & _1563;
    assign _1565 = _1564 ? _1391 : _1061;
    assign _1560 = _1381 == _1569;
    assign _1561 = _1376 & _1560;
    assign _1566 = _1561 ? _1394 : _1565;
    assign _1557 = _299 == _1569;
    assign _1558 = _1376 & _1557;
    assign _1568 = _1558 ? _1099 : _1566;
    assign _1574 = _285 ? _1573 : _1568;
    assign _17 = _1574;
    always @(posedge _277) begin
        if (_275)
            _1061 <= _1099;
        else
            _1061 <= _17;
    end
    assign _1588 = 8'b11110101;
    assign _1589 = _280 == _1588;
    assign _1592 = _1589 ? _6252 : _1099;
    assign _1582 = _1386 == _1588;
    assign _1583 = _1376 & _1582;
    assign _1584 = _1583 ? _1391 : _1058;
    assign _1579 = _1381 == _1588;
    assign _1580 = _1376 & _1579;
    assign _1585 = _1580 ? _1394 : _1584;
    assign _1576 = _299 == _1588;
    assign _1577 = _1376 & _1576;
    assign _1587 = _1577 ? _1099 : _1585;
    assign _1593 = _285 ? _1592 : _1587;
    assign _18 = _1593;
    always @(posedge _277) begin
        if (_275)
            _1058 <= _1099;
        else
            _1058 <= _18;
    end
    assign _1607 = 8'b11110100;
    assign _1608 = _280 == _1607;
    assign _1611 = _1608 ? _6252 : _1099;
    assign _1601 = _1386 == _1607;
    assign _1602 = _1376 & _1601;
    assign _1603 = _1602 ? _1391 : _1055;
    assign _1598 = _1381 == _1607;
    assign _1599 = _1376 & _1598;
    assign _1604 = _1599 ? _1394 : _1603;
    assign _1595 = _299 == _1607;
    assign _1596 = _1376 & _1595;
    assign _1606 = _1596 ? _1099 : _1604;
    assign _1612 = _285 ? _1611 : _1606;
    assign _19 = _1612;
    always @(posedge _277) begin
        if (_275)
            _1055 <= _1099;
        else
            _1055 <= _19;
    end
    assign _1626 = 8'b11110011;
    assign _1627 = _280 == _1626;
    assign _1630 = _1627 ? _6252 : _1099;
    assign _1620 = _1386 == _1626;
    assign _1621 = _1376 & _1620;
    assign _1622 = _1621 ? _1391 : _1052;
    assign _1617 = _1381 == _1626;
    assign _1618 = _1376 & _1617;
    assign _1623 = _1618 ? _1394 : _1622;
    assign _1614 = _299 == _1626;
    assign _1615 = _1376 & _1614;
    assign _1625 = _1615 ? _1099 : _1623;
    assign _1631 = _285 ? _1630 : _1625;
    assign _20 = _1631;
    always @(posedge _277) begin
        if (_275)
            _1052 <= _1099;
        else
            _1052 <= _20;
    end
    assign _1645 = 8'b11110010;
    assign _1646 = _280 == _1645;
    assign _1649 = _1646 ? _6252 : _1099;
    assign _1639 = _1386 == _1645;
    assign _1640 = _1376 & _1639;
    assign _1641 = _1640 ? _1391 : _1049;
    assign _1636 = _1381 == _1645;
    assign _1637 = _1376 & _1636;
    assign _1642 = _1637 ? _1394 : _1641;
    assign _1633 = _299 == _1645;
    assign _1634 = _1376 & _1633;
    assign _1644 = _1634 ? _1099 : _1642;
    assign _1650 = _285 ? _1649 : _1644;
    assign _21 = _1650;
    always @(posedge _277) begin
        if (_275)
            _1049 <= _1099;
        else
            _1049 <= _21;
    end
    assign _1664 = 8'b11110001;
    assign _1665 = _280 == _1664;
    assign _1668 = _1665 ? _6252 : _1099;
    assign _1658 = _1386 == _1664;
    assign _1659 = _1376 & _1658;
    assign _1660 = _1659 ? _1391 : _1046;
    assign _1655 = _1381 == _1664;
    assign _1656 = _1376 & _1655;
    assign _1661 = _1656 ? _1394 : _1660;
    assign _1652 = _299 == _1664;
    assign _1653 = _1376 & _1652;
    assign _1663 = _1653 ? _1099 : _1661;
    assign _1669 = _285 ? _1668 : _1663;
    assign _22 = _1669;
    always @(posedge _277) begin
        if (_275)
            _1046 <= _1099;
        else
            _1046 <= _22;
    end
    assign _1683 = 8'b11110000;
    assign _1684 = _280 == _1683;
    assign _1687 = _1684 ? _6252 : _1099;
    assign _1677 = _1386 == _1683;
    assign _1678 = _1376 & _1677;
    assign _1679 = _1678 ? _1391 : _1043;
    assign _1674 = _1381 == _1683;
    assign _1675 = _1376 & _1674;
    assign _1680 = _1675 ? _1394 : _1679;
    assign _1671 = _299 == _1683;
    assign _1672 = _1376 & _1671;
    assign _1682 = _1672 ? _1099 : _1680;
    assign _1688 = _285 ? _1687 : _1682;
    assign _23 = _1688;
    always @(posedge _277) begin
        if (_275)
            _1043 <= _1099;
        else
            _1043 <= _23;
    end
    assign _1702 = 8'b11101111;
    assign _1703 = _280 == _1702;
    assign _1706 = _1703 ? _6252 : _1099;
    assign _1696 = _1386 == _1702;
    assign _1697 = _1376 & _1696;
    assign _1698 = _1697 ? _1391 : _1040;
    assign _1693 = _1381 == _1702;
    assign _1694 = _1376 & _1693;
    assign _1699 = _1694 ? _1394 : _1698;
    assign _1690 = _299 == _1702;
    assign _1691 = _1376 & _1690;
    assign _1701 = _1691 ? _1099 : _1699;
    assign _1707 = _285 ? _1706 : _1701;
    assign _24 = _1707;
    always @(posedge _277) begin
        if (_275)
            _1040 <= _1099;
        else
            _1040 <= _24;
    end
    assign _1721 = 8'b11101110;
    assign _1722 = _280 == _1721;
    assign _1725 = _1722 ? _6252 : _1099;
    assign _1715 = _1386 == _1721;
    assign _1716 = _1376 & _1715;
    assign _1717 = _1716 ? _1391 : _1037;
    assign _1712 = _1381 == _1721;
    assign _1713 = _1376 & _1712;
    assign _1718 = _1713 ? _1394 : _1717;
    assign _1709 = _299 == _1721;
    assign _1710 = _1376 & _1709;
    assign _1720 = _1710 ? _1099 : _1718;
    assign _1726 = _285 ? _1725 : _1720;
    assign _25 = _1726;
    always @(posedge _277) begin
        if (_275)
            _1037 <= _1099;
        else
            _1037 <= _25;
    end
    assign _1740 = 8'b11101101;
    assign _1741 = _280 == _1740;
    assign _1744 = _1741 ? _6252 : _1099;
    assign _1734 = _1386 == _1740;
    assign _1735 = _1376 & _1734;
    assign _1736 = _1735 ? _1391 : _1034;
    assign _1731 = _1381 == _1740;
    assign _1732 = _1376 & _1731;
    assign _1737 = _1732 ? _1394 : _1736;
    assign _1728 = _299 == _1740;
    assign _1729 = _1376 & _1728;
    assign _1739 = _1729 ? _1099 : _1737;
    assign _1745 = _285 ? _1744 : _1739;
    assign _26 = _1745;
    always @(posedge _277) begin
        if (_275)
            _1034 <= _1099;
        else
            _1034 <= _26;
    end
    assign _1759 = 8'b11101100;
    assign _1760 = _280 == _1759;
    assign _1763 = _1760 ? _6252 : _1099;
    assign _1753 = _1386 == _1759;
    assign _1754 = _1376 & _1753;
    assign _1755 = _1754 ? _1391 : _1031;
    assign _1750 = _1381 == _1759;
    assign _1751 = _1376 & _1750;
    assign _1756 = _1751 ? _1394 : _1755;
    assign _1747 = _299 == _1759;
    assign _1748 = _1376 & _1747;
    assign _1758 = _1748 ? _1099 : _1756;
    assign _1764 = _285 ? _1763 : _1758;
    assign _27 = _1764;
    always @(posedge _277) begin
        if (_275)
            _1031 <= _1099;
        else
            _1031 <= _27;
    end
    assign _1778 = 8'b11101011;
    assign _1779 = _280 == _1778;
    assign _1782 = _1779 ? _6252 : _1099;
    assign _1772 = _1386 == _1778;
    assign _1773 = _1376 & _1772;
    assign _1774 = _1773 ? _1391 : _1028;
    assign _1769 = _1381 == _1778;
    assign _1770 = _1376 & _1769;
    assign _1775 = _1770 ? _1394 : _1774;
    assign _1766 = _299 == _1778;
    assign _1767 = _1376 & _1766;
    assign _1777 = _1767 ? _1099 : _1775;
    assign _1783 = _285 ? _1782 : _1777;
    assign _28 = _1783;
    always @(posedge _277) begin
        if (_275)
            _1028 <= _1099;
        else
            _1028 <= _28;
    end
    assign _1797 = 8'b11101010;
    assign _1798 = _280 == _1797;
    assign _1801 = _1798 ? _6252 : _1099;
    assign _1791 = _1386 == _1797;
    assign _1792 = _1376 & _1791;
    assign _1793 = _1792 ? _1391 : _1025;
    assign _1788 = _1381 == _1797;
    assign _1789 = _1376 & _1788;
    assign _1794 = _1789 ? _1394 : _1793;
    assign _1785 = _299 == _1797;
    assign _1786 = _1376 & _1785;
    assign _1796 = _1786 ? _1099 : _1794;
    assign _1802 = _285 ? _1801 : _1796;
    assign _29 = _1802;
    always @(posedge _277) begin
        if (_275)
            _1025 <= _1099;
        else
            _1025 <= _29;
    end
    assign _1816 = 8'b11101001;
    assign _1817 = _280 == _1816;
    assign _1820 = _1817 ? _6252 : _1099;
    assign _1810 = _1386 == _1816;
    assign _1811 = _1376 & _1810;
    assign _1812 = _1811 ? _1391 : _1022;
    assign _1807 = _1381 == _1816;
    assign _1808 = _1376 & _1807;
    assign _1813 = _1808 ? _1394 : _1812;
    assign _1804 = _299 == _1816;
    assign _1805 = _1376 & _1804;
    assign _1815 = _1805 ? _1099 : _1813;
    assign _1821 = _285 ? _1820 : _1815;
    assign _30 = _1821;
    always @(posedge _277) begin
        if (_275)
            _1022 <= _1099;
        else
            _1022 <= _30;
    end
    assign _1835 = 8'b11101000;
    assign _1836 = _280 == _1835;
    assign _1839 = _1836 ? _6252 : _1099;
    assign _1829 = _1386 == _1835;
    assign _1830 = _1376 & _1829;
    assign _1831 = _1830 ? _1391 : _1019;
    assign _1826 = _1381 == _1835;
    assign _1827 = _1376 & _1826;
    assign _1832 = _1827 ? _1394 : _1831;
    assign _1823 = _299 == _1835;
    assign _1824 = _1376 & _1823;
    assign _1834 = _1824 ? _1099 : _1832;
    assign _1840 = _285 ? _1839 : _1834;
    assign _31 = _1840;
    always @(posedge _277) begin
        if (_275)
            _1019 <= _1099;
        else
            _1019 <= _31;
    end
    assign _1854 = 8'b11100111;
    assign _1855 = _280 == _1854;
    assign _1858 = _1855 ? _6252 : _1099;
    assign _1848 = _1386 == _1854;
    assign _1849 = _1376 & _1848;
    assign _1850 = _1849 ? _1391 : _1016;
    assign _1845 = _1381 == _1854;
    assign _1846 = _1376 & _1845;
    assign _1851 = _1846 ? _1394 : _1850;
    assign _1842 = _299 == _1854;
    assign _1843 = _1376 & _1842;
    assign _1853 = _1843 ? _1099 : _1851;
    assign _1859 = _285 ? _1858 : _1853;
    assign _32 = _1859;
    always @(posedge _277) begin
        if (_275)
            _1016 <= _1099;
        else
            _1016 <= _32;
    end
    assign _1873 = 8'b11100110;
    assign _1874 = _280 == _1873;
    assign _1877 = _1874 ? _6252 : _1099;
    assign _1867 = _1386 == _1873;
    assign _1868 = _1376 & _1867;
    assign _1869 = _1868 ? _1391 : _1013;
    assign _1864 = _1381 == _1873;
    assign _1865 = _1376 & _1864;
    assign _1870 = _1865 ? _1394 : _1869;
    assign _1861 = _299 == _1873;
    assign _1862 = _1376 & _1861;
    assign _1872 = _1862 ? _1099 : _1870;
    assign _1878 = _285 ? _1877 : _1872;
    assign _33 = _1878;
    always @(posedge _277) begin
        if (_275)
            _1013 <= _1099;
        else
            _1013 <= _33;
    end
    assign _1892 = 8'b11100101;
    assign _1893 = _280 == _1892;
    assign _1896 = _1893 ? _6252 : _1099;
    assign _1886 = _1386 == _1892;
    assign _1887 = _1376 & _1886;
    assign _1888 = _1887 ? _1391 : _1010;
    assign _1883 = _1381 == _1892;
    assign _1884 = _1376 & _1883;
    assign _1889 = _1884 ? _1394 : _1888;
    assign _1880 = _299 == _1892;
    assign _1881 = _1376 & _1880;
    assign _1891 = _1881 ? _1099 : _1889;
    assign _1897 = _285 ? _1896 : _1891;
    assign _34 = _1897;
    always @(posedge _277) begin
        if (_275)
            _1010 <= _1099;
        else
            _1010 <= _34;
    end
    assign _1911 = 8'b11100100;
    assign _1912 = _280 == _1911;
    assign _1915 = _1912 ? _6252 : _1099;
    assign _1905 = _1386 == _1911;
    assign _1906 = _1376 & _1905;
    assign _1907 = _1906 ? _1391 : _1007;
    assign _1902 = _1381 == _1911;
    assign _1903 = _1376 & _1902;
    assign _1908 = _1903 ? _1394 : _1907;
    assign _1899 = _299 == _1911;
    assign _1900 = _1376 & _1899;
    assign _1910 = _1900 ? _1099 : _1908;
    assign _1916 = _285 ? _1915 : _1910;
    assign _35 = _1916;
    always @(posedge _277) begin
        if (_275)
            _1007 <= _1099;
        else
            _1007 <= _35;
    end
    assign _1930 = 8'b11100011;
    assign _1931 = _280 == _1930;
    assign _1934 = _1931 ? _6252 : _1099;
    assign _1924 = _1386 == _1930;
    assign _1925 = _1376 & _1924;
    assign _1926 = _1925 ? _1391 : _1004;
    assign _1921 = _1381 == _1930;
    assign _1922 = _1376 & _1921;
    assign _1927 = _1922 ? _1394 : _1926;
    assign _1918 = _299 == _1930;
    assign _1919 = _1376 & _1918;
    assign _1929 = _1919 ? _1099 : _1927;
    assign _1935 = _285 ? _1934 : _1929;
    assign _36 = _1935;
    always @(posedge _277) begin
        if (_275)
            _1004 <= _1099;
        else
            _1004 <= _36;
    end
    assign _1949 = 8'b11100010;
    assign _1950 = _280 == _1949;
    assign _1953 = _1950 ? _6252 : _1099;
    assign _1943 = _1386 == _1949;
    assign _1944 = _1376 & _1943;
    assign _1945 = _1944 ? _1391 : _1001;
    assign _1940 = _1381 == _1949;
    assign _1941 = _1376 & _1940;
    assign _1946 = _1941 ? _1394 : _1945;
    assign _1937 = _299 == _1949;
    assign _1938 = _1376 & _1937;
    assign _1948 = _1938 ? _1099 : _1946;
    assign _1954 = _285 ? _1953 : _1948;
    assign _37 = _1954;
    always @(posedge _277) begin
        if (_275)
            _1001 <= _1099;
        else
            _1001 <= _37;
    end
    assign _1968 = 8'b11100001;
    assign _1969 = _280 == _1968;
    assign _1972 = _1969 ? _6252 : _1099;
    assign _1962 = _1386 == _1968;
    assign _1963 = _1376 & _1962;
    assign _1964 = _1963 ? _1391 : _998;
    assign _1959 = _1381 == _1968;
    assign _1960 = _1376 & _1959;
    assign _1965 = _1960 ? _1394 : _1964;
    assign _1956 = _299 == _1968;
    assign _1957 = _1376 & _1956;
    assign _1967 = _1957 ? _1099 : _1965;
    assign _1973 = _285 ? _1972 : _1967;
    assign _38 = _1973;
    always @(posedge _277) begin
        if (_275)
            _998 <= _1099;
        else
            _998 <= _38;
    end
    assign _1987 = 8'b11100000;
    assign _1988 = _280 == _1987;
    assign _1991 = _1988 ? _6252 : _1099;
    assign _1981 = _1386 == _1987;
    assign _1982 = _1376 & _1981;
    assign _1983 = _1982 ? _1391 : _995;
    assign _1978 = _1381 == _1987;
    assign _1979 = _1376 & _1978;
    assign _1984 = _1979 ? _1394 : _1983;
    assign _1975 = _299 == _1987;
    assign _1976 = _1376 & _1975;
    assign _1986 = _1976 ? _1099 : _1984;
    assign _1992 = _285 ? _1991 : _1986;
    assign _39 = _1992;
    always @(posedge _277) begin
        if (_275)
            _995 <= _1099;
        else
            _995 <= _39;
    end
    assign _2006 = 8'b11011111;
    assign _2007 = _280 == _2006;
    assign _2010 = _2007 ? _6252 : _1099;
    assign _2000 = _1386 == _2006;
    assign _2001 = _1376 & _2000;
    assign _2002 = _2001 ? _1391 : _992;
    assign _1997 = _1381 == _2006;
    assign _1998 = _1376 & _1997;
    assign _2003 = _1998 ? _1394 : _2002;
    assign _1994 = _299 == _2006;
    assign _1995 = _1376 & _1994;
    assign _2005 = _1995 ? _1099 : _2003;
    assign _2011 = _285 ? _2010 : _2005;
    assign _40 = _2011;
    always @(posedge _277) begin
        if (_275)
            _992 <= _1099;
        else
            _992 <= _40;
    end
    assign _2025 = 8'b11011110;
    assign _2026 = _280 == _2025;
    assign _2029 = _2026 ? _6252 : _1099;
    assign _2019 = _1386 == _2025;
    assign _2020 = _1376 & _2019;
    assign _2021 = _2020 ? _1391 : _989;
    assign _2016 = _1381 == _2025;
    assign _2017 = _1376 & _2016;
    assign _2022 = _2017 ? _1394 : _2021;
    assign _2013 = _299 == _2025;
    assign _2014 = _1376 & _2013;
    assign _2024 = _2014 ? _1099 : _2022;
    assign _2030 = _285 ? _2029 : _2024;
    assign _41 = _2030;
    always @(posedge _277) begin
        if (_275)
            _989 <= _1099;
        else
            _989 <= _41;
    end
    assign _2044 = 8'b11011101;
    assign _2045 = _280 == _2044;
    assign _2048 = _2045 ? _6252 : _1099;
    assign _2038 = _1386 == _2044;
    assign _2039 = _1376 & _2038;
    assign _2040 = _2039 ? _1391 : _986;
    assign _2035 = _1381 == _2044;
    assign _2036 = _1376 & _2035;
    assign _2041 = _2036 ? _1394 : _2040;
    assign _2032 = _299 == _2044;
    assign _2033 = _1376 & _2032;
    assign _2043 = _2033 ? _1099 : _2041;
    assign _2049 = _285 ? _2048 : _2043;
    assign _42 = _2049;
    always @(posedge _277) begin
        if (_275)
            _986 <= _1099;
        else
            _986 <= _42;
    end
    assign _2063 = 8'b11011100;
    assign _2064 = _280 == _2063;
    assign _2067 = _2064 ? _6252 : _1099;
    assign _2057 = _1386 == _2063;
    assign _2058 = _1376 & _2057;
    assign _2059 = _2058 ? _1391 : _983;
    assign _2054 = _1381 == _2063;
    assign _2055 = _1376 & _2054;
    assign _2060 = _2055 ? _1394 : _2059;
    assign _2051 = _299 == _2063;
    assign _2052 = _1376 & _2051;
    assign _2062 = _2052 ? _1099 : _2060;
    assign _2068 = _285 ? _2067 : _2062;
    assign _43 = _2068;
    always @(posedge _277) begin
        if (_275)
            _983 <= _1099;
        else
            _983 <= _43;
    end
    assign _2082 = 8'b11011011;
    assign _2083 = _280 == _2082;
    assign _2086 = _2083 ? _6252 : _1099;
    assign _2076 = _1386 == _2082;
    assign _2077 = _1376 & _2076;
    assign _2078 = _2077 ? _1391 : _980;
    assign _2073 = _1381 == _2082;
    assign _2074 = _1376 & _2073;
    assign _2079 = _2074 ? _1394 : _2078;
    assign _2070 = _299 == _2082;
    assign _2071 = _1376 & _2070;
    assign _2081 = _2071 ? _1099 : _2079;
    assign _2087 = _285 ? _2086 : _2081;
    assign _44 = _2087;
    always @(posedge _277) begin
        if (_275)
            _980 <= _1099;
        else
            _980 <= _44;
    end
    assign _2101 = 8'b11011010;
    assign _2102 = _280 == _2101;
    assign _2105 = _2102 ? _6252 : _1099;
    assign _2095 = _1386 == _2101;
    assign _2096 = _1376 & _2095;
    assign _2097 = _2096 ? _1391 : _977;
    assign _2092 = _1381 == _2101;
    assign _2093 = _1376 & _2092;
    assign _2098 = _2093 ? _1394 : _2097;
    assign _2089 = _299 == _2101;
    assign _2090 = _1376 & _2089;
    assign _2100 = _2090 ? _1099 : _2098;
    assign _2106 = _285 ? _2105 : _2100;
    assign _45 = _2106;
    always @(posedge _277) begin
        if (_275)
            _977 <= _1099;
        else
            _977 <= _45;
    end
    assign _2120 = 8'b11011001;
    assign _2121 = _280 == _2120;
    assign _2124 = _2121 ? _6252 : _1099;
    assign _2114 = _1386 == _2120;
    assign _2115 = _1376 & _2114;
    assign _2116 = _2115 ? _1391 : _974;
    assign _2111 = _1381 == _2120;
    assign _2112 = _1376 & _2111;
    assign _2117 = _2112 ? _1394 : _2116;
    assign _2108 = _299 == _2120;
    assign _2109 = _1376 & _2108;
    assign _2119 = _2109 ? _1099 : _2117;
    assign _2125 = _285 ? _2124 : _2119;
    assign _46 = _2125;
    always @(posedge _277) begin
        if (_275)
            _974 <= _1099;
        else
            _974 <= _46;
    end
    assign _2139 = 8'b11011000;
    assign _2140 = _280 == _2139;
    assign _2143 = _2140 ? _6252 : _1099;
    assign _2133 = _1386 == _2139;
    assign _2134 = _1376 & _2133;
    assign _2135 = _2134 ? _1391 : _971;
    assign _2130 = _1381 == _2139;
    assign _2131 = _1376 & _2130;
    assign _2136 = _2131 ? _1394 : _2135;
    assign _2127 = _299 == _2139;
    assign _2128 = _1376 & _2127;
    assign _2138 = _2128 ? _1099 : _2136;
    assign _2144 = _285 ? _2143 : _2138;
    assign _47 = _2144;
    always @(posedge _277) begin
        if (_275)
            _971 <= _1099;
        else
            _971 <= _47;
    end
    assign _2158 = 8'b11010111;
    assign _2159 = _280 == _2158;
    assign _2162 = _2159 ? _6252 : _1099;
    assign _2152 = _1386 == _2158;
    assign _2153 = _1376 & _2152;
    assign _2154 = _2153 ? _1391 : _968;
    assign _2149 = _1381 == _2158;
    assign _2150 = _1376 & _2149;
    assign _2155 = _2150 ? _1394 : _2154;
    assign _2146 = _299 == _2158;
    assign _2147 = _1376 & _2146;
    assign _2157 = _2147 ? _1099 : _2155;
    assign _2163 = _285 ? _2162 : _2157;
    assign _48 = _2163;
    always @(posedge _277) begin
        if (_275)
            _968 <= _1099;
        else
            _968 <= _48;
    end
    assign _2177 = 8'b11010110;
    assign _2178 = _280 == _2177;
    assign _2181 = _2178 ? _6252 : _1099;
    assign _2171 = _1386 == _2177;
    assign _2172 = _1376 & _2171;
    assign _2173 = _2172 ? _1391 : _965;
    assign _2168 = _1381 == _2177;
    assign _2169 = _1376 & _2168;
    assign _2174 = _2169 ? _1394 : _2173;
    assign _2165 = _299 == _2177;
    assign _2166 = _1376 & _2165;
    assign _2176 = _2166 ? _1099 : _2174;
    assign _2182 = _285 ? _2181 : _2176;
    assign _49 = _2182;
    always @(posedge _277) begin
        if (_275)
            _965 <= _1099;
        else
            _965 <= _49;
    end
    assign _2196 = 8'b11010101;
    assign _2197 = _280 == _2196;
    assign _2200 = _2197 ? _6252 : _1099;
    assign _2190 = _1386 == _2196;
    assign _2191 = _1376 & _2190;
    assign _2192 = _2191 ? _1391 : _962;
    assign _2187 = _1381 == _2196;
    assign _2188 = _1376 & _2187;
    assign _2193 = _2188 ? _1394 : _2192;
    assign _2184 = _299 == _2196;
    assign _2185 = _1376 & _2184;
    assign _2195 = _2185 ? _1099 : _2193;
    assign _2201 = _285 ? _2200 : _2195;
    assign _50 = _2201;
    always @(posedge _277) begin
        if (_275)
            _962 <= _1099;
        else
            _962 <= _50;
    end
    assign _2215 = 8'b11010100;
    assign _2216 = _280 == _2215;
    assign _2219 = _2216 ? _6252 : _1099;
    assign _2209 = _1386 == _2215;
    assign _2210 = _1376 & _2209;
    assign _2211 = _2210 ? _1391 : _959;
    assign _2206 = _1381 == _2215;
    assign _2207 = _1376 & _2206;
    assign _2212 = _2207 ? _1394 : _2211;
    assign _2203 = _299 == _2215;
    assign _2204 = _1376 & _2203;
    assign _2214 = _2204 ? _1099 : _2212;
    assign _2220 = _285 ? _2219 : _2214;
    assign _51 = _2220;
    always @(posedge _277) begin
        if (_275)
            _959 <= _1099;
        else
            _959 <= _51;
    end
    assign _2234 = 8'b11010011;
    assign _2235 = _280 == _2234;
    assign _2238 = _2235 ? _6252 : _1099;
    assign _2228 = _1386 == _2234;
    assign _2229 = _1376 & _2228;
    assign _2230 = _2229 ? _1391 : _956;
    assign _2225 = _1381 == _2234;
    assign _2226 = _1376 & _2225;
    assign _2231 = _2226 ? _1394 : _2230;
    assign _2222 = _299 == _2234;
    assign _2223 = _1376 & _2222;
    assign _2233 = _2223 ? _1099 : _2231;
    assign _2239 = _285 ? _2238 : _2233;
    assign _52 = _2239;
    always @(posedge _277) begin
        if (_275)
            _956 <= _1099;
        else
            _956 <= _52;
    end
    assign _2253 = 8'b11010010;
    assign _2254 = _280 == _2253;
    assign _2257 = _2254 ? _6252 : _1099;
    assign _2247 = _1386 == _2253;
    assign _2248 = _1376 & _2247;
    assign _2249 = _2248 ? _1391 : _953;
    assign _2244 = _1381 == _2253;
    assign _2245 = _1376 & _2244;
    assign _2250 = _2245 ? _1394 : _2249;
    assign _2241 = _299 == _2253;
    assign _2242 = _1376 & _2241;
    assign _2252 = _2242 ? _1099 : _2250;
    assign _2258 = _285 ? _2257 : _2252;
    assign _53 = _2258;
    always @(posedge _277) begin
        if (_275)
            _953 <= _1099;
        else
            _953 <= _53;
    end
    assign _2272 = 8'b11010001;
    assign _2273 = _280 == _2272;
    assign _2276 = _2273 ? _6252 : _1099;
    assign _2266 = _1386 == _2272;
    assign _2267 = _1376 & _2266;
    assign _2268 = _2267 ? _1391 : _950;
    assign _2263 = _1381 == _2272;
    assign _2264 = _1376 & _2263;
    assign _2269 = _2264 ? _1394 : _2268;
    assign _2260 = _299 == _2272;
    assign _2261 = _1376 & _2260;
    assign _2271 = _2261 ? _1099 : _2269;
    assign _2277 = _285 ? _2276 : _2271;
    assign _54 = _2277;
    always @(posedge _277) begin
        if (_275)
            _950 <= _1099;
        else
            _950 <= _54;
    end
    assign _2291 = 8'b11010000;
    assign _2292 = _280 == _2291;
    assign _2295 = _2292 ? _6252 : _1099;
    assign _2285 = _1386 == _2291;
    assign _2286 = _1376 & _2285;
    assign _2287 = _2286 ? _1391 : _947;
    assign _2282 = _1381 == _2291;
    assign _2283 = _1376 & _2282;
    assign _2288 = _2283 ? _1394 : _2287;
    assign _2279 = _299 == _2291;
    assign _2280 = _1376 & _2279;
    assign _2290 = _2280 ? _1099 : _2288;
    assign _2296 = _285 ? _2295 : _2290;
    assign _55 = _2296;
    always @(posedge _277) begin
        if (_275)
            _947 <= _1099;
        else
            _947 <= _55;
    end
    assign _2310 = 8'b11001111;
    assign _2311 = _280 == _2310;
    assign _2314 = _2311 ? _6252 : _1099;
    assign _2304 = _1386 == _2310;
    assign _2305 = _1376 & _2304;
    assign _2306 = _2305 ? _1391 : _944;
    assign _2301 = _1381 == _2310;
    assign _2302 = _1376 & _2301;
    assign _2307 = _2302 ? _1394 : _2306;
    assign _2298 = _299 == _2310;
    assign _2299 = _1376 & _2298;
    assign _2309 = _2299 ? _1099 : _2307;
    assign _2315 = _285 ? _2314 : _2309;
    assign _56 = _2315;
    always @(posedge _277) begin
        if (_275)
            _944 <= _1099;
        else
            _944 <= _56;
    end
    assign _2329 = 8'b11001110;
    assign _2330 = _280 == _2329;
    assign _2333 = _2330 ? _6252 : _1099;
    assign _2323 = _1386 == _2329;
    assign _2324 = _1376 & _2323;
    assign _2325 = _2324 ? _1391 : _941;
    assign _2320 = _1381 == _2329;
    assign _2321 = _1376 & _2320;
    assign _2326 = _2321 ? _1394 : _2325;
    assign _2317 = _299 == _2329;
    assign _2318 = _1376 & _2317;
    assign _2328 = _2318 ? _1099 : _2326;
    assign _2334 = _285 ? _2333 : _2328;
    assign _57 = _2334;
    always @(posedge _277) begin
        if (_275)
            _941 <= _1099;
        else
            _941 <= _57;
    end
    assign _2348 = 8'b11001101;
    assign _2349 = _280 == _2348;
    assign _2352 = _2349 ? _6252 : _1099;
    assign _2342 = _1386 == _2348;
    assign _2343 = _1376 & _2342;
    assign _2344 = _2343 ? _1391 : _938;
    assign _2339 = _1381 == _2348;
    assign _2340 = _1376 & _2339;
    assign _2345 = _2340 ? _1394 : _2344;
    assign _2336 = _299 == _2348;
    assign _2337 = _1376 & _2336;
    assign _2347 = _2337 ? _1099 : _2345;
    assign _2353 = _285 ? _2352 : _2347;
    assign _58 = _2353;
    always @(posedge _277) begin
        if (_275)
            _938 <= _1099;
        else
            _938 <= _58;
    end
    assign _2367 = 8'b11001100;
    assign _2368 = _280 == _2367;
    assign _2371 = _2368 ? _6252 : _1099;
    assign _2361 = _1386 == _2367;
    assign _2362 = _1376 & _2361;
    assign _2363 = _2362 ? _1391 : _935;
    assign _2358 = _1381 == _2367;
    assign _2359 = _1376 & _2358;
    assign _2364 = _2359 ? _1394 : _2363;
    assign _2355 = _299 == _2367;
    assign _2356 = _1376 & _2355;
    assign _2366 = _2356 ? _1099 : _2364;
    assign _2372 = _285 ? _2371 : _2366;
    assign _59 = _2372;
    always @(posedge _277) begin
        if (_275)
            _935 <= _1099;
        else
            _935 <= _59;
    end
    assign _2386 = 8'b11001011;
    assign _2387 = _280 == _2386;
    assign _2390 = _2387 ? _6252 : _1099;
    assign _2380 = _1386 == _2386;
    assign _2381 = _1376 & _2380;
    assign _2382 = _2381 ? _1391 : _932;
    assign _2377 = _1381 == _2386;
    assign _2378 = _1376 & _2377;
    assign _2383 = _2378 ? _1394 : _2382;
    assign _2374 = _299 == _2386;
    assign _2375 = _1376 & _2374;
    assign _2385 = _2375 ? _1099 : _2383;
    assign _2391 = _285 ? _2390 : _2385;
    assign _60 = _2391;
    always @(posedge _277) begin
        if (_275)
            _932 <= _1099;
        else
            _932 <= _60;
    end
    assign _2405 = 8'b11001010;
    assign _2406 = _280 == _2405;
    assign _2409 = _2406 ? _6252 : _1099;
    assign _2399 = _1386 == _2405;
    assign _2400 = _1376 & _2399;
    assign _2401 = _2400 ? _1391 : _929;
    assign _2396 = _1381 == _2405;
    assign _2397 = _1376 & _2396;
    assign _2402 = _2397 ? _1394 : _2401;
    assign _2393 = _299 == _2405;
    assign _2394 = _1376 & _2393;
    assign _2404 = _2394 ? _1099 : _2402;
    assign _2410 = _285 ? _2409 : _2404;
    assign _61 = _2410;
    always @(posedge _277) begin
        if (_275)
            _929 <= _1099;
        else
            _929 <= _61;
    end
    assign _2424 = 8'b11001001;
    assign _2425 = _280 == _2424;
    assign _2428 = _2425 ? _6252 : _1099;
    assign _2418 = _1386 == _2424;
    assign _2419 = _1376 & _2418;
    assign _2420 = _2419 ? _1391 : _926;
    assign _2415 = _1381 == _2424;
    assign _2416 = _1376 & _2415;
    assign _2421 = _2416 ? _1394 : _2420;
    assign _2412 = _299 == _2424;
    assign _2413 = _1376 & _2412;
    assign _2423 = _2413 ? _1099 : _2421;
    assign _2429 = _285 ? _2428 : _2423;
    assign _62 = _2429;
    always @(posedge _277) begin
        if (_275)
            _926 <= _1099;
        else
            _926 <= _62;
    end
    assign _2443 = 8'b11001000;
    assign _2444 = _280 == _2443;
    assign _2447 = _2444 ? _6252 : _1099;
    assign _2437 = _1386 == _2443;
    assign _2438 = _1376 & _2437;
    assign _2439 = _2438 ? _1391 : _923;
    assign _2434 = _1381 == _2443;
    assign _2435 = _1376 & _2434;
    assign _2440 = _2435 ? _1394 : _2439;
    assign _2431 = _299 == _2443;
    assign _2432 = _1376 & _2431;
    assign _2442 = _2432 ? _1099 : _2440;
    assign _2448 = _285 ? _2447 : _2442;
    assign _63 = _2448;
    always @(posedge _277) begin
        if (_275)
            _923 <= _1099;
        else
            _923 <= _63;
    end
    assign _2462 = 8'b11000111;
    assign _2463 = _280 == _2462;
    assign _2466 = _2463 ? _6252 : _1099;
    assign _2456 = _1386 == _2462;
    assign _2457 = _1376 & _2456;
    assign _2458 = _2457 ? _1391 : _920;
    assign _2453 = _1381 == _2462;
    assign _2454 = _1376 & _2453;
    assign _2459 = _2454 ? _1394 : _2458;
    assign _2450 = _299 == _2462;
    assign _2451 = _1376 & _2450;
    assign _2461 = _2451 ? _1099 : _2459;
    assign _2467 = _285 ? _2466 : _2461;
    assign _64 = _2467;
    always @(posedge _277) begin
        if (_275)
            _920 <= _1099;
        else
            _920 <= _64;
    end
    assign _2481 = 8'b11000110;
    assign _2482 = _280 == _2481;
    assign _2485 = _2482 ? _6252 : _1099;
    assign _2475 = _1386 == _2481;
    assign _2476 = _1376 & _2475;
    assign _2477 = _2476 ? _1391 : _917;
    assign _2472 = _1381 == _2481;
    assign _2473 = _1376 & _2472;
    assign _2478 = _2473 ? _1394 : _2477;
    assign _2469 = _299 == _2481;
    assign _2470 = _1376 & _2469;
    assign _2480 = _2470 ? _1099 : _2478;
    assign _2486 = _285 ? _2485 : _2480;
    assign _65 = _2486;
    always @(posedge _277) begin
        if (_275)
            _917 <= _1099;
        else
            _917 <= _65;
    end
    assign _2500 = 8'b11000101;
    assign _2501 = _280 == _2500;
    assign _2504 = _2501 ? _6252 : _1099;
    assign _2494 = _1386 == _2500;
    assign _2495 = _1376 & _2494;
    assign _2496 = _2495 ? _1391 : _914;
    assign _2491 = _1381 == _2500;
    assign _2492 = _1376 & _2491;
    assign _2497 = _2492 ? _1394 : _2496;
    assign _2488 = _299 == _2500;
    assign _2489 = _1376 & _2488;
    assign _2499 = _2489 ? _1099 : _2497;
    assign _2505 = _285 ? _2504 : _2499;
    assign _66 = _2505;
    always @(posedge _277) begin
        if (_275)
            _914 <= _1099;
        else
            _914 <= _66;
    end
    assign _2519 = 8'b11000100;
    assign _2520 = _280 == _2519;
    assign _2523 = _2520 ? _6252 : _1099;
    assign _2513 = _1386 == _2519;
    assign _2514 = _1376 & _2513;
    assign _2515 = _2514 ? _1391 : _911;
    assign _2510 = _1381 == _2519;
    assign _2511 = _1376 & _2510;
    assign _2516 = _2511 ? _1394 : _2515;
    assign _2507 = _299 == _2519;
    assign _2508 = _1376 & _2507;
    assign _2518 = _2508 ? _1099 : _2516;
    assign _2524 = _285 ? _2523 : _2518;
    assign _67 = _2524;
    always @(posedge _277) begin
        if (_275)
            _911 <= _1099;
        else
            _911 <= _67;
    end
    assign _2538 = 8'b11000011;
    assign _2539 = _280 == _2538;
    assign _2542 = _2539 ? _6252 : _1099;
    assign _2532 = _1386 == _2538;
    assign _2533 = _1376 & _2532;
    assign _2534 = _2533 ? _1391 : _908;
    assign _2529 = _1381 == _2538;
    assign _2530 = _1376 & _2529;
    assign _2535 = _2530 ? _1394 : _2534;
    assign _2526 = _299 == _2538;
    assign _2527 = _1376 & _2526;
    assign _2537 = _2527 ? _1099 : _2535;
    assign _2543 = _285 ? _2542 : _2537;
    assign _68 = _2543;
    always @(posedge _277) begin
        if (_275)
            _908 <= _1099;
        else
            _908 <= _68;
    end
    assign _2557 = 8'b11000010;
    assign _2558 = _280 == _2557;
    assign _2561 = _2558 ? _6252 : _1099;
    assign _2551 = _1386 == _2557;
    assign _2552 = _1376 & _2551;
    assign _2553 = _2552 ? _1391 : _905;
    assign _2548 = _1381 == _2557;
    assign _2549 = _1376 & _2548;
    assign _2554 = _2549 ? _1394 : _2553;
    assign _2545 = _299 == _2557;
    assign _2546 = _1376 & _2545;
    assign _2556 = _2546 ? _1099 : _2554;
    assign _2562 = _285 ? _2561 : _2556;
    assign _69 = _2562;
    always @(posedge _277) begin
        if (_275)
            _905 <= _1099;
        else
            _905 <= _69;
    end
    assign _2576 = 8'b11000001;
    assign _2577 = _280 == _2576;
    assign _2580 = _2577 ? _6252 : _1099;
    assign _2570 = _1386 == _2576;
    assign _2571 = _1376 & _2570;
    assign _2572 = _2571 ? _1391 : _902;
    assign _2567 = _1381 == _2576;
    assign _2568 = _1376 & _2567;
    assign _2573 = _2568 ? _1394 : _2572;
    assign _2564 = _299 == _2576;
    assign _2565 = _1376 & _2564;
    assign _2575 = _2565 ? _1099 : _2573;
    assign _2581 = _285 ? _2580 : _2575;
    assign _70 = _2581;
    always @(posedge _277) begin
        if (_275)
            _902 <= _1099;
        else
            _902 <= _70;
    end
    assign _2595 = 8'b11000000;
    assign _2596 = _280 == _2595;
    assign _2599 = _2596 ? _6252 : _1099;
    assign _2589 = _1386 == _2595;
    assign _2590 = _1376 & _2589;
    assign _2591 = _2590 ? _1391 : _899;
    assign _2586 = _1381 == _2595;
    assign _2587 = _1376 & _2586;
    assign _2592 = _2587 ? _1394 : _2591;
    assign _2583 = _299 == _2595;
    assign _2584 = _1376 & _2583;
    assign _2594 = _2584 ? _1099 : _2592;
    assign _2600 = _285 ? _2599 : _2594;
    assign _71 = _2600;
    always @(posedge _277) begin
        if (_275)
            _899 <= _1099;
        else
            _899 <= _71;
    end
    assign _2614 = 8'b10111111;
    assign _2615 = _280 == _2614;
    assign _2618 = _2615 ? _6252 : _1099;
    assign _2608 = _1386 == _2614;
    assign _2609 = _1376 & _2608;
    assign _2610 = _2609 ? _1391 : _896;
    assign _2605 = _1381 == _2614;
    assign _2606 = _1376 & _2605;
    assign _2611 = _2606 ? _1394 : _2610;
    assign _2602 = _299 == _2614;
    assign _2603 = _1376 & _2602;
    assign _2613 = _2603 ? _1099 : _2611;
    assign _2619 = _285 ? _2618 : _2613;
    assign _72 = _2619;
    always @(posedge _277) begin
        if (_275)
            _896 <= _1099;
        else
            _896 <= _72;
    end
    assign _2633 = 8'b10111110;
    assign _2634 = _280 == _2633;
    assign _2637 = _2634 ? _6252 : _1099;
    assign _2627 = _1386 == _2633;
    assign _2628 = _1376 & _2627;
    assign _2629 = _2628 ? _1391 : _893;
    assign _2624 = _1381 == _2633;
    assign _2625 = _1376 & _2624;
    assign _2630 = _2625 ? _1394 : _2629;
    assign _2621 = _299 == _2633;
    assign _2622 = _1376 & _2621;
    assign _2632 = _2622 ? _1099 : _2630;
    assign _2638 = _285 ? _2637 : _2632;
    assign _73 = _2638;
    always @(posedge _277) begin
        if (_275)
            _893 <= _1099;
        else
            _893 <= _73;
    end
    assign _2652 = 8'b10111101;
    assign _2653 = _280 == _2652;
    assign _2656 = _2653 ? _6252 : _1099;
    assign _2646 = _1386 == _2652;
    assign _2647 = _1376 & _2646;
    assign _2648 = _2647 ? _1391 : _890;
    assign _2643 = _1381 == _2652;
    assign _2644 = _1376 & _2643;
    assign _2649 = _2644 ? _1394 : _2648;
    assign _2640 = _299 == _2652;
    assign _2641 = _1376 & _2640;
    assign _2651 = _2641 ? _1099 : _2649;
    assign _2657 = _285 ? _2656 : _2651;
    assign _74 = _2657;
    always @(posedge _277) begin
        if (_275)
            _890 <= _1099;
        else
            _890 <= _74;
    end
    assign _2671 = 8'b10111100;
    assign _2672 = _280 == _2671;
    assign _2675 = _2672 ? _6252 : _1099;
    assign _2665 = _1386 == _2671;
    assign _2666 = _1376 & _2665;
    assign _2667 = _2666 ? _1391 : _887;
    assign _2662 = _1381 == _2671;
    assign _2663 = _1376 & _2662;
    assign _2668 = _2663 ? _1394 : _2667;
    assign _2659 = _299 == _2671;
    assign _2660 = _1376 & _2659;
    assign _2670 = _2660 ? _1099 : _2668;
    assign _2676 = _285 ? _2675 : _2670;
    assign _75 = _2676;
    always @(posedge _277) begin
        if (_275)
            _887 <= _1099;
        else
            _887 <= _75;
    end
    assign _2690 = 8'b10111011;
    assign _2691 = _280 == _2690;
    assign _2694 = _2691 ? _6252 : _1099;
    assign _2684 = _1386 == _2690;
    assign _2685 = _1376 & _2684;
    assign _2686 = _2685 ? _1391 : _884;
    assign _2681 = _1381 == _2690;
    assign _2682 = _1376 & _2681;
    assign _2687 = _2682 ? _1394 : _2686;
    assign _2678 = _299 == _2690;
    assign _2679 = _1376 & _2678;
    assign _2689 = _2679 ? _1099 : _2687;
    assign _2695 = _285 ? _2694 : _2689;
    assign _76 = _2695;
    always @(posedge _277) begin
        if (_275)
            _884 <= _1099;
        else
            _884 <= _76;
    end
    assign _2709 = 8'b10111010;
    assign _2710 = _280 == _2709;
    assign _2713 = _2710 ? _6252 : _1099;
    assign _2703 = _1386 == _2709;
    assign _2704 = _1376 & _2703;
    assign _2705 = _2704 ? _1391 : _881;
    assign _2700 = _1381 == _2709;
    assign _2701 = _1376 & _2700;
    assign _2706 = _2701 ? _1394 : _2705;
    assign _2697 = _299 == _2709;
    assign _2698 = _1376 & _2697;
    assign _2708 = _2698 ? _1099 : _2706;
    assign _2714 = _285 ? _2713 : _2708;
    assign _77 = _2714;
    always @(posedge _277) begin
        if (_275)
            _881 <= _1099;
        else
            _881 <= _77;
    end
    assign _2728 = 8'b10111001;
    assign _2729 = _280 == _2728;
    assign _2732 = _2729 ? _6252 : _1099;
    assign _2722 = _1386 == _2728;
    assign _2723 = _1376 & _2722;
    assign _2724 = _2723 ? _1391 : _878;
    assign _2719 = _1381 == _2728;
    assign _2720 = _1376 & _2719;
    assign _2725 = _2720 ? _1394 : _2724;
    assign _2716 = _299 == _2728;
    assign _2717 = _1376 & _2716;
    assign _2727 = _2717 ? _1099 : _2725;
    assign _2733 = _285 ? _2732 : _2727;
    assign _78 = _2733;
    always @(posedge _277) begin
        if (_275)
            _878 <= _1099;
        else
            _878 <= _78;
    end
    assign _2747 = 8'b10111000;
    assign _2748 = _280 == _2747;
    assign _2751 = _2748 ? _6252 : _1099;
    assign _2741 = _1386 == _2747;
    assign _2742 = _1376 & _2741;
    assign _2743 = _2742 ? _1391 : _875;
    assign _2738 = _1381 == _2747;
    assign _2739 = _1376 & _2738;
    assign _2744 = _2739 ? _1394 : _2743;
    assign _2735 = _299 == _2747;
    assign _2736 = _1376 & _2735;
    assign _2746 = _2736 ? _1099 : _2744;
    assign _2752 = _285 ? _2751 : _2746;
    assign _79 = _2752;
    always @(posedge _277) begin
        if (_275)
            _875 <= _1099;
        else
            _875 <= _79;
    end
    assign _2766 = 8'b10110111;
    assign _2767 = _280 == _2766;
    assign _2770 = _2767 ? _6252 : _1099;
    assign _2760 = _1386 == _2766;
    assign _2761 = _1376 & _2760;
    assign _2762 = _2761 ? _1391 : _872;
    assign _2757 = _1381 == _2766;
    assign _2758 = _1376 & _2757;
    assign _2763 = _2758 ? _1394 : _2762;
    assign _2754 = _299 == _2766;
    assign _2755 = _1376 & _2754;
    assign _2765 = _2755 ? _1099 : _2763;
    assign _2771 = _285 ? _2770 : _2765;
    assign _80 = _2771;
    always @(posedge _277) begin
        if (_275)
            _872 <= _1099;
        else
            _872 <= _80;
    end
    assign _2785 = 8'b10110110;
    assign _2786 = _280 == _2785;
    assign _2789 = _2786 ? _6252 : _1099;
    assign _2779 = _1386 == _2785;
    assign _2780 = _1376 & _2779;
    assign _2781 = _2780 ? _1391 : _869;
    assign _2776 = _1381 == _2785;
    assign _2777 = _1376 & _2776;
    assign _2782 = _2777 ? _1394 : _2781;
    assign _2773 = _299 == _2785;
    assign _2774 = _1376 & _2773;
    assign _2784 = _2774 ? _1099 : _2782;
    assign _2790 = _285 ? _2789 : _2784;
    assign _81 = _2790;
    always @(posedge _277) begin
        if (_275)
            _869 <= _1099;
        else
            _869 <= _81;
    end
    assign _2804 = 8'b10110101;
    assign _2805 = _280 == _2804;
    assign _2808 = _2805 ? _6252 : _1099;
    assign _2798 = _1386 == _2804;
    assign _2799 = _1376 & _2798;
    assign _2800 = _2799 ? _1391 : _866;
    assign _2795 = _1381 == _2804;
    assign _2796 = _1376 & _2795;
    assign _2801 = _2796 ? _1394 : _2800;
    assign _2792 = _299 == _2804;
    assign _2793 = _1376 & _2792;
    assign _2803 = _2793 ? _1099 : _2801;
    assign _2809 = _285 ? _2808 : _2803;
    assign _82 = _2809;
    always @(posedge _277) begin
        if (_275)
            _866 <= _1099;
        else
            _866 <= _82;
    end
    assign _2823 = 8'b10110100;
    assign _2824 = _280 == _2823;
    assign _2827 = _2824 ? _6252 : _1099;
    assign _2817 = _1386 == _2823;
    assign _2818 = _1376 & _2817;
    assign _2819 = _2818 ? _1391 : _863;
    assign _2814 = _1381 == _2823;
    assign _2815 = _1376 & _2814;
    assign _2820 = _2815 ? _1394 : _2819;
    assign _2811 = _299 == _2823;
    assign _2812 = _1376 & _2811;
    assign _2822 = _2812 ? _1099 : _2820;
    assign _2828 = _285 ? _2827 : _2822;
    assign _83 = _2828;
    always @(posedge _277) begin
        if (_275)
            _863 <= _1099;
        else
            _863 <= _83;
    end
    assign _2842 = 8'b10110011;
    assign _2843 = _280 == _2842;
    assign _2846 = _2843 ? _6252 : _1099;
    assign _2836 = _1386 == _2842;
    assign _2837 = _1376 & _2836;
    assign _2838 = _2837 ? _1391 : _860;
    assign _2833 = _1381 == _2842;
    assign _2834 = _1376 & _2833;
    assign _2839 = _2834 ? _1394 : _2838;
    assign _2830 = _299 == _2842;
    assign _2831 = _1376 & _2830;
    assign _2841 = _2831 ? _1099 : _2839;
    assign _2847 = _285 ? _2846 : _2841;
    assign _84 = _2847;
    always @(posedge _277) begin
        if (_275)
            _860 <= _1099;
        else
            _860 <= _84;
    end
    assign _2861 = 8'b10110010;
    assign _2862 = _280 == _2861;
    assign _2865 = _2862 ? _6252 : _1099;
    assign _2855 = _1386 == _2861;
    assign _2856 = _1376 & _2855;
    assign _2857 = _2856 ? _1391 : _857;
    assign _2852 = _1381 == _2861;
    assign _2853 = _1376 & _2852;
    assign _2858 = _2853 ? _1394 : _2857;
    assign _2849 = _299 == _2861;
    assign _2850 = _1376 & _2849;
    assign _2860 = _2850 ? _1099 : _2858;
    assign _2866 = _285 ? _2865 : _2860;
    assign _85 = _2866;
    always @(posedge _277) begin
        if (_275)
            _857 <= _1099;
        else
            _857 <= _85;
    end
    assign _2880 = 8'b10110001;
    assign _2881 = _280 == _2880;
    assign _2884 = _2881 ? _6252 : _1099;
    assign _2874 = _1386 == _2880;
    assign _2875 = _1376 & _2874;
    assign _2876 = _2875 ? _1391 : _854;
    assign _2871 = _1381 == _2880;
    assign _2872 = _1376 & _2871;
    assign _2877 = _2872 ? _1394 : _2876;
    assign _2868 = _299 == _2880;
    assign _2869 = _1376 & _2868;
    assign _2879 = _2869 ? _1099 : _2877;
    assign _2885 = _285 ? _2884 : _2879;
    assign _86 = _2885;
    always @(posedge _277) begin
        if (_275)
            _854 <= _1099;
        else
            _854 <= _86;
    end
    assign _2899 = 8'b10110000;
    assign _2900 = _280 == _2899;
    assign _2903 = _2900 ? _6252 : _1099;
    assign _2893 = _1386 == _2899;
    assign _2894 = _1376 & _2893;
    assign _2895 = _2894 ? _1391 : _851;
    assign _2890 = _1381 == _2899;
    assign _2891 = _1376 & _2890;
    assign _2896 = _2891 ? _1394 : _2895;
    assign _2887 = _299 == _2899;
    assign _2888 = _1376 & _2887;
    assign _2898 = _2888 ? _1099 : _2896;
    assign _2904 = _285 ? _2903 : _2898;
    assign _87 = _2904;
    always @(posedge _277) begin
        if (_275)
            _851 <= _1099;
        else
            _851 <= _87;
    end
    assign _2918 = 8'b10101111;
    assign _2919 = _280 == _2918;
    assign _2922 = _2919 ? _6252 : _1099;
    assign _2912 = _1386 == _2918;
    assign _2913 = _1376 & _2912;
    assign _2914 = _2913 ? _1391 : _848;
    assign _2909 = _1381 == _2918;
    assign _2910 = _1376 & _2909;
    assign _2915 = _2910 ? _1394 : _2914;
    assign _2906 = _299 == _2918;
    assign _2907 = _1376 & _2906;
    assign _2917 = _2907 ? _1099 : _2915;
    assign _2923 = _285 ? _2922 : _2917;
    assign _88 = _2923;
    always @(posedge _277) begin
        if (_275)
            _848 <= _1099;
        else
            _848 <= _88;
    end
    assign _2937 = 8'b10101110;
    assign _2938 = _280 == _2937;
    assign _2941 = _2938 ? _6252 : _1099;
    assign _2931 = _1386 == _2937;
    assign _2932 = _1376 & _2931;
    assign _2933 = _2932 ? _1391 : _845;
    assign _2928 = _1381 == _2937;
    assign _2929 = _1376 & _2928;
    assign _2934 = _2929 ? _1394 : _2933;
    assign _2925 = _299 == _2937;
    assign _2926 = _1376 & _2925;
    assign _2936 = _2926 ? _1099 : _2934;
    assign _2942 = _285 ? _2941 : _2936;
    assign _89 = _2942;
    always @(posedge _277) begin
        if (_275)
            _845 <= _1099;
        else
            _845 <= _89;
    end
    assign _2956 = 8'b10101101;
    assign _2957 = _280 == _2956;
    assign _2960 = _2957 ? _6252 : _1099;
    assign _2950 = _1386 == _2956;
    assign _2951 = _1376 & _2950;
    assign _2952 = _2951 ? _1391 : _842;
    assign _2947 = _1381 == _2956;
    assign _2948 = _1376 & _2947;
    assign _2953 = _2948 ? _1394 : _2952;
    assign _2944 = _299 == _2956;
    assign _2945 = _1376 & _2944;
    assign _2955 = _2945 ? _1099 : _2953;
    assign _2961 = _285 ? _2960 : _2955;
    assign _90 = _2961;
    always @(posedge _277) begin
        if (_275)
            _842 <= _1099;
        else
            _842 <= _90;
    end
    assign _2975 = 8'b10101100;
    assign _2976 = _280 == _2975;
    assign _2979 = _2976 ? _6252 : _1099;
    assign _2969 = _1386 == _2975;
    assign _2970 = _1376 & _2969;
    assign _2971 = _2970 ? _1391 : _839;
    assign _2966 = _1381 == _2975;
    assign _2967 = _1376 & _2966;
    assign _2972 = _2967 ? _1394 : _2971;
    assign _2963 = _299 == _2975;
    assign _2964 = _1376 & _2963;
    assign _2974 = _2964 ? _1099 : _2972;
    assign _2980 = _285 ? _2979 : _2974;
    assign _91 = _2980;
    always @(posedge _277) begin
        if (_275)
            _839 <= _1099;
        else
            _839 <= _91;
    end
    assign _2994 = 8'b10101011;
    assign _2995 = _280 == _2994;
    assign _2998 = _2995 ? _6252 : _1099;
    assign _2988 = _1386 == _2994;
    assign _2989 = _1376 & _2988;
    assign _2990 = _2989 ? _1391 : _836;
    assign _2985 = _1381 == _2994;
    assign _2986 = _1376 & _2985;
    assign _2991 = _2986 ? _1394 : _2990;
    assign _2982 = _299 == _2994;
    assign _2983 = _1376 & _2982;
    assign _2993 = _2983 ? _1099 : _2991;
    assign _2999 = _285 ? _2998 : _2993;
    assign _92 = _2999;
    always @(posedge _277) begin
        if (_275)
            _836 <= _1099;
        else
            _836 <= _92;
    end
    assign _3013 = 8'b10101010;
    assign _3014 = _280 == _3013;
    assign _3017 = _3014 ? _6252 : _1099;
    assign _3007 = _1386 == _3013;
    assign _3008 = _1376 & _3007;
    assign _3009 = _3008 ? _1391 : _833;
    assign _3004 = _1381 == _3013;
    assign _3005 = _1376 & _3004;
    assign _3010 = _3005 ? _1394 : _3009;
    assign _3001 = _299 == _3013;
    assign _3002 = _1376 & _3001;
    assign _3012 = _3002 ? _1099 : _3010;
    assign _3018 = _285 ? _3017 : _3012;
    assign _93 = _3018;
    always @(posedge _277) begin
        if (_275)
            _833 <= _1099;
        else
            _833 <= _93;
    end
    assign _3032 = 8'b10101001;
    assign _3033 = _280 == _3032;
    assign _3036 = _3033 ? _6252 : _1099;
    assign _3026 = _1386 == _3032;
    assign _3027 = _1376 & _3026;
    assign _3028 = _3027 ? _1391 : _830;
    assign _3023 = _1381 == _3032;
    assign _3024 = _1376 & _3023;
    assign _3029 = _3024 ? _1394 : _3028;
    assign _3020 = _299 == _3032;
    assign _3021 = _1376 & _3020;
    assign _3031 = _3021 ? _1099 : _3029;
    assign _3037 = _285 ? _3036 : _3031;
    assign _94 = _3037;
    always @(posedge _277) begin
        if (_275)
            _830 <= _1099;
        else
            _830 <= _94;
    end
    assign _3051 = 8'b10101000;
    assign _3052 = _280 == _3051;
    assign _3055 = _3052 ? _6252 : _1099;
    assign _3045 = _1386 == _3051;
    assign _3046 = _1376 & _3045;
    assign _3047 = _3046 ? _1391 : _827;
    assign _3042 = _1381 == _3051;
    assign _3043 = _1376 & _3042;
    assign _3048 = _3043 ? _1394 : _3047;
    assign _3039 = _299 == _3051;
    assign _3040 = _1376 & _3039;
    assign _3050 = _3040 ? _1099 : _3048;
    assign _3056 = _285 ? _3055 : _3050;
    assign _95 = _3056;
    always @(posedge _277) begin
        if (_275)
            _827 <= _1099;
        else
            _827 <= _95;
    end
    assign _3070 = 8'b10100111;
    assign _3071 = _280 == _3070;
    assign _3074 = _3071 ? _6252 : _1099;
    assign _3064 = _1386 == _3070;
    assign _3065 = _1376 & _3064;
    assign _3066 = _3065 ? _1391 : _824;
    assign _3061 = _1381 == _3070;
    assign _3062 = _1376 & _3061;
    assign _3067 = _3062 ? _1394 : _3066;
    assign _3058 = _299 == _3070;
    assign _3059 = _1376 & _3058;
    assign _3069 = _3059 ? _1099 : _3067;
    assign _3075 = _285 ? _3074 : _3069;
    assign _96 = _3075;
    always @(posedge _277) begin
        if (_275)
            _824 <= _1099;
        else
            _824 <= _96;
    end
    assign _3089 = 8'b10100110;
    assign _3090 = _280 == _3089;
    assign _3093 = _3090 ? _6252 : _1099;
    assign _3083 = _1386 == _3089;
    assign _3084 = _1376 & _3083;
    assign _3085 = _3084 ? _1391 : _821;
    assign _3080 = _1381 == _3089;
    assign _3081 = _1376 & _3080;
    assign _3086 = _3081 ? _1394 : _3085;
    assign _3077 = _299 == _3089;
    assign _3078 = _1376 & _3077;
    assign _3088 = _3078 ? _1099 : _3086;
    assign _3094 = _285 ? _3093 : _3088;
    assign _97 = _3094;
    always @(posedge _277) begin
        if (_275)
            _821 <= _1099;
        else
            _821 <= _97;
    end
    assign _3108 = 8'b10100101;
    assign _3109 = _280 == _3108;
    assign _3112 = _3109 ? _6252 : _1099;
    assign _3102 = _1386 == _3108;
    assign _3103 = _1376 & _3102;
    assign _3104 = _3103 ? _1391 : _818;
    assign _3099 = _1381 == _3108;
    assign _3100 = _1376 & _3099;
    assign _3105 = _3100 ? _1394 : _3104;
    assign _3096 = _299 == _3108;
    assign _3097 = _1376 & _3096;
    assign _3107 = _3097 ? _1099 : _3105;
    assign _3113 = _285 ? _3112 : _3107;
    assign _98 = _3113;
    always @(posedge _277) begin
        if (_275)
            _818 <= _1099;
        else
            _818 <= _98;
    end
    assign _3127 = 8'b10100100;
    assign _3128 = _280 == _3127;
    assign _3131 = _3128 ? _6252 : _1099;
    assign _3121 = _1386 == _3127;
    assign _3122 = _1376 & _3121;
    assign _3123 = _3122 ? _1391 : _815;
    assign _3118 = _1381 == _3127;
    assign _3119 = _1376 & _3118;
    assign _3124 = _3119 ? _1394 : _3123;
    assign _3115 = _299 == _3127;
    assign _3116 = _1376 & _3115;
    assign _3126 = _3116 ? _1099 : _3124;
    assign _3132 = _285 ? _3131 : _3126;
    assign _99 = _3132;
    always @(posedge _277) begin
        if (_275)
            _815 <= _1099;
        else
            _815 <= _99;
    end
    assign _3146 = 8'b10100011;
    assign _3147 = _280 == _3146;
    assign _3150 = _3147 ? _6252 : _1099;
    assign _3140 = _1386 == _3146;
    assign _3141 = _1376 & _3140;
    assign _3142 = _3141 ? _1391 : _812;
    assign _3137 = _1381 == _3146;
    assign _3138 = _1376 & _3137;
    assign _3143 = _3138 ? _1394 : _3142;
    assign _3134 = _299 == _3146;
    assign _3135 = _1376 & _3134;
    assign _3145 = _3135 ? _1099 : _3143;
    assign _3151 = _285 ? _3150 : _3145;
    assign _100 = _3151;
    always @(posedge _277) begin
        if (_275)
            _812 <= _1099;
        else
            _812 <= _100;
    end
    assign _3165 = 8'b10100010;
    assign _3166 = _280 == _3165;
    assign _3169 = _3166 ? _6252 : _1099;
    assign _3159 = _1386 == _3165;
    assign _3160 = _1376 & _3159;
    assign _3161 = _3160 ? _1391 : _809;
    assign _3156 = _1381 == _3165;
    assign _3157 = _1376 & _3156;
    assign _3162 = _3157 ? _1394 : _3161;
    assign _3153 = _299 == _3165;
    assign _3154 = _1376 & _3153;
    assign _3164 = _3154 ? _1099 : _3162;
    assign _3170 = _285 ? _3169 : _3164;
    assign _101 = _3170;
    always @(posedge _277) begin
        if (_275)
            _809 <= _1099;
        else
            _809 <= _101;
    end
    assign _3184 = 8'b10100001;
    assign _3185 = _280 == _3184;
    assign _3188 = _3185 ? _6252 : _1099;
    assign _3178 = _1386 == _3184;
    assign _3179 = _1376 & _3178;
    assign _3180 = _3179 ? _1391 : _806;
    assign _3175 = _1381 == _3184;
    assign _3176 = _1376 & _3175;
    assign _3181 = _3176 ? _1394 : _3180;
    assign _3172 = _299 == _3184;
    assign _3173 = _1376 & _3172;
    assign _3183 = _3173 ? _1099 : _3181;
    assign _3189 = _285 ? _3188 : _3183;
    assign _102 = _3189;
    always @(posedge _277) begin
        if (_275)
            _806 <= _1099;
        else
            _806 <= _102;
    end
    assign _3203 = 8'b10100000;
    assign _3204 = _280 == _3203;
    assign _3207 = _3204 ? _6252 : _1099;
    assign _3197 = _1386 == _3203;
    assign _3198 = _1376 & _3197;
    assign _3199 = _3198 ? _1391 : _803;
    assign _3194 = _1381 == _3203;
    assign _3195 = _1376 & _3194;
    assign _3200 = _3195 ? _1394 : _3199;
    assign _3191 = _299 == _3203;
    assign _3192 = _1376 & _3191;
    assign _3202 = _3192 ? _1099 : _3200;
    assign _3208 = _285 ? _3207 : _3202;
    assign _103 = _3208;
    always @(posedge _277) begin
        if (_275)
            _803 <= _1099;
        else
            _803 <= _103;
    end
    assign _3222 = 8'b10011111;
    assign _3223 = _280 == _3222;
    assign _3226 = _3223 ? _6252 : _1099;
    assign _3216 = _1386 == _3222;
    assign _3217 = _1376 & _3216;
    assign _3218 = _3217 ? _1391 : _800;
    assign _3213 = _1381 == _3222;
    assign _3214 = _1376 & _3213;
    assign _3219 = _3214 ? _1394 : _3218;
    assign _3210 = _299 == _3222;
    assign _3211 = _1376 & _3210;
    assign _3221 = _3211 ? _1099 : _3219;
    assign _3227 = _285 ? _3226 : _3221;
    assign _104 = _3227;
    always @(posedge _277) begin
        if (_275)
            _800 <= _1099;
        else
            _800 <= _104;
    end
    assign _3241 = 8'b10011110;
    assign _3242 = _280 == _3241;
    assign _3245 = _3242 ? _6252 : _1099;
    assign _3235 = _1386 == _3241;
    assign _3236 = _1376 & _3235;
    assign _3237 = _3236 ? _1391 : _797;
    assign _3232 = _1381 == _3241;
    assign _3233 = _1376 & _3232;
    assign _3238 = _3233 ? _1394 : _3237;
    assign _3229 = _299 == _3241;
    assign _3230 = _1376 & _3229;
    assign _3240 = _3230 ? _1099 : _3238;
    assign _3246 = _285 ? _3245 : _3240;
    assign _105 = _3246;
    always @(posedge _277) begin
        if (_275)
            _797 <= _1099;
        else
            _797 <= _105;
    end
    assign _3260 = 8'b10011101;
    assign _3261 = _280 == _3260;
    assign _3264 = _3261 ? _6252 : _1099;
    assign _3254 = _1386 == _3260;
    assign _3255 = _1376 & _3254;
    assign _3256 = _3255 ? _1391 : _794;
    assign _3251 = _1381 == _3260;
    assign _3252 = _1376 & _3251;
    assign _3257 = _3252 ? _1394 : _3256;
    assign _3248 = _299 == _3260;
    assign _3249 = _1376 & _3248;
    assign _3259 = _3249 ? _1099 : _3257;
    assign _3265 = _285 ? _3264 : _3259;
    assign _106 = _3265;
    always @(posedge _277) begin
        if (_275)
            _794 <= _1099;
        else
            _794 <= _106;
    end
    assign _3279 = 8'b10011100;
    assign _3280 = _280 == _3279;
    assign _3283 = _3280 ? _6252 : _1099;
    assign _3273 = _1386 == _3279;
    assign _3274 = _1376 & _3273;
    assign _3275 = _3274 ? _1391 : _791;
    assign _3270 = _1381 == _3279;
    assign _3271 = _1376 & _3270;
    assign _3276 = _3271 ? _1394 : _3275;
    assign _3267 = _299 == _3279;
    assign _3268 = _1376 & _3267;
    assign _3278 = _3268 ? _1099 : _3276;
    assign _3284 = _285 ? _3283 : _3278;
    assign _107 = _3284;
    always @(posedge _277) begin
        if (_275)
            _791 <= _1099;
        else
            _791 <= _107;
    end
    assign _3298 = 8'b10011011;
    assign _3299 = _280 == _3298;
    assign _3302 = _3299 ? _6252 : _1099;
    assign _3292 = _1386 == _3298;
    assign _3293 = _1376 & _3292;
    assign _3294 = _3293 ? _1391 : _788;
    assign _3289 = _1381 == _3298;
    assign _3290 = _1376 & _3289;
    assign _3295 = _3290 ? _1394 : _3294;
    assign _3286 = _299 == _3298;
    assign _3287 = _1376 & _3286;
    assign _3297 = _3287 ? _1099 : _3295;
    assign _3303 = _285 ? _3302 : _3297;
    assign _108 = _3303;
    always @(posedge _277) begin
        if (_275)
            _788 <= _1099;
        else
            _788 <= _108;
    end
    assign _3317 = 8'b10011010;
    assign _3318 = _280 == _3317;
    assign _3321 = _3318 ? _6252 : _1099;
    assign _3311 = _1386 == _3317;
    assign _3312 = _1376 & _3311;
    assign _3313 = _3312 ? _1391 : _785;
    assign _3308 = _1381 == _3317;
    assign _3309 = _1376 & _3308;
    assign _3314 = _3309 ? _1394 : _3313;
    assign _3305 = _299 == _3317;
    assign _3306 = _1376 & _3305;
    assign _3316 = _3306 ? _1099 : _3314;
    assign _3322 = _285 ? _3321 : _3316;
    assign _109 = _3322;
    always @(posedge _277) begin
        if (_275)
            _785 <= _1099;
        else
            _785 <= _109;
    end
    assign _3336 = 8'b10011001;
    assign _3337 = _280 == _3336;
    assign _3340 = _3337 ? _6252 : _1099;
    assign _3330 = _1386 == _3336;
    assign _3331 = _1376 & _3330;
    assign _3332 = _3331 ? _1391 : _782;
    assign _3327 = _1381 == _3336;
    assign _3328 = _1376 & _3327;
    assign _3333 = _3328 ? _1394 : _3332;
    assign _3324 = _299 == _3336;
    assign _3325 = _1376 & _3324;
    assign _3335 = _3325 ? _1099 : _3333;
    assign _3341 = _285 ? _3340 : _3335;
    assign _110 = _3341;
    always @(posedge _277) begin
        if (_275)
            _782 <= _1099;
        else
            _782 <= _110;
    end
    assign _3355 = 8'b10011000;
    assign _3356 = _280 == _3355;
    assign _3359 = _3356 ? _6252 : _1099;
    assign _3349 = _1386 == _3355;
    assign _3350 = _1376 & _3349;
    assign _3351 = _3350 ? _1391 : _779;
    assign _3346 = _1381 == _3355;
    assign _3347 = _1376 & _3346;
    assign _3352 = _3347 ? _1394 : _3351;
    assign _3343 = _299 == _3355;
    assign _3344 = _1376 & _3343;
    assign _3354 = _3344 ? _1099 : _3352;
    assign _3360 = _285 ? _3359 : _3354;
    assign _111 = _3360;
    always @(posedge _277) begin
        if (_275)
            _779 <= _1099;
        else
            _779 <= _111;
    end
    assign _3374 = 8'b10010111;
    assign _3375 = _280 == _3374;
    assign _3378 = _3375 ? _6252 : _1099;
    assign _3368 = _1386 == _3374;
    assign _3369 = _1376 & _3368;
    assign _3370 = _3369 ? _1391 : _776;
    assign _3365 = _1381 == _3374;
    assign _3366 = _1376 & _3365;
    assign _3371 = _3366 ? _1394 : _3370;
    assign _3362 = _299 == _3374;
    assign _3363 = _1376 & _3362;
    assign _3373 = _3363 ? _1099 : _3371;
    assign _3379 = _285 ? _3378 : _3373;
    assign _112 = _3379;
    always @(posedge _277) begin
        if (_275)
            _776 <= _1099;
        else
            _776 <= _112;
    end
    assign _3393 = 8'b10010110;
    assign _3394 = _280 == _3393;
    assign _3397 = _3394 ? _6252 : _1099;
    assign _3387 = _1386 == _3393;
    assign _3388 = _1376 & _3387;
    assign _3389 = _3388 ? _1391 : _773;
    assign _3384 = _1381 == _3393;
    assign _3385 = _1376 & _3384;
    assign _3390 = _3385 ? _1394 : _3389;
    assign _3381 = _299 == _3393;
    assign _3382 = _1376 & _3381;
    assign _3392 = _3382 ? _1099 : _3390;
    assign _3398 = _285 ? _3397 : _3392;
    assign _113 = _3398;
    always @(posedge _277) begin
        if (_275)
            _773 <= _1099;
        else
            _773 <= _113;
    end
    assign _3412 = 8'b10010101;
    assign _3413 = _280 == _3412;
    assign _3416 = _3413 ? _6252 : _1099;
    assign _3406 = _1386 == _3412;
    assign _3407 = _1376 & _3406;
    assign _3408 = _3407 ? _1391 : _770;
    assign _3403 = _1381 == _3412;
    assign _3404 = _1376 & _3403;
    assign _3409 = _3404 ? _1394 : _3408;
    assign _3400 = _299 == _3412;
    assign _3401 = _1376 & _3400;
    assign _3411 = _3401 ? _1099 : _3409;
    assign _3417 = _285 ? _3416 : _3411;
    assign _114 = _3417;
    always @(posedge _277) begin
        if (_275)
            _770 <= _1099;
        else
            _770 <= _114;
    end
    assign _3431 = 8'b10010100;
    assign _3432 = _280 == _3431;
    assign _3435 = _3432 ? _6252 : _1099;
    assign _3425 = _1386 == _3431;
    assign _3426 = _1376 & _3425;
    assign _3427 = _3426 ? _1391 : _767;
    assign _3422 = _1381 == _3431;
    assign _3423 = _1376 & _3422;
    assign _3428 = _3423 ? _1394 : _3427;
    assign _3419 = _299 == _3431;
    assign _3420 = _1376 & _3419;
    assign _3430 = _3420 ? _1099 : _3428;
    assign _3436 = _285 ? _3435 : _3430;
    assign _115 = _3436;
    always @(posedge _277) begin
        if (_275)
            _767 <= _1099;
        else
            _767 <= _115;
    end
    assign _3450 = 8'b10010011;
    assign _3451 = _280 == _3450;
    assign _3454 = _3451 ? _6252 : _1099;
    assign _3444 = _1386 == _3450;
    assign _3445 = _1376 & _3444;
    assign _3446 = _3445 ? _1391 : _764;
    assign _3441 = _1381 == _3450;
    assign _3442 = _1376 & _3441;
    assign _3447 = _3442 ? _1394 : _3446;
    assign _3438 = _299 == _3450;
    assign _3439 = _1376 & _3438;
    assign _3449 = _3439 ? _1099 : _3447;
    assign _3455 = _285 ? _3454 : _3449;
    assign _116 = _3455;
    always @(posedge _277) begin
        if (_275)
            _764 <= _1099;
        else
            _764 <= _116;
    end
    assign _3469 = 8'b10010010;
    assign _3470 = _280 == _3469;
    assign _3473 = _3470 ? _6252 : _1099;
    assign _3463 = _1386 == _3469;
    assign _3464 = _1376 & _3463;
    assign _3465 = _3464 ? _1391 : _761;
    assign _3460 = _1381 == _3469;
    assign _3461 = _1376 & _3460;
    assign _3466 = _3461 ? _1394 : _3465;
    assign _3457 = _299 == _3469;
    assign _3458 = _1376 & _3457;
    assign _3468 = _3458 ? _1099 : _3466;
    assign _3474 = _285 ? _3473 : _3468;
    assign _117 = _3474;
    always @(posedge _277) begin
        if (_275)
            _761 <= _1099;
        else
            _761 <= _117;
    end
    assign _3488 = 8'b10010001;
    assign _3489 = _280 == _3488;
    assign _3492 = _3489 ? _6252 : _1099;
    assign _3482 = _1386 == _3488;
    assign _3483 = _1376 & _3482;
    assign _3484 = _3483 ? _1391 : _758;
    assign _3479 = _1381 == _3488;
    assign _3480 = _1376 & _3479;
    assign _3485 = _3480 ? _1394 : _3484;
    assign _3476 = _299 == _3488;
    assign _3477 = _1376 & _3476;
    assign _3487 = _3477 ? _1099 : _3485;
    assign _3493 = _285 ? _3492 : _3487;
    assign _118 = _3493;
    always @(posedge _277) begin
        if (_275)
            _758 <= _1099;
        else
            _758 <= _118;
    end
    assign _3507 = 8'b10010000;
    assign _3508 = _280 == _3507;
    assign _3511 = _3508 ? _6252 : _1099;
    assign _3501 = _1386 == _3507;
    assign _3502 = _1376 & _3501;
    assign _3503 = _3502 ? _1391 : _755;
    assign _3498 = _1381 == _3507;
    assign _3499 = _1376 & _3498;
    assign _3504 = _3499 ? _1394 : _3503;
    assign _3495 = _299 == _3507;
    assign _3496 = _1376 & _3495;
    assign _3506 = _3496 ? _1099 : _3504;
    assign _3512 = _285 ? _3511 : _3506;
    assign _119 = _3512;
    always @(posedge _277) begin
        if (_275)
            _755 <= _1099;
        else
            _755 <= _119;
    end
    assign _3526 = 8'b10001111;
    assign _3527 = _280 == _3526;
    assign _3530 = _3527 ? _6252 : _1099;
    assign _3520 = _1386 == _3526;
    assign _3521 = _1376 & _3520;
    assign _3522 = _3521 ? _1391 : _752;
    assign _3517 = _1381 == _3526;
    assign _3518 = _1376 & _3517;
    assign _3523 = _3518 ? _1394 : _3522;
    assign _3514 = _299 == _3526;
    assign _3515 = _1376 & _3514;
    assign _3525 = _3515 ? _1099 : _3523;
    assign _3531 = _285 ? _3530 : _3525;
    assign _120 = _3531;
    always @(posedge _277) begin
        if (_275)
            _752 <= _1099;
        else
            _752 <= _120;
    end
    assign _3545 = 8'b10001110;
    assign _3546 = _280 == _3545;
    assign _3549 = _3546 ? _6252 : _1099;
    assign _3539 = _1386 == _3545;
    assign _3540 = _1376 & _3539;
    assign _3541 = _3540 ? _1391 : _749;
    assign _3536 = _1381 == _3545;
    assign _3537 = _1376 & _3536;
    assign _3542 = _3537 ? _1394 : _3541;
    assign _3533 = _299 == _3545;
    assign _3534 = _1376 & _3533;
    assign _3544 = _3534 ? _1099 : _3542;
    assign _3550 = _285 ? _3549 : _3544;
    assign _121 = _3550;
    always @(posedge _277) begin
        if (_275)
            _749 <= _1099;
        else
            _749 <= _121;
    end
    assign _3564 = 8'b10001101;
    assign _3565 = _280 == _3564;
    assign _3568 = _3565 ? _6252 : _1099;
    assign _3558 = _1386 == _3564;
    assign _3559 = _1376 & _3558;
    assign _3560 = _3559 ? _1391 : _746;
    assign _3555 = _1381 == _3564;
    assign _3556 = _1376 & _3555;
    assign _3561 = _3556 ? _1394 : _3560;
    assign _3552 = _299 == _3564;
    assign _3553 = _1376 & _3552;
    assign _3563 = _3553 ? _1099 : _3561;
    assign _3569 = _285 ? _3568 : _3563;
    assign _122 = _3569;
    always @(posedge _277) begin
        if (_275)
            _746 <= _1099;
        else
            _746 <= _122;
    end
    assign _3583 = 8'b10001100;
    assign _3584 = _280 == _3583;
    assign _3587 = _3584 ? _6252 : _1099;
    assign _3577 = _1386 == _3583;
    assign _3578 = _1376 & _3577;
    assign _3579 = _3578 ? _1391 : _743;
    assign _3574 = _1381 == _3583;
    assign _3575 = _1376 & _3574;
    assign _3580 = _3575 ? _1394 : _3579;
    assign _3571 = _299 == _3583;
    assign _3572 = _1376 & _3571;
    assign _3582 = _3572 ? _1099 : _3580;
    assign _3588 = _285 ? _3587 : _3582;
    assign _123 = _3588;
    always @(posedge _277) begin
        if (_275)
            _743 <= _1099;
        else
            _743 <= _123;
    end
    assign _3602 = 8'b10001011;
    assign _3603 = _280 == _3602;
    assign _3606 = _3603 ? _6252 : _1099;
    assign _3596 = _1386 == _3602;
    assign _3597 = _1376 & _3596;
    assign _3598 = _3597 ? _1391 : _740;
    assign _3593 = _1381 == _3602;
    assign _3594 = _1376 & _3593;
    assign _3599 = _3594 ? _1394 : _3598;
    assign _3590 = _299 == _3602;
    assign _3591 = _1376 & _3590;
    assign _3601 = _3591 ? _1099 : _3599;
    assign _3607 = _285 ? _3606 : _3601;
    assign _124 = _3607;
    always @(posedge _277) begin
        if (_275)
            _740 <= _1099;
        else
            _740 <= _124;
    end
    assign _3621 = 8'b10001010;
    assign _3622 = _280 == _3621;
    assign _3625 = _3622 ? _6252 : _1099;
    assign _3615 = _1386 == _3621;
    assign _3616 = _1376 & _3615;
    assign _3617 = _3616 ? _1391 : _737;
    assign _3612 = _1381 == _3621;
    assign _3613 = _1376 & _3612;
    assign _3618 = _3613 ? _1394 : _3617;
    assign _3609 = _299 == _3621;
    assign _3610 = _1376 & _3609;
    assign _3620 = _3610 ? _1099 : _3618;
    assign _3626 = _285 ? _3625 : _3620;
    assign _125 = _3626;
    always @(posedge _277) begin
        if (_275)
            _737 <= _1099;
        else
            _737 <= _125;
    end
    assign _3640 = 8'b10001001;
    assign _3641 = _280 == _3640;
    assign _3644 = _3641 ? _6252 : _1099;
    assign _3634 = _1386 == _3640;
    assign _3635 = _1376 & _3634;
    assign _3636 = _3635 ? _1391 : _734;
    assign _3631 = _1381 == _3640;
    assign _3632 = _1376 & _3631;
    assign _3637 = _3632 ? _1394 : _3636;
    assign _3628 = _299 == _3640;
    assign _3629 = _1376 & _3628;
    assign _3639 = _3629 ? _1099 : _3637;
    assign _3645 = _285 ? _3644 : _3639;
    assign _126 = _3645;
    always @(posedge _277) begin
        if (_275)
            _734 <= _1099;
        else
            _734 <= _126;
    end
    assign _3659 = 8'b10001000;
    assign _3660 = _280 == _3659;
    assign _3663 = _3660 ? _6252 : _1099;
    assign _3653 = _1386 == _3659;
    assign _3654 = _1376 & _3653;
    assign _3655 = _3654 ? _1391 : _731;
    assign _3650 = _1381 == _3659;
    assign _3651 = _1376 & _3650;
    assign _3656 = _3651 ? _1394 : _3655;
    assign _3647 = _299 == _3659;
    assign _3648 = _1376 & _3647;
    assign _3658 = _3648 ? _1099 : _3656;
    assign _3664 = _285 ? _3663 : _3658;
    assign _127 = _3664;
    always @(posedge _277) begin
        if (_275)
            _731 <= _1099;
        else
            _731 <= _127;
    end
    assign _3678 = 8'b10000111;
    assign _3679 = _280 == _3678;
    assign _3682 = _3679 ? _6252 : _1099;
    assign _3672 = _1386 == _3678;
    assign _3673 = _1376 & _3672;
    assign _3674 = _3673 ? _1391 : _728;
    assign _3669 = _1381 == _3678;
    assign _3670 = _1376 & _3669;
    assign _3675 = _3670 ? _1394 : _3674;
    assign _3666 = _299 == _3678;
    assign _3667 = _1376 & _3666;
    assign _3677 = _3667 ? _1099 : _3675;
    assign _3683 = _285 ? _3682 : _3677;
    assign _128 = _3683;
    always @(posedge _277) begin
        if (_275)
            _728 <= _1099;
        else
            _728 <= _128;
    end
    assign _3697 = 8'b10000110;
    assign _3698 = _280 == _3697;
    assign _3701 = _3698 ? _6252 : _1099;
    assign _3691 = _1386 == _3697;
    assign _3692 = _1376 & _3691;
    assign _3693 = _3692 ? _1391 : _725;
    assign _3688 = _1381 == _3697;
    assign _3689 = _1376 & _3688;
    assign _3694 = _3689 ? _1394 : _3693;
    assign _3685 = _299 == _3697;
    assign _3686 = _1376 & _3685;
    assign _3696 = _3686 ? _1099 : _3694;
    assign _3702 = _285 ? _3701 : _3696;
    assign _129 = _3702;
    always @(posedge _277) begin
        if (_275)
            _725 <= _1099;
        else
            _725 <= _129;
    end
    assign _3716 = 8'b10000101;
    assign _3717 = _280 == _3716;
    assign _3720 = _3717 ? _6252 : _1099;
    assign _3710 = _1386 == _3716;
    assign _3711 = _1376 & _3710;
    assign _3712 = _3711 ? _1391 : _722;
    assign _3707 = _1381 == _3716;
    assign _3708 = _1376 & _3707;
    assign _3713 = _3708 ? _1394 : _3712;
    assign _3704 = _299 == _3716;
    assign _3705 = _1376 & _3704;
    assign _3715 = _3705 ? _1099 : _3713;
    assign _3721 = _285 ? _3720 : _3715;
    assign _130 = _3721;
    always @(posedge _277) begin
        if (_275)
            _722 <= _1099;
        else
            _722 <= _130;
    end
    assign _3735 = 8'b10000100;
    assign _3736 = _280 == _3735;
    assign _3739 = _3736 ? _6252 : _1099;
    assign _3729 = _1386 == _3735;
    assign _3730 = _1376 & _3729;
    assign _3731 = _3730 ? _1391 : _719;
    assign _3726 = _1381 == _3735;
    assign _3727 = _1376 & _3726;
    assign _3732 = _3727 ? _1394 : _3731;
    assign _3723 = _299 == _3735;
    assign _3724 = _1376 & _3723;
    assign _3734 = _3724 ? _1099 : _3732;
    assign _3740 = _285 ? _3739 : _3734;
    assign _131 = _3740;
    always @(posedge _277) begin
        if (_275)
            _719 <= _1099;
        else
            _719 <= _131;
    end
    assign _3754 = 8'b10000011;
    assign _3755 = _280 == _3754;
    assign _3758 = _3755 ? _6252 : _1099;
    assign _3748 = _1386 == _3754;
    assign _3749 = _1376 & _3748;
    assign _3750 = _3749 ? _1391 : _716;
    assign _3745 = _1381 == _3754;
    assign _3746 = _1376 & _3745;
    assign _3751 = _3746 ? _1394 : _3750;
    assign _3742 = _299 == _3754;
    assign _3743 = _1376 & _3742;
    assign _3753 = _3743 ? _1099 : _3751;
    assign _3759 = _285 ? _3758 : _3753;
    assign _132 = _3759;
    always @(posedge _277) begin
        if (_275)
            _716 <= _1099;
        else
            _716 <= _132;
    end
    assign _3773 = 8'b10000010;
    assign _3774 = _280 == _3773;
    assign _3777 = _3774 ? _6252 : _1099;
    assign _3767 = _1386 == _3773;
    assign _3768 = _1376 & _3767;
    assign _3769 = _3768 ? _1391 : _713;
    assign _3764 = _1381 == _3773;
    assign _3765 = _1376 & _3764;
    assign _3770 = _3765 ? _1394 : _3769;
    assign _3761 = _299 == _3773;
    assign _3762 = _1376 & _3761;
    assign _3772 = _3762 ? _1099 : _3770;
    assign _3778 = _285 ? _3777 : _3772;
    assign _133 = _3778;
    always @(posedge _277) begin
        if (_275)
            _713 <= _1099;
        else
            _713 <= _133;
    end
    assign _3792 = 8'b10000001;
    assign _3793 = _280 == _3792;
    assign _3796 = _3793 ? _6252 : _1099;
    assign _3786 = _1386 == _3792;
    assign _3787 = _1376 & _3786;
    assign _3788 = _3787 ? _1391 : _710;
    assign _3783 = _1381 == _3792;
    assign _3784 = _1376 & _3783;
    assign _3789 = _3784 ? _1394 : _3788;
    assign _3780 = _299 == _3792;
    assign _3781 = _1376 & _3780;
    assign _3791 = _3781 ? _1099 : _3789;
    assign _3797 = _285 ? _3796 : _3791;
    assign _134 = _3797;
    always @(posedge _277) begin
        if (_275)
            _710 <= _1099;
        else
            _710 <= _134;
    end
    assign _3811 = 8'b10000000;
    assign _3812 = _280 == _3811;
    assign _3815 = _3812 ? _6252 : _1099;
    assign _3805 = _1386 == _3811;
    assign _3806 = _1376 & _3805;
    assign _3807 = _3806 ? _1391 : _707;
    assign _3802 = _1381 == _3811;
    assign _3803 = _1376 & _3802;
    assign _3808 = _3803 ? _1394 : _3807;
    assign _3799 = _299 == _3811;
    assign _3800 = _1376 & _3799;
    assign _3810 = _3800 ? _1099 : _3808;
    assign _3816 = _285 ? _3815 : _3810;
    assign _135 = _3816;
    always @(posedge _277) begin
        if (_275)
            _707 <= _1099;
        else
            _707 <= _135;
    end
    assign _3830 = 8'b01111111;
    assign _3831 = _280 == _3830;
    assign _3834 = _3831 ? _6252 : _1099;
    assign _3824 = _1386 == _3830;
    assign _3825 = _1376 & _3824;
    assign _3826 = _3825 ? _1391 : _704;
    assign _3821 = _1381 == _3830;
    assign _3822 = _1376 & _3821;
    assign _3827 = _3822 ? _1394 : _3826;
    assign _3818 = _299 == _3830;
    assign _3819 = _1376 & _3818;
    assign _3829 = _3819 ? _1099 : _3827;
    assign _3835 = _285 ? _3834 : _3829;
    assign _136 = _3835;
    always @(posedge _277) begin
        if (_275)
            _704 <= _1099;
        else
            _704 <= _136;
    end
    assign _3849 = 8'b01111110;
    assign _3850 = _280 == _3849;
    assign _3853 = _3850 ? _6252 : _1099;
    assign _3843 = _1386 == _3849;
    assign _3844 = _1376 & _3843;
    assign _3845 = _3844 ? _1391 : _701;
    assign _3840 = _1381 == _3849;
    assign _3841 = _1376 & _3840;
    assign _3846 = _3841 ? _1394 : _3845;
    assign _3837 = _299 == _3849;
    assign _3838 = _1376 & _3837;
    assign _3848 = _3838 ? _1099 : _3846;
    assign _3854 = _285 ? _3853 : _3848;
    assign _137 = _3854;
    always @(posedge _277) begin
        if (_275)
            _701 <= _1099;
        else
            _701 <= _137;
    end
    assign _3868 = 8'b01111101;
    assign _3869 = _280 == _3868;
    assign _3872 = _3869 ? _6252 : _1099;
    assign _3862 = _1386 == _3868;
    assign _3863 = _1376 & _3862;
    assign _3864 = _3863 ? _1391 : _698;
    assign _3859 = _1381 == _3868;
    assign _3860 = _1376 & _3859;
    assign _3865 = _3860 ? _1394 : _3864;
    assign _3856 = _299 == _3868;
    assign _3857 = _1376 & _3856;
    assign _3867 = _3857 ? _1099 : _3865;
    assign _3873 = _285 ? _3872 : _3867;
    assign _138 = _3873;
    always @(posedge _277) begin
        if (_275)
            _698 <= _1099;
        else
            _698 <= _138;
    end
    assign _3887 = 8'b01111100;
    assign _3888 = _280 == _3887;
    assign _3891 = _3888 ? _6252 : _1099;
    assign _3881 = _1386 == _3887;
    assign _3882 = _1376 & _3881;
    assign _3883 = _3882 ? _1391 : _695;
    assign _3878 = _1381 == _3887;
    assign _3879 = _1376 & _3878;
    assign _3884 = _3879 ? _1394 : _3883;
    assign _3875 = _299 == _3887;
    assign _3876 = _1376 & _3875;
    assign _3886 = _3876 ? _1099 : _3884;
    assign _3892 = _285 ? _3891 : _3886;
    assign _139 = _3892;
    always @(posedge _277) begin
        if (_275)
            _695 <= _1099;
        else
            _695 <= _139;
    end
    assign _3906 = 8'b01111011;
    assign _3907 = _280 == _3906;
    assign _3910 = _3907 ? _6252 : _1099;
    assign _3900 = _1386 == _3906;
    assign _3901 = _1376 & _3900;
    assign _3902 = _3901 ? _1391 : _692;
    assign _3897 = _1381 == _3906;
    assign _3898 = _1376 & _3897;
    assign _3903 = _3898 ? _1394 : _3902;
    assign _3894 = _299 == _3906;
    assign _3895 = _1376 & _3894;
    assign _3905 = _3895 ? _1099 : _3903;
    assign _3911 = _285 ? _3910 : _3905;
    assign _140 = _3911;
    always @(posedge _277) begin
        if (_275)
            _692 <= _1099;
        else
            _692 <= _140;
    end
    assign _3925 = 8'b01111010;
    assign _3926 = _280 == _3925;
    assign _3929 = _3926 ? _6252 : _1099;
    assign _3919 = _1386 == _3925;
    assign _3920 = _1376 & _3919;
    assign _3921 = _3920 ? _1391 : _689;
    assign _3916 = _1381 == _3925;
    assign _3917 = _1376 & _3916;
    assign _3922 = _3917 ? _1394 : _3921;
    assign _3913 = _299 == _3925;
    assign _3914 = _1376 & _3913;
    assign _3924 = _3914 ? _1099 : _3922;
    assign _3930 = _285 ? _3929 : _3924;
    assign _141 = _3930;
    always @(posedge _277) begin
        if (_275)
            _689 <= _1099;
        else
            _689 <= _141;
    end
    assign _3944 = 8'b01111001;
    assign _3945 = _280 == _3944;
    assign _3948 = _3945 ? _6252 : _1099;
    assign _3938 = _1386 == _3944;
    assign _3939 = _1376 & _3938;
    assign _3940 = _3939 ? _1391 : _686;
    assign _3935 = _1381 == _3944;
    assign _3936 = _1376 & _3935;
    assign _3941 = _3936 ? _1394 : _3940;
    assign _3932 = _299 == _3944;
    assign _3933 = _1376 & _3932;
    assign _3943 = _3933 ? _1099 : _3941;
    assign _3949 = _285 ? _3948 : _3943;
    assign _142 = _3949;
    always @(posedge _277) begin
        if (_275)
            _686 <= _1099;
        else
            _686 <= _142;
    end
    assign _3963 = 8'b01111000;
    assign _3964 = _280 == _3963;
    assign _3967 = _3964 ? _6252 : _1099;
    assign _3957 = _1386 == _3963;
    assign _3958 = _1376 & _3957;
    assign _3959 = _3958 ? _1391 : _683;
    assign _3954 = _1381 == _3963;
    assign _3955 = _1376 & _3954;
    assign _3960 = _3955 ? _1394 : _3959;
    assign _3951 = _299 == _3963;
    assign _3952 = _1376 & _3951;
    assign _3962 = _3952 ? _1099 : _3960;
    assign _3968 = _285 ? _3967 : _3962;
    assign _143 = _3968;
    always @(posedge _277) begin
        if (_275)
            _683 <= _1099;
        else
            _683 <= _143;
    end
    assign _3982 = 8'b01110111;
    assign _3983 = _280 == _3982;
    assign _3986 = _3983 ? _6252 : _1099;
    assign _3976 = _1386 == _3982;
    assign _3977 = _1376 & _3976;
    assign _3978 = _3977 ? _1391 : _680;
    assign _3973 = _1381 == _3982;
    assign _3974 = _1376 & _3973;
    assign _3979 = _3974 ? _1394 : _3978;
    assign _3970 = _299 == _3982;
    assign _3971 = _1376 & _3970;
    assign _3981 = _3971 ? _1099 : _3979;
    assign _3987 = _285 ? _3986 : _3981;
    assign _144 = _3987;
    always @(posedge _277) begin
        if (_275)
            _680 <= _1099;
        else
            _680 <= _144;
    end
    assign _4001 = 8'b01110110;
    assign _4002 = _280 == _4001;
    assign _4005 = _4002 ? _6252 : _1099;
    assign _3995 = _1386 == _4001;
    assign _3996 = _1376 & _3995;
    assign _3997 = _3996 ? _1391 : _677;
    assign _3992 = _1381 == _4001;
    assign _3993 = _1376 & _3992;
    assign _3998 = _3993 ? _1394 : _3997;
    assign _3989 = _299 == _4001;
    assign _3990 = _1376 & _3989;
    assign _4000 = _3990 ? _1099 : _3998;
    assign _4006 = _285 ? _4005 : _4000;
    assign _145 = _4006;
    always @(posedge _277) begin
        if (_275)
            _677 <= _1099;
        else
            _677 <= _145;
    end
    assign _4020 = 8'b01110101;
    assign _4021 = _280 == _4020;
    assign _4024 = _4021 ? _6252 : _1099;
    assign _4014 = _1386 == _4020;
    assign _4015 = _1376 & _4014;
    assign _4016 = _4015 ? _1391 : _674;
    assign _4011 = _1381 == _4020;
    assign _4012 = _1376 & _4011;
    assign _4017 = _4012 ? _1394 : _4016;
    assign _4008 = _299 == _4020;
    assign _4009 = _1376 & _4008;
    assign _4019 = _4009 ? _1099 : _4017;
    assign _4025 = _285 ? _4024 : _4019;
    assign _146 = _4025;
    always @(posedge _277) begin
        if (_275)
            _674 <= _1099;
        else
            _674 <= _146;
    end
    assign _4039 = 8'b01110100;
    assign _4040 = _280 == _4039;
    assign _4043 = _4040 ? _6252 : _1099;
    assign _4033 = _1386 == _4039;
    assign _4034 = _1376 & _4033;
    assign _4035 = _4034 ? _1391 : _671;
    assign _4030 = _1381 == _4039;
    assign _4031 = _1376 & _4030;
    assign _4036 = _4031 ? _1394 : _4035;
    assign _4027 = _299 == _4039;
    assign _4028 = _1376 & _4027;
    assign _4038 = _4028 ? _1099 : _4036;
    assign _4044 = _285 ? _4043 : _4038;
    assign _147 = _4044;
    always @(posedge _277) begin
        if (_275)
            _671 <= _1099;
        else
            _671 <= _147;
    end
    assign _4058 = 8'b01110011;
    assign _4059 = _280 == _4058;
    assign _4062 = _4059 ? _6252 : _1099;
    assign _4052 = _1386 == _4058;
    assign _4053 = _1376 & _4052;
    assign _4054 = _4053 ? _1391 : _668;
    assign _4049 = _1381 == _4058;
    assign _4050 = _1376 & _4049;
    assign _4055 = _4050 ? _1394 : _4054;
    assign _4046 = _299 == _4058;
    assign _4047 = _1376 & _4046;
    assign _4057 = _4047 ? _1099 : _4055;
    assign _4063 = _285 ? _4062 : _4057;
    assign _148 = _4063;
    always @(posedge _277) begin
        if (_275)
            _668 <= _1099;
        else
            _668 <= _148;
    end
    assign _4077 = 8'b01110010;
    assign _4078 = _280 == _4077;
    assign _4081 = _4078 ? _6252 : _1099;
    assign _4071 = _1386 == _4077;
    assign _4072 = _1376 & _4071;
    assign _4073 = _4072 ? _1391 : _665;
    assign _4068 = _1381 == _4077;
    assign _4069 = _1376 & _4068;
    assign _4074 = _4069 ? _1394 : _4073;
    assign _4065 = _299 == _4077;
    assign _4066 = _1376 & _4065;
    assign _4076 = _4066 ? _1099 : _4074;
    assign _4082 = _285 ? _4081 : _4076;
    assign _149 = _4082;
    always @(posedge _277) begin
        if (_275)
            _665 <= _1099;
        else
            _665 <= _149;
    end
    assign _4096 = 8'b01110001;
    assign _4097 = _280 == _4096;
    assign _4100 = _4097 ? _6252 : _1099;
    assign _4090 = _1386 == _4096;
    assign _4091 = _1376 & _4090;
    assign _4092 = _4091 ? _1391 : _662;
    assign _4087 = _1381 == _4096;
    assign _4088 = _1376 & _4087;
    assign _4093 = _4088 ? _1394 : _4092;
    assign _4084 = _299 == _4096;
    assign _4085 = _1376 & _4084;
    assign _4095 = _4085 ? _1099 : _4093;
    assign _4101 = _285 ? _4100 : _4095;
    assign _150 = _4101;
    always @(posedge _277) begin
        if (_275)
            _662 <= _1099;
        else
            _662 <= _150;
    end
    assign _4115 = 8'b01110000;
    assign _4116 = _280 == _4115;
    assign _4119 = _4116 ? _6252 : _1099;
    assign _4109 = _1386 == _4115;
    assign _4110 = _1376 & _4109;
    assign _4111 = _4110 ? _1391 : _659;
    assign _4106 = _1381 == _4115;
    assign _4107 = _1376 & _4106;
    assign _4112 = _4107 ? _1394 : _4111;
    assign _4103 = _299 == _4115;
    assign _4104 = _1376 & _4103;
    assign _4114 = _4104 ? _1099 : _4112;
    assign _4120 = _285 ? _4119 : _4114;
    assign _151 = _4120;
    always @(posedge _277) begin
        if (_275)
            _659 <= _1099;
        else
            _659 <= _151;
    end
    assign _4134 = 8'b01101111;
    assign _4135 = _280 == _4134;
    assign _4138 = _4135 ? _6252 : _1099;
    assign _4128 = _1386 == _4134;
    assign _4129 = _1376 & _4128;
    assign _4130 = _4129 ? _1391 : _656;
    assign _4125 = _1381 == _4134;
    assign _4126 = _1376 & _4125;
    assign _4131 = _4126 ? _1394 : _4130;
    assign _4122 = _299 == _4134;
    assign _4123 = _1376 & _4122;
    assign _4133 = _4123 ? _1099 : _4131;
    assign _4139 = _285 ? _4138 : _4133;
    assign _152 = _4139;
    always @(posedge _277) begin
        if (_275)
            _656 <= _1099;
        else
            _656 <= _152;
    end
    assign _4153 = 8'b01101110;
    assign _4154 = _280 == _4153;
    assign _4157 = _4154 ? _6252 : _1099;
    assign _4147 = _1386 == _4153;
    assign _4148 = _1376 & _4147;
    assign _4149 = _4148 ? _1391 : _653;
    assign _4144 = _1381 == _4153;
    assign _4145 = _1376 & _4144;
    assign _4150 = _4145 ? _1394 : _4149;
    assign _4141 = _299 == _4153;
    assign _4142 = _1376 & _4141;
    assign _4152 = _4142 ? _1099 : _4150;
    assign _4158 = _285 ? _4157 : _4152;
    assign _153 = _4158;
    always @(posedge _277) begin
        if (_275)
            _653 <= _1099;
        else
            _653 <= _153;
    end
    assign _4172 = 8'b01101101;
    assign _4173 = _280 == _4172;
    assign _4176 = _4173 ? _6252 : _1099;
    assign _4166 = _1386 == _4172;
    assign _4167 = _1376 & _4166;
    assign _4168 = _4167 ? _1391 : _650;
    assign _4163 = _1381 == _4172;
    assign _4164 = _1376 & _4163;
    assign _4169 = _4164 ? _1394 : _4168;
    assign _4160 = _299 == _4172;
    assign _4161 = _1376 & _4160;
    assign _4171 = _4161 ? _1099 : _4169;
    assign _4177 = _285 ? _4176 : _4171;
    assign _154 = _4177;
    always @(posedge _277) begin
        if (_275)
            _650 <= _1099;
        else
            _650 <= _154;
    end
    assign _4191 = 8'b01101100;
    assign _4192 = _280 == _4191;
    assign _4195 = _4192 ? _6252 : _1099;
    assign _4185 = _1386 == _4191;
    assign _4186 = _1376 & _4185;
    assign _4187 = _4186 ? _1391 : _647;
    assign _4182 = _1381 == _4191;
    assign _4183 = _1376 & _4182;
    assign _4188 = _4183 ? _1394 : _4187;
    assign _4179 = _299 == _4191;
    assign _4180 = _1376 & _4179;
    assign _4190 = _4180 ? _1099 : _4188;
    assign _4196 = _285 ? _4195 : _4190;
    assign _155 = _4196;
    always @(posedge _277) begin
        if (_275)
            _647 <= _1099;
        else
            _647 <= _155;
    end
    assign _4210 = 8'b01101011;
    assign _4211 = _280 == _4210;
    assign _4214 = _4211 ? _6252 : _1099;
    assign _4204 = _1386 == _4210;
    assign _4205 = _1376 & _4204;
    assign _4206 = _4205 ? _1391 : _644;
    assign _4201 = _1381 == _4210;
    assign _4202 = _1376 & _4201;
    assign _4207 = _4202 ? _1394 : _4206;
    assign _4198 = _299 == _4210;
    assign _4199 = _1376 & _4198;
    assign _4209 = _4199 ? _1099 : _4207;
    assign _4215 = _285 ? _4214 : _4209;
    assign _156 = _4215;
    always @(posedge _277) begin
        if (_275)
            _644 <= _1099;
        else
            _644 <= _156;
    end
    assign _4229 = 8'b01101010;
    assign _4230 = _280 == _4229;
    assign _4233 = _4230 ? _6252 : _1099;
    assign _4223 = _1386 == _4229;
    assign _4224 = _1376 & _4223;
    assign _4225 = _4224 ? _1391 : _641;
    assign _4220 = _1381 == _4229;
    assign _4221 = _1376 & _4220;
    assign _4226 = _4221 ? _1394 : _4225;
    assign _4217 = _299 == _4229;
    assign _4218 = _1376 & _4217;
    assign _4228 = _4218 ? _1099 : _4226;
    assign _4234 = _285 ? _4233 : _4228;
    assign _157 = _4234;
    always @(posedge _277) begin
        if (_275)
            _641 <= _1099;
        else
            _641 <= _157;
    end
    assign _4248 = 8'b01101001;
    assign _4249 = _280 == _4248;
    assign _4252 = _4249 ? _6252 : _1099;
    assign _4242 = _1386 == _4248;
    assign _4243 = _1376 & _4242;
    assign _4244 = _4243 ? _1391 : _638;
    assign _4239 = _1381 == _4248;
    assign _4240 = _1376 & _4239;
    assign _4245 = _4240 ? _1394 : _4244;
    assign _4236 = _299 == _4248;
    assign _4237 = _1376 & _4236;
    assign _4247 = _4237 ? _1099 : _4245;
    assign _4253 = _285 ? _4252 : _4247;
    assign _158 = _4253;
    always @(posedge _277) begin
        if (_275)
            _638 <= _1099;
        else
            _638 <= _158;
    end
    assign _4267 = 8'b01101000;
    assign _4268 = _280 == _4267;
    assign _4271 = _4268 ? _6252 : _1099;
    assign _4261 = _1386 == _4267;
    assign _4262 = _1376 & _4261;
    assign _4263 = _4262 ? _1391 : _635;
    assign _4258 = _1381 == _4267;
    assign _4259 = _1376 & _4258;
    assign _4264 = _4259 ? _1394 : _4263;
    assign _4255 = _299 == _4267;
    assign _4256 = _1376 & _4255;
    assign _4266 = _4256 ? _1099 : _4264;
    assign _4272 = _285 ? _4271 : _4266;
    assign _159 = _4272;
    always @(posedge _277) begin
        if (_275)
            _635 <= _1099;
        else
            _635 <= _159;
    end
    assign _4286 = 8'b01100111;
    assign _4287 = _280 == _4286;
    assign _4290 = _4287 ? _6252 : _1099;
    assign _4280 = _1386 == _4286;
    assign _4281 = _1376 & _4280;
    assign _4282 = _4281 ? _1391 : _632;
    assign _4277 = _1381 == _4286;
    assign _4278 = _1376 & _4277;
    assign _4283 = _4278 ? _1394 : _4282;
    assign _4274 = _299 == _4286;
    assign _4275 = _1376 & _4274;
    assign _4285 = _4275 ? _1099 : _4283;
    assign _4291 = _285 ? _4290 : _4285;
    assign _160 = _4291;
    always @(posedge _277) begin
        if (_275)
            _632 <= _1099;
        else
            _632 <= _160;
    end
    assign _4305 = 8'b01100110;
    assign _4306 = _280 == _4305;
    assign _4309 = _4306 ? _6252 : _1099;
    assign _4299 = _1386 == _4305;
    assign _4300 = _1376 & _4299;
    assign _4301 = _4300 ? _1391 : _629;
    assign _4296 = _1381 == _4305;
    assign _4297 = _1376 & _4296;
    assign _4302 = _4297 ? _1394 : _4301;
    assign _4293 = _299 == _4305;
    assign _4294 = _1376 & _4293;
    assign _4304 = _4294 ? _1099 : _4302;
    assign _4310 = _285 ? _4309 : _4304;
    assign _161 = _4310;
    always @(posedge _277) begin
        if (_275)
            _629 <= _1099;
        else
            _629 <= _161;
    end
    assign _4324 = 8'b01100101;
    assign _4325 = _280 == _4324;
    assign _4328 = _4325 ? _6252 : _1099;
    assign _4318 = _1386 == _4324;
    assign _4319 = _1376 & _4318;
    assign _4320 = _4319 ? _1391 : _626;
    assign _4315 = _1381 == _4324;
    assign _4316 = _1376 & _4315;
    assign _4321 = _4316 ? _1394 : _4320;
    assign _4312 = _299 == _4324;
    assign _4313 = _1376 & _4312;
    assign _4323 = _4313 ? _1099 : _4321;
    assign _4329 = _285 ? _4328 : _4323;
    assign _162 = _4329;
    always @(posedge _277) begin
        if (_275)
            _626 <= _1099;
        else
            _626 <= _162;
    end
    assign _4343 = 8'b01100100;
    assign _4344 = _280 == _4343;
    assign _4347 = _4344 ? _6252 : _1099;
    assign _4337 = _1386 == _4343;
    assign _4338 = _1376 & _4337;
    assign _4339 = _4338 ? _1391 : _623;
    assign _4334 = _1381 == _4343;
    assign _4335 = _1376 & _4334;
    assign _4340 = _4335 ? _1394 : _4339;
    assign _4331 = _299 == _4343;
    assign _4332 = _1376 & _4331;
    assign _4342 = _4332 ? _1099 : _4340;
    assign _4348 = _285 ? _4347 : _4342;
    assign _163 = _4348;
    always @(posedge _277) begin
        if (_275)
            _623 <= _1099;
        else
            _623 <= _163;
    end
    assign _4362 = 8'b01100011;
    assign _4363 = _280 == _4362;
    assign _4366 = _4363 ? _6252 : _1099;
    assign _4356 = _1386 == _4362;
    assign _4357 = _1376 & _4356;
    assign _4358 = _4357 ? _1391 : _620;
    assign _4353 = _1381 == _4362;
    assign _4354 = _1376 & _4353;
    assign _4359 = _4354 ? _1394 : _4358;
    assign _4350 = _299 == _4362;
    assign _4351 = _1376 & _4350;
    assign _4361 = _4351 ? _1099 : _4359;
    assign _4367 = _285 ? _4366 : _4361;
    assign _164 = _4367;
    always @(posedge _277) begin
        if (_275)
            _620 <= _1099;
        else
            _620 <= _164;
    end
    assign _4381 = 8'b01100010;
    assign _4382 = _280 == _4381;
    assign _4385 = _4382 ? _6252 : _1099;
    assign _4375 = _1386 == _4381;
    assign _4376 = _1376 & _4375;
    assign _4377 = _4376 ? _1391 : _617;
    assign _4372 = _1381 == _4381;
    assign _4373 = _1376 & _4372;
    assign _4378 = _4373 ? _1394 : _4377;
    assign _4369 = _299 == _4381;
    assign _4370 = _1376 & _4369;
    assign _4380 = _4370 ? _1099 : _4378;
    assign _4386 = _285 ? _4385 : _4380;
    assign _165 = _4386;
    always @(posedge _277) begin
        if (_275)
            _617 <= _1099;
        else
            _617 <= _165;
    end
    assign _4400 = 8'b01100001;
    assign _4401 = _280 == _4400;
    assign _4404 = _4401 ? _6252 : _1099;
    assign _4394 = _1386 == _4400;
    assign _4395 = _1376 & _4394;
    assign _4396 = _4395 ? _1391 : _614;
    assign _4391 = _1381 == _4400;
    assign _4392 = _1376 & _4391;
    assign _4397 = _4392 ? _1394 : _4396;
    assign _4388 = _299 == _4400;
    assign _4389 = _1376 & _4388;
    assign _4399 = _4389 ? _1099 : _4397;
    assign _4405 = _285 ? _4404 : _4399;
    assign _166 = _4405;
    always @(posedge _277) begin
        if (_275)
            _614 <= _1099;
        else
            _614 <= _166;
    end
    assign _4419 = 8'b01100000;
    assign _4420 = _280 == _4419;
    assign _4423 = _4420 ? _6252 : _1099;
    assign _4413 = _1386 == _4419;
    assign _4414 = _1376 & _4413;
    assign _4415 = _4414 ? _1391 : _611;
    assign _4410 = _1381 == _4419;
    assign _4411 = _1376 & _4410;
    assign _4416 = _4411 ? _1394 : _4415;
    assign _4407 = _299 == _4419;
    assign _4408 = _1376 & _4407;
    assign _4418 = _4408 ? _1099 : _4416;
    assign _4424 = _285 ? _4423 : _4418;
    assign _167 = _4424;
    always @(posedge _277) begin
        if (_275)
            _611 <= _1099;
        else
            _611 <= _167;
    end
    assign _4438 = 8'b01011111;
    assign _4439 = _280 == _4438;
    assign _4442 = _4439 ? _6252 : _1099;
    assign _4432 = _1386 == _4438;
    assign _4433 = _1376 & _4432;
    assign _4434 = _4433 ? _1391 : _608;
    assign _4429 = _1381 == _4438;
    assign _4430 = _1376 & _4429;
    assign _4435 = _4430 ? _1394 : _4434;
    assign _4426 = _299 == _4438;
    assign _4427 = _1376 & _4426;
    assign _4437 = _4427 ? _1099 : _4435;
    assign _4443 = _285 ? _4442 : _4437;
    assign _168 = _4443;
    always @(posedge _277) begin
        if (_275)
            _608 <= _1099;
        else
            _608 <= _168;
    end
    assign _4457 = 8'b01011110;
    assign _4458 = _280 == _4457;
    assign _4461 = _4458 ? _6252 : _1099;
    assign _4451 = _1386 == _4457;
    assign _4452 = _1376 & _4451;
    assign _4453 = _4452 ? _1391 : _605;
    assign _4448 = _1381 == _4457;
    assign _4449 = _1376 & _4448;
    assign _4454 = _4449 ? _1394 : _4453;
    assign _4445 = _299 == _4457;
    assign _4446 = _1376 & _4445;
    assign _4456 = _4446 ? _1099 : _4454;
    assign _4462 = _285 ? _4461 : _4456;
    assign _169 = _4462;
    always @(posedge _277) begin
        if (_275)
            _605 <= _1099;
        else
            _605 <= _169;
    end
    assign _4476 = 8'b01011101;
    assign _4477 = _280 == _4476;
    assign _4480 = _4477 ? _6252 : _1099;
    assign _4470 = _1386 == _4476;
    assign _4471 = _1376 & _4470;
    assign _4472 = _4471 ? _1391 : _602;
    assign _4467 = _1381 == _4476;
    assign _4468 = _1376 & _4467;
    assign _4473 = _4468 ? _1394 : _4472;
    assign _4464 = _299 == _4476;
    assign _4465 = _1376 & _4464;
    assign _4475 = _4465 ? _1099 : _4473;
    assign _4481 = _285 ? _4480 : _4475;
    assign _170 = _4481;
    always @(posedge _277) begin
        if (_275)
            _602 <= _1099;
        else
            _602 <= _170;
    end
    assign _4495 = 8'b01011100;
    assign _4496 = _280 == _4495;
    assign _4499 = _4496 ? _6252 : _1099;
    assign _4489 = _1386 == _4495;
    assign _4490 = _1376 & _4489;
    assign _4491 = _4490 ? _1391 : _599;
    assign _4486 = _1381 == _4495;
    assign _4487 = _1376 & _4486;
    assign _4492 = _4487 ? _1394 : _4491;
    assign _4483 = _299 == _4495;
    assign _4484 = _1376 & _4483;
    assign _4494 = _4484 ? _1099 : _4492;
    assign _4500 = _285 ? _4499 : _4494;
    assign _171 = _4500;
    always @(posedge _277) begin
        if (_275)
            _599 <= _1099;
        else
            _599 <= _171;
    end
    assign _4514 = 8'b01011011;
    assign _4515 = _280 == _4514;
    assign _4518 = _4515 ? _6252 : _1099;
    assign _4508 = _1386 == _4514;
    assign _4509 = _1376 & _4508;
    assign _4510 = _4509 ? _1391 : _596;
    assign _4505 = _1381 == _4514;
    assign _4506 = _1376 & _4505;
    assign _4511 = _4506 ? _1394 : _4510;
    assign _4502 = _299 == _4514;
    assign _4503 = _1376 & _4502;
    assign _4513 = _4503 ? _1099 : _4511;
    assign _4519 = _285 ? _4518 : _4513;
    assign _172 = _4519;
    always @(posedge _277) begin
        if (_275)
            _596 <= _1099;
        else
            _596 <= _172;
    end
    assign _4533 = 8'b01011010;
    assign _4534 = _280 == _4533;
    assign _4537 = _4534 ? _6252 : _1099;
    assign _4527 = _1386 == _4533;
    assign _4528 = _1376 & _4527;
    assign _4529 = _4528 ? _1391 : _593;
    assign _4524 = _1381 == _4533;
    assign _4525 = _1376 & _4524;
    assign _4530 = _4525 ? _1394 : _4529;
    assign _4521 = _299 == _4533;
    assign _4522 = _1376 & _4521;
    assign _4532 = _4522 ? _1099 : _4530;
    assign _4538 = _285 ? _4537 : _4532;
    assign _173 = _4538;
    always @(posedge _277) begin
        if (_275)
            _593 <= _1099;
        else
            _593 <= _173;
    end
    assign _4552 = 8'b01011001;
    assign _4553 = _280 == _4552;
    assign _4556 = _4553 ? _6252 : _1099;
    assign _4546 = _1386 == _4552;
    assign _4547 = _1376 & _4546;
    assign _4548 = _4547 ? _1391 : _590;
    assign _4543 = _1381 == _4552;
    assign _4544 = _1376 & _4543;
    assign _4549 = _4544 ? _1394 : _4548;
    assign _4540 = _299 == _4552;
    assign _4541 = _1376 & _4540;
    assign _4551 = _4541 ? _1099 : _4549;
    assign _4557 = _285 ? _4556 : _4551;
    assign _174 = _4557;
    always @(posedge _277) begin
        if (_275)
            _590 <= _1099;
        else
            _590 <= _174;
    end
    assign _4571 = 8'b01011000;
    assign _4572 = _280 == _4571;
    assign _4575 = _4572 ? _6252 : _1099;
    assign _4565 = _1386 == _4571;
    assign _4566 = _1376 & _4565;
    assign _4567 = _4566 ? _1391 : _587;
    assign _4562 = _1381 == _4571;
    assign _4563 = _1376 & _4562;
    assign _4568 = _4563 ? _1394 : _4567;
    assign _4559 = _299 == _4571;
    assign _4560 = _1376 & _4559;
    assign _4570 = _4560 ? _1099 : _4568;
    assign _4576 = _285 ? _4575 : _4570;
    assign _175 = _4576;
    always @(posedge _277) begin
        if (_275)
            _587 <= _1099;
        else
            _587 <= _175;
    end
    assign _4590 = 8'b01010111;
    assign _4591 = _280 == _4590;
    assign _4594 = _4591 ? _6252 : _1099;
    assign _4584 = _1386 == _4590;
    assign _4585 = _1376 & _4584;
    assign _4586 = _4585 ? _1391 : _584;
    assign _4581 = _1381 == _4590;
    assign _4582 = _1376 & _4581;
    assign _4587 = _4582 ? _1394 : _4586;
    assign _4578 = _299 == _4590;
    assign _4579 = _1376 & _4578;
    assign _4589 = _4579 ? _1099 : _4587;
    assign _4595 = _285 ? _4594 : _4589;
    assign _176 = _4595;
    always @(posedge _277) begin
        if (_275)
            _584 <= _1099;
        else
            _584 <= _176;
    end
    assign _4609 = 8'b01010110;
    assign _4610 = _280 == _4609;
    assign _4613 = _4610 ? _6252 : _1099;
    assign _4603 = _1386 == _4609;
    assign _4604 = _1376 & _4603;
    assign _4605 = _4604 ? _1391 : _581;
    assign _4600 = _1381 == _4609;
    assign _4601 = _1376 & _4600;
    assign _4606 = _4601 ? _1394 : _4605;
    assign _4597 = _299 == _4609;
    assign _4598 = _1376 & _4597;
    assign _4608 = _4598 ? _1099 : _4606;
    assign _4614 = _285 ? _4613 : _4608;
    assign _177 = _4614;
    always @(posedge _277) begin
        if (_275)
            _581 <= _1099;
        else
            _581 <= _177;
    end
    assign _4628 = 8'b01010101;
    assign _4629 = _280 == _4628;
    assign _4632 = _4629 ? _6252 : _1099;
    assign _4622 = _1386 == _4628;
    assign _4623 = _1376 & _4622;
    assign _4624 = _4623 ? _1391 : _578;
    assign _4619 = _1381 == _4628;
    assign _4620 = _1376 & _4619;
    assign _4625 = _4620 ? _1394 : _4624;
    assign _4616 = _299 == _4628;
    assign _4617 = _1376 & _4616;
    assign _4627 = _4617 ? _1099 : _4625;
    assign _4633 = _285 ? _4632 : _4627;
    assign _178 = _4633;
    always @(posedge _277) begin
        if (_275)
            _578 <= _1099;
        else
            _578 <= _178;
    end
    assign _4647 = 8'b01010100;
    assign _4648 = _280 == _4647;
    assign _4651 = _4648 ? _6252 : _1099;
    assign _4641 = _1386 == _4647;
    assign _4642 = _1376 & _4641;
    assign _4643 = _4642 ? _1391 : _575;
    assign _4638 = _1381 == _4647;
    assign _4639 = _1376 & _4638;
    assign _4644 = _4639 ? _1394 : _4643;
    assign _4635 = _299 == _4647;
    assign _4636 = _1376 & _4635;
    assign _4646 = _4636 ? _1099 : _4644;
    assign _4652 = _285 ? _4651 : _4646;
    assign _179 = _4652;
    always @(posedge _277) begin
        if (_275)
            _575 <= _1099;
        else
            _575 <= _179;
    end
    assign _4666 = 8'b01010011;
    assign _4667 = _280 == _4666;
    assign _4670 = _4667 ? _6252 : _1099;
    assign _4660 = _1386 == _4666;
    assign _4661 = _1376 & _4660;
    assign _4662 = _4661 ? _1391 : _572;
    assign _4657 = _1381 == _4666;
    assign _4658 = _1376 & _4657;
    assign _4663 = _4658 ? _1394 : _4662;
    assign _4654 = _299 == _4666;
    assign _4655 = _1376 & _4654;
    assign _4665 = _4655 ? _1099 : _4663;
    assign _4671 = _285 ? _4670 : _4665;
    assign _180 = _4671;
    always @(posedge _277) begin
        if (_275)
            _572 <= _1099;
        else
            _572 <= _180;
    end
    assign _4685 = 8'b01010010;
    assign _4686 = _280 == _4685;
    assign _4689 = _4686 ? _6252 : _1099;
    assign _4679 = _1386 == _4685;
    assign _4680 = _1376 & _4679;
    assign _4681 = _4680 ? _1391 : _569;
    assign _4676 = _1381 == _4685;
    assign _4677 = _1376 & _4676;
    assign _4682 = _4677 ? _1394 : _4681;
    assign _4673 = _299 == _4685;
    assign _4674 = _1376 & _4673;
    assign _4684 = _4674 ? _1099 : _4682;
    assign _4690 = _285 ? _4689 : _4684;
    assign _181 = _4690;
    always @(posedge _277) begin
        if (_275)
            _569 <= _1099;
        else
            _569 <= _181;
    end
    assign _4704 = 8'b01010001;
    assign _4705 = _280 == _4704;
    assign _4708 = _4705 ? _6252 : _1099;
    assign _4698 = _1386 == _4704;
    assign _4699 = _1376 & _4698;
    assign _4700 = _4699 ? _1391 : _566;
    assign _4695 = _1381 == _4704;
    assign _4696 = _1376 & _4695;
    assign _4701 = _4696 ? _1394 : _4700;
    assign _4692 = _299 == _4704;
    assign _4693 = _1376 & _4692;
    assign _4703 = _4693 ? _1099 : _4701;
    assign _4709 = _285 ? _4708 : _4703;
    assign _182 = _4709;
    always @(posedge _277) begin
        if (_275)
            _566 <= _1099;
        else
            _566 <= _182;
    end
    assign _4723 = 8'b01010000;
    assign _4724 = _280 == _4723;
    assign _4727 = _4724 ? _6252 : _1099;
    assign _4717 = _1386 == _4723;
    assign _4718 = _1376 & _4717;
    assign _4719 = _4718 ? _1391 : _563;
    assign _4714 = _1381 == _4723;
    assign _4715 = _1376 & _4714;
    assign _4720 = _4715 ? _1394 : _4719;
    assign _4711 = _299 == _4723;
    assign _4712 = _1376 & _4711;
    assign _4722 = _4712 ? _1099 : _4720;
    assign _4728 = _285 ? _4727 : _4722;
    assign _183 = _4728;
    always @(posedge _277) begin
        if (_275)
            _563 <= _1099;
        else
            _563 <= _183;
    end
    assign _4742 = 8'b01001111;
    assign _4743 = _280 == _4742;
    assign _4746 = _4743 ? _6252 : _1099;
    assign _4736 = _1386 == _4742;
    assign _4737 = _1376 & _4736;
    assign _4738 = _4737 ? _1391 : _560;
    assign _4733 = _1381 == _4742;
    assign _4734 = _1376 & _4733;
    assign _4739 = _4734 ? _1394 : _4738;
    assign _4730 = _299 == _4742;
    assign _4731 = _1376 & _4730;
    assign _4741 = _4731 ? _1099 : _4739;
    assign _4747 = _285 ? _4746 : _4741;
    assign _184 = _4747;
    always @(posedge _277) begin
        if (_275)
            _560 <= _1099;
        else
            _560 <= _184;
    end
    assign _4761 = 8'b01001110;
    assign _4762 = _280 == _4761;
    assign _4765 = _4762 ? _6252 : _1099;
    assign _4755 = _1386 == _4761;
    assign _4756 = _1376 & _4755;
    assign _4757 = _4756 ? _1391 : _557;
    assign _4752 = _1381 == _4761;
    assign _4753 = _1376 & _4752;
    assign _4758 = _4753 ? _1394 : _4757;
    assign _4749 = _299 == _4761;
    assign _4750 = _1376 & _4749;
    assign _4760 = _4750 ? _1099 : _4758;
    assign _4766 = _285 ? _4765 : _4760;
    assign _185 = _4766;
    always @(posedge _277) begin
        if (_275)
            _557 <= _1099;
        else
            _557 <= _185;
    end
    assign _4780 = 8'b01001101;
    assign _4781 = _280 == _4780;
    assign _4784 = _4781 ? _6252 : _1099;
    assign _4774 = _1386 == _4780;
    assign _4775 = _1376 & _4774;
    assign _4776 = _4775 ? _1391 : _554;
    assign _4771 = _1381 == _4780;
    assign _4772 = _1376 & _4771;
    assign _4777 = _4772 ? _1394 : _4776;
    assign _4768 = _299 == _4780;
    assign _4769 = _1376 & _4768;
    assign _4779 = _4769 ? _1099 : _4777;
    assign _4785 = _285 ? _4784 : _4779;
    assign _186 = _4785;
    always @(posedge _277) begin
        if (_275)
            _554 <= _1099;
        else
            _554 <= _186;
    end
    assign _4799 = 8'b01001100;
    assign _4800 = _280 == _4799;
    assign _4803 = _4800 ? _6252 : _1099;
    assign _4793 = _1386 == _4799;
    assign _4794 = _1376 & _4793;
    assign _4795 = _4794 ? _1391 : _551;
    assign _4790 = _1381 == _4799;
    assign _4791 = _1376 & _4790;
    assign _4796 = _4791 ? _1394 : _4795;
    assign _4787 = _299 == _4799;
    assign _4788 = _1376 & _4787;
    assign _4798 = _4788 ? _1099 : _4796;
    assign _4804 = _285 ? _4803 : _4798;
    assign _187 = _4804;
    always @(posedge _277) begin
        if (_275)
            _551 <= _1099;
        else
            _551 <= _187;
    end
    assign _4818 = 8'b01001011;
    assign _4819 = _280 == _4818;
    assign _4822 = _4819 ? _6252 : _1099;
    assign _4812 = _1386 == _4818;
    assign _4813 = _1376 & _4812;
    assign _4814 = _4813 ? _1391 : _548;
    assign _4809 = _1381 == _4818;
    assign _4810 = _1376 & _4809;
    assign _4815 = _4810 ? _1394 : _4814;
    assign _4806 = _299 == _4818;
    assign _4807 = _1376 & _4806;
    assign _4817 = _4807 ? _1099 : _4815;
    assign _4823 = _285 ? _4822 : _4817;
    assign _188 = _4823;
    always @(posedge _277) begin
        if (_275)
            _548 <= _1099;
        else
            _548 <= _188;
    end
    assign _4837 = 8'b01001010;
    assign _4838 = _280 == _4837;
    assign _4841 = _4838 ? _6252 : _1099;
    assign _4831 = _1386 == _4837;
    assign _4832 = _1376 & _4831;
    assign _4833 = _4832 ? _1391 : _545;
    assign _4828 = _1381 == _4837;
    assign _4829 = _1376 & _4828;
    assign _4834 = _4829 ? _1394 : _4833;
    assign _4825 = _299 == _4837;
    assign _4826 = _1376 & _4825;
    assign _4836 = _4826 ? _1099 : _4834;
    assign _4842 = _285 ? _4841 : _4836;
    assign _189 = _4842;
    always @(posedge _277) begin
        if (_275)
            _545 <= _1099;
        else
            _545 <= _189;
    end
    assign _4856 = 8'b01001001;
    assign _4857 = _280 == _4856;
    assign _4860 = _4857 ? _6252 : _1099;
    assign _4850 = _1386 == _4856;
    assign _4851 = _1376 & _4850;
    assign _4852 = _4851 ? _1391 : _542;
    assign _4847 = _1381 == _4856;
    assign _4848 = _1376 & _4847;
    assign _4853 = _4848 ? _1394 : _4852;
    assign _4844 = _299 == _4856;
    assign _4845 = _1376 & _4844;
    assign _4855 = _4845 ? _1099 : _4853;
    assign _4861 = _285 ? _4860 : _4855;
    assign _190 = _4861;
    always @(posedge _277) begin
        if (_275)
            _542 <= _1099;
        else
            _542 <= _190;
    end
    assign _4875 = 8'b01001000;
    assign _4876 = _280 == _4875;
    assign _4879 = _4876 ? _6252 : _1099;
    assign _4869 = _1386 == _4875;
    assign _4870 = _1376 & _4869;
    assign _4871 = _4870 ? _1391 : _539;
    assign _4866 = _1381 == _4875;
    assign _4867 = _1376 & _4866;
    assign _4872 = _4867 ? _1394 : _4871;
    assign _4863 = _299 == _4875;
    assign _4864 = _1376 & _4863;
    assign _4874 = _4864 ? _1099 : _4872;
    assign _4880 = _285 ? _4879 : _4874;
    assign _191 = _4880;
    always @(posedge _277) begin
        if (_275)
            _539 <= _1099;
        else
            _539 <= _191;
    end
    assign _4894 = 8'b01000111;
    assign _4895 = _280 == _4894;
    assign _4898 = _4895 ? _6252 : _1099;
    assign _4888 = _1386 == _4894;
    assign _4889 = _1376 & _4888;
    assign _4890 = _4889 ? _1391 : _536;
    assign _4885 = _1381 == _4894;
    assign _4886 = _1376 & _4885;
    assign _4891 = _4886 ? _1394 : _4890;
    assign _4882 = _299 == _4894;
    assign _4883 = _1376 & _4882;
    assign _4893 = _4883 ? _1099 : _4891;
    assign _4899 = _285 ? _4898 : _4893;
    assign _192 = _4899;
    always @(posedge _277) begin
        if (_275)
            _536 <= _1099;
        else
            _536 <= _192;
    end
    assign _4913 = 8'b01000110;
    assign _4914 = _280 == _4913;
    assign _4917 = _4914 ? _6252 : _1099;
    assign _4907 = _1386 == _4913;
    assign _4908 = _1376 & _4907;
    assign _4909 = _4908 ? _1391 : _533;
    assign _4904 = _1381 == _4913;
    assign _4905 = _1376 & _4904;
    assign _4910 = _4905 ? _1394 : _4909;
    assign _4901 = _299 == _4913;
    assign _4902 = _1376 & _4901;
    assign _4912 = _4902 ? _1099 : _4910;
    assign _4918 = _285 ? _4917 : _4912;
    assign _193 = _4918;
    always @(posedge _277) begin
        if (_275)
            _533 <= _1099;
        else
            _533 <= _193;
    end
    assign _4932 = 8'b01000101;
    assign _4933 = _280 == _4932;
    assign _4936 = _4933 ? _6252 : _1099;
    assign _4926 = _1386 == _4932;
    assign _4927 = _1376 & _4926;
    assign _4928 = _4927 ? _1391 : _530;
    assign _4923 = _1381 == _4932;
    assign _4924 = _1376 & _4923;
    assign _4929 = _4924 ? _1394 : _4928;
    assign _4920 = _299 == _4932;
    assign _4921 = _1376 & _4920;
    assign _4931 = _4921 ? _1099 : _4929;
    assign _4937 = _285 ? _4936 : _4931;
    assign _194 = _4937;
    always @(posedge _277) begin
        if (_275)
            _530 <= _1099;
        else
            _530 <= _194;
    end
    assign _4951 = 8'b01000100;
    assign _4952 = _280 == _4951;
    assign _4955 = _4952 ? _6252 : _1099;
    assign _4945 = _1386 == _4951;
    assign _4946 = _1376 & _4945;
    assign _4947 = _4946 ? _1391 : _527;
    assign _4942 = _1381 == _4951;
    assign _4943 = _1376 & _4942;
    assign _4948 = _4943 ? _1394 : _4947;
    assign _4939 = _299 == _4951;
    assign _4940 = _1376 & _4939;
    assign _4950 = _4940 ? _1099 : _4948;
    assign _4956 = _285 ? _4955 : _4950;
    assign _195 = _4956;
    always @(posedge _277) begin
        if (_275)
            _527 <= _1099;
        else
            _527 <= _195;
    end
    assign _4970 = 8'b01000011;
    assign _4971 = _280 == _4970;
    assign _4974 = _4971 ? _6252 : _1099;
    assign _4964 = _1386 == _4970;
    assign _4965 = _1376 & _4964;
    assign _4966 = _4965 ? _1391 : _524;
    assign _4961 = _1381 == _4970;
    assign _4962 = _1376 & _4961;
    assign _4967 = _4962 ? _1394 : _4966;
    assign _4958 = _299 == _4970;
    assign _4959 = _1376 & _4958;
    assign _4969 = _4959 ? _1099 : _4967;
    assign _4975 = _285 ? _4974 : _4969;
    assign _196 = _4975;
    always @(posedge _277) begin
        if (_275)
            _524 <= _1099;
        else
            _524 <= _196;
    end
    assign _4989 = 8'b01000010;
    assign _4990 = _280 == _4989;
    assign _4993 = _4990 ? _6252 : _1099;
    assign _4983 = _1386 == _4989;
    assign _4984 = _1376 & _4983;
    assign _4985 = _4984 ? _1391 : _521;
    assign _4980 = _1381 == _4989;
    assign _4981 = _1376 & _4980;
    assign _4986 = _4981 ? _1394 : _4985;
    assign _4977 = _299 == _4989;
    assign _4978 = _1376 & _4977;
    assign _4988 = _4978 ? _1099 : _4986;
    assign _4994 = _285 ? _4993 : _4988;
    assign _197 = _4994;
    always @(posedge _277) begin
        if (_275)
            _521 <= _1099;
        else
            _521 <= _197;
    end
    assign _5008 = 8'b01000001;
    assign _5009 = _280 == _5008;
    assign _5012 = _5009 ? _6252 : _1099;
    assign _5002 = _1386 == _5008;
    assign _5003 = _1376 & _5002;
    assign _5004 = _5003 ? _1391 : _518;
    assign _4999 = _1381 == _5008;
    assign _5000 = _1376 & _4999;
    assign _5005 = _5000 ? _1394 : _5004;
    assign _4996 = _299 == _5008;
    assign _4997 = _1376 & _4996;
    assign _5007 = _4997 ? _1099 : _5005;
    assign _5013 = _285 ? _5012 : _5007;
    assign _198 = _5013;
    always @(posedge _277) begin
        if (_275)
            _518 <= _1099;
        else
            _518 <= _198;
    end
    assign _5027 = 8'b01000000;
    assign _5028 = _280 == _5027;
    assign _5031 = _5028 ? _6252 : _1099;
    assign _5021 = _1386 == _5027;
    assign _5022 = _1376 & _5021;
    assign _5023 = _5022 ? _1391 : _515;
    assign _5018 = _1381 == _5027;
    assign _5019 = _1376 & _5018;
    assign _5024 = _5019 ? _1394 : _5023;
    assign _5015 = _299 == _5027;
    assign _5016 = _1376 & _5015;
    assign _5026 = _5016 ? _1099 : _5024;
    assign _5032 = _285 ? _5031 : _5026;
    assign _199 = _5032;
    always @(posedge _277) begin
        if (_275)
            _515 <= _1099;
        else
            _515 <= _199;
    end
    assign _5046 = 8'b00111111;
    assign _5047 = _280 == _5046;
    assign _5050 = _5047 ? _6252 : _1099;
    assign _5040 = _1386 == _5046;
    assign _5041 = _1376 & _5040;
    assign _5042 = _5041 ? _1391 : _512;
    assign _5037 = _1381 == _5046;
    assign _5038 = _1376 & _5037;
    assign _5043 = _5038 ? _1394 : _5042;
    assign _5034 = _299 == _5046;
    assign _5035 = _1376 & _5034;
    assign _5045 = _5035 ? _1099 : _5043;
    assign _5051 = _285 ? _5050 : _5045;
    assign _200 = _5051;
    always @(posedge _277) begin
        if (_275)
            _512 <= _1099;
        else
            _512 <= _200;
    end
    assign _5065 = 8'b00111110;
    assign _5066 = _280 == _5065;
    assign _5069 = _5066 ? _6252 : _1099;
    assign _5059 = _1386 == _5065;
    assign _5060 = _1376 & _5059;
    assign _5061 = _5060 ? _1391 : _509;
    assign _5056 = _1381 == _5065;
    assign _5057 = _1376 & _5056;
    assign _5062 = _5057 ? _1394 : _5061;
    assign _5053 = _299 == _5065;
    assign _5054 = _1376 & _5053;
    assign _5064 = _5054 ? _1099 : _5062;
    assign _5070 = _285 ? _5069 : _5064;
    assign _201 = _5070;
    always @(posedge _277) begin
        if (_275)
            _509 <= _1099;
        else
            _509 <= _201;
    end
    assign _5084 = 8'b00111101;
    assign _5085 = _280 == _5084;
    assign _5088 = _5085 ? _6252 : _1099;
    assign _5078 = _1386 == _5084;
    assign _5079 = _1376 & _5078;
    assign _5080 = _5079 ? _1391 : _506;
    assign _5075 = _1381 == _5084;
    assign _5076 = _1376 & _5075;
    assign _5081 = _5076 ? _1394 : _5080;
    assign _5072 = _299 == _5084;
    assign _5073 = _1376 & _5072;
    assign _5083 = _5073 ? _1099 : _5081;
    assign _5089 = _285 ? _5088 : _5083;
    assign _202 = _5089;
    always @(posedge _277) begin
        if (_275)
            _506 <= _1099;
        else
            _506 <= _202;
    end
    assign _5103 = 8'b00111100;
    assign _5104 = _280 == _5103;
    assign _5107 = _5104 ? _6252 : _1099;
    assign _5097 = _1386 == _5103;
    assign _5098 = _1376 & _5097;
    assign _5099 = _5098 ? _1391 : _503;
    assign _5094 = _1381 == _5103;
    assign _5095 = _1376 & _5094;
    assign _5100 = _5095 ? _1394 : _5099;
    assign _5091 = _299 == _5103;
    assign _5092 = _1376 & _5091;
    assign _5102 = _5092 ? _1099 : _5100;
    assign _5108 = _285 ? _5107 : _5102;
    assign _203 = _5108;
    always @(posedge _277) begin
        if (_275)
            _503 <= _1099;
        else
            _503 <= _203;
    end
    assign _5122 = 8'b00111011;
    assign _5123 = _280 == _5122;
    assign _5126 = _5123 ? _6252 : _1099;
    assign _5116 = _1386 == _5122;
    assign _5117 = _1376 & _5116;
    assign _5118 = _5117 ? _1391 : _500;
    assign _5113 = _1381 == _5122;
    assign _5114 = _1376 & _5113;
    assign _5119 = _5114 ? _1394 : _5118;
    assign _5110 = _299 == _5122;
    assign _5111 = _1376 & _5110;
    assign _5121 = _5111 ? _1099 : _5119;
    assign _5127 = _285 ? _5126 : _5121;
    assign _204 = _5127;
    always @(posedge _277) begin
        if (_275)
            _500 <= _1099;
        else
            _500 <= _204;
    end
    assign _5141 = 8'b00111010;
    assign _5142 = _280 == _5141;
    assign _5145 = _5142 ? _6252 : _1099;
    assign _5135 = _1386 == _5141;
    assign _5136 = _1376 & _5135;
    assign _5137 = _5136 ? _1391 : _497;
    assign _5132 = _1381 == _5141;
    assign _5133 = _1376 & _5132;
    assign _5138 = _5133 ? _1394 : _5137;
    assign _5129 = _299 == _5141;
    assign _5130 = _1376 & _5129;
    assign _5140 = _5130 ? _1099 : _5138;
    assign _5146 = _285 ? _5145 : _5140;
    assign _205 = _5146;
    always @(posedge _277) begin
        if (_275)
            _497 <= _1099;
        else
            _497 <= _205;
    end
    assign _5160 = 8'b00111001;
    assign _5161 = _280 == _5160;
    assign _5164 = _5161 ? _6252 : _1099;
    assign _5154 = _1386 == _5160;
    assign _5155 = _1376 & _5154;
    assign _5156 = _5155 ? _1391 : _494;
    assign _5151 = _1381 == _5160;
    assign _5152 = _1376 & _5151;
    assign _5157 = _5152 ? _1394 : _5156;
    assign _5148 = _299 == _5160;
    assign _5149 = _1376 & _5148;
    assign _5159 = _5149 ? _1099 : _5157;
    assign _5165 = _285 ? _5164 : _5159;
    assign _206 = _5165;
    always @(posedge _277) begin
        if (_275)
            _494 <= _1099;
        else
            _494 <= _206;
    end
    assign _5179 = 8'b00111000;
    assign _5180 = _280 == _5179;
    assign _5183 = _5180 ? _6252 : _1099;
    assign _5173 = _1386 == _5179;
    assign _5174 = _1376 & _5173;
    assign _5175 = _5174 ? _1391 : _491;
    assign _5170 = _1381 == _5179;
    assign _5171 = _1376 & _5170;
    assign _5176 = _5171 ? _1394 : _5175;
    assign _5167 = _299 == _5179;
    assign _5168 = _1376 & _5167;
    assign _5178 = _5168 ? _1099 : _5176;
    assign _5184 = _285 ? _5183 : _5178;
    assign _207 = _5184;
    always @(posedge _277) begin
        if (_275)
            _491 <= _1099;
        else
            _491 <= _207;
    end
    assign _5198 = 8'b00110111;
    assign _5199 = _280 == _5198;
    assign _5202 = _5199 ? _6252 : _1099;
    assign _5192 = _1386 == _5198;
    assign _5193 = _1376 & _5192;
    assign _5194 = _5193 ? _1391 : _488;
    assign _5189 = _1381 == _5198;
    assign _5190 = _1376 & _5189;
    assign _5195 = _5190 ? _1394 : _5194;
    assign _5186 = _299 == _5198;
    assign _5187 = _1376 & _5186;
    assign _5197 = _5187 ? _1099 : _5195;
    assign _5203 = _285 ? _5202 : _5197;
    assign _208 = _5203;
    always @(posedge _277) begin
        if (_275)
            _488 <= _1099;
        else
            _488 <= _208;
    end
    assign _5217 = 8'b00110110;
    assign _5218 = _280 == _5217;
    assign _5221 = _5218 ? _6252 : _1099;
    assign _5211 = _1386 == _5217;
    assign _5212 = _1376 & _5211;
    assign _5213 = _5212 ? _1391 : _485;
    assign _5208 = _1381 == _5217;
    assign _5209 = _1376 & _5208;
    assign _5214 = _5209 ? _1394 : _5213;
    assign _5205 = _299 == _5217;
    assign _5206 = _1376 & _5205;
    assign _5216 = _5206 ? _1099 : _5214;
    assign _5222 = _285 ? _5221 : _5216;
    assign _209 = _5222;
    always @(posedge _277) begin
        if (_275)
            _485 <= _1099;
        else
            _485 <= _209;
    end
    assign _5236 = 8'b00110101;
    assign _5237 = _280 == _5236;
    assign _5240 = _5237 ? _6252 : _1099;
    assign _5230 = _1386 == _5236;
    assign _5231 = _1376 & _5230;
    assign _5232 = _5231 ? _1391 : _482;
    assign _5227 = _1381 == _5236;
    assign _5228 = _1376 & _5227;
    assign _5233 = _5228 ? _1394 : _5232;
    assign _5224 = _299 == _5236;
    assign _5225 = _1376 & _5224;
    assign _5235 = _5225 ? _1099 : _5233;
    assign _5241 = _285 ? _5240 : _5235;
    assign _210 = _5241;
    always @(posedge _277) begin
        if (_275)
            _482 <= _1099;
        else
            _482 <= _210;
    end
    assign _5255 = 8'b00110100;
    assign _5256 = _280 == _5255;
    assign _5259 = _5256 ? _6252 : _1099;
    assign _5249 = _1386 == _5255;
    assign _5250 = _1376 & _5249;
    assign _5251 = _5250 ? _1391 : _479;
    assign _5246 = _1381 == _5255;
    assign _5247 = _1376 & _5246;
    assign _5252 = _5247 ? _1394 : _5251;
    assign _5243 = _299 == _5255;
    assign _5244 = _1376 & _5243;
    assign _5254 = _5244 ? _1099 : _5252;
    assign _5260 = _285 ? _5259 : _5254;
    assign _211 = _5260;
    always @(posedge _277) begin
        if (_275)
            _479 <= _1099;
        else
            _479 <= _211;
    end
    assign _5274 = 8'b00110011;
    assign _5275 = _280 == _5274;
    assign _5278 = _5275 ? _6252 : _1099;
    assign _5268 = _1386 == _5274;
    assign _5269 = _1376 & _5268;
    assign _5270 = _5269 ? _1391 : _476;
    assign _5265 = _1381 == _5274;
    assign _5266 = _1376 & _5265;
    assign _5271 = _5266 ? _1394 : _5270;
    assign _5262 = _299 == _5274;
    assign _5263 = _1376 & _5262;
    assign _5273 = _5263 ? _1099 : _5271;
    assign _5279 = _285 ? _5278 : _5273;
    assign _212 = _5279;
    always @(posedge _277) begin
        if (_275)
            _476 <= _1099;
        else
            _476 <= _212;
    end
    assign _5293 = 8'b00110010;
    assign _5294 = _280 == _5293;
    assign _5297 = _5294 ? _6252 : _1099;
    assign _5287 = _1386 == _5293;
    assign _5288 = _1376 & _5287;
    assign _5289 = _5288 ? _1391 : _473;
    assign _5284 = _1381 == _5293;
    assign _5285 = _1376 & _5284;
    assign _5290 = _5285 ? _1394 : _5289;
    assign _5281 = _299 == _5293;
    assign _5282 = _1376 & _5281;
    assign _5292 = _5282 ? _1099 : _5290;
    assign _5298 = _285 ? _5297 : _5292;
    assign _213 = _5298;
    always @(posedge _277) begin
        if (_275)
            _473 <= _1099;
        else
            _473 <= _213;
    end
    assign _5312 = 8'b00110001;
    assign _5313 = _280 == _5312;
    assign _5316 = _5313 ? _6252 : _1099;
    assign _5306 = _1386 == _5312;
    assign _5307 = _1376 & _5306;
    assign _5308 = _5307 ? _1391 : _470;
    assign _5303 = _1381 == _5312;
    assign _5304 = _1376 & _5303;
    assign _5309 = _5304 ? _1394 : _5308;
    assign _5300 = _299 == _5312;
    assign _5301 = _1376 & _5300;
    assign _5311 = _5301 ? _1099 : _5309;
    assign _5317 = _285 ? _5316 : _5311;
    assign _214 = _5317;
    always @(posedge _277) begin
        if (_275)
            _470 <= _1099;
        else
            _470 <= _214;
    end
    assign _5331 = 8'b00110000;
    assign _5332 = _280 == _5331;
    assign _5335 = _5332 ? _6252 : _1099;
    assign _5325 = _1386 == _5331;
    assign _5326 = _1376 & _5325;
    assign _5327 = _5326 ? _1391 : _467;
    assign _5322 = _1381 == _5331;
    assign _5323 = _1376 & _5322;
    assign _5328 = _5323 ? _1394 : _5327;
    assign _5319 = _299 == _5331;
    assign _5320 = _1376 & _5319;
    assign _5330 = _5320 ? _1099 : _5328;
    assign _5336 = _285 ? _5335 : _5330;
    assign _215 = _5336;
    always @(posedge _277) begin
        if (_275)
            _467 <= _1099;
        else
            _467 <= _215;
    end
    assign _5350 = 8'b00101111;
    assign _5351 = _280 == _5350;
    assign _5354 = _5351 ? _6252 : _1099;
    assign _5344 = _1386 == _5350;
    assign _5345 = _1376 & _5344;
    assign _5346 = _5345 ? _1391 : _464;
    assign _5341 = _1381 == _5350;
    assign _5342 = _1376 & _5341;
    assign _5347 = _5342 ? _1394 : _5346;
    assign _5338 = _299 == _5350;
    assign _5339 = _1376 & _5338;
    assign _5349 = _5339 ? _1099 : _5347;
    assign _5355 = _285 ? _5354 : _5349;
    assign _216 = _5355;
    always @(posedge _277) begin
        if (_275)
            _464 <= _1099;
        else
            _464 <= _216;
    end
    assign _5369 = 8'b00101110;
    assign _5370 = _280 == _5369;
    assign _5373 = _5370 ? _6252 : _1099;
    assign _5363 = _1386 == _5369;
    assign _5364 = _1376 & _5363;
    assign _5365 = _5364 ? _1391 : _461;
    assign _5360 = _1381 == _5369;
    assign _5361 = _1376 & _5360;
    assign _5366 = _5361 ? _1394 : _5365;
    assign _5357 = _299 == _5369;
    assign _5358 = _1376 & _5357;
    assign _5368 = _5358 ? _1099 : _5366;
    assign _5374 = _285 ? _5373 : _5368;
    assign _217 = _5374;
    always @(posedge _277) begin
        if (_275)
            _461 <= _1099;
        else
            _461 <= _217;
    end
    assign _5388 = 8'b00101101;
    assign _5389 = _280 == _5388;
    assign _5392 = _5389 ? _6252 : _1099;
    assign _5382 = _1386 == _5388;
    assign _5383 = _1376 & _5382;
    assign _5384 = _5383 ? _1391 : _458;
    assign _5379 = _1381 == _5388;
    assign _5380 = _1376 & _5379;
    assign _5385 = _5380 ? _1394 : _5384;
    assign _5376 = _299 == _5388;
    assign _5377 = _1376 & _5376;
    assign _5387 = _5377 ? _1099 : _5385;
    assign _5393 = _285 ? _5392 : _5387;
    assign _218 = _5393;
    always @(posedge _277) begin
        if (_275)
            _458 <= _1099;
        else
            _458 <= _218;
    end
    assign _5407 = 8'b00101100;
    assign _5408 = _280 == _5407;
    assign _5411 = _5408 ? _6252 : _1099;
    assign _5401 = _1386 == _5407;
    assign _5402 = _1376 & _5401;
    assign _5403 = _5402 ? _1391 : _455;
    assign _5398 = _1381 == _5407;
    assign _5399 = _1376 & _5398;
    assign _5404 = _5399 ? _1394 : _5403;
    assign _5395 = _299 == _5407;
    assign _5396 = _1376 & _5395;
    assign _5406 = _5396 ? _1099 : _5404;
    assign _5412 = _285 ? _5411 : _5406;
    assign _219 = _5412;
    always @(posedge _277) begin
        if (_275)
            _455 <= _1099;
        else
            _455 <= _219;
    end
    assign _5426 = 8'b00101011;
    assign _5427 = _280 == _5426;
    assign _5430 = _5427 ? _6252 : _1099;
    assign _5420 = _1386 == _5426;
    assign _5421 = _1376 & _5420;
    assign _5422 = _5421 ? _1391 : _452;
    assign _5417 = _1381 == _5426;
    assign _5418 = _1376 & _5417;
    assign _5423 = _5418 ? _1394 : _5422;
    assign _5414 = _299 == _5426;
    assign _5415 = _1376 & _5414;
    assign _5425 = _5415 ? _1099 : _5423;
    assign _5431 = _285 ? _5430 : _5425;
    assign _220 = _5431;
    always @(posedge _277) begin
        if (_275)
            _452 <= _1099;
        else
            _452 <= _220;
    end
    assign _5445 = 8'b00101010;
    assign _5446 = _280 == _5445;
    assign _5449 = _5446 ? _6252 : _1099;
    assign _5439 = _1386 == _5445;
    assign _5440 = _1376 & _5439;
    assign _5441 = _5440 ? _1391 : _449;
    assign _5436 = _1381 == _5445;
    assign _5437 = _1376 & _5436;
    assign _5442 = _5437 ? _1394 : _5441;
    assign _5433 = _299 == _5445;
    assign _5434 = _1376 & _5433;
    assign _5444 = _5434 ? _1099 : _5442;
    assign _5450 = _285 ? _5449 : _5444;
    assign _221 = _5450;
    always @(posedge _277) begin
        if (_275)
            _449 <= _1099;
        else
            _449 <= _221;
    end
    assign _5464 = 8'b00101001;
    assign _5465 = _280 == _5464;
    assign _5468 = _5465 ? _6252 : _1099;
    assign _5458 = _1386 == _5464;
    assign _5459 = _1376 & _5458;
    assign _5460 = _5459 ? _1391 : _446;
    assign _5455 = _1381 == _5464;
    assign _5456 = _1376 & _5455;
    assign _5461 = _5456 ? _1394 : _5460;
    assign _5452 = _299 == _5464;
    assign _5453 = _1376 & _5452;
    assign _5463 = _5453 ? _1099 : _5461;
    assign _5469 = _285 ? _5468 : _5463;
    assign _222 = _5469;
    always @(posedge _277) begin
        if (_275)
            _446 <= _1099;
        else
            _446 <= _222;
    end
    assign _5483 = 8'b00101000;
    assign _5484 = _280 == _5483;
    assign _5487 = _5484 ? _6252 : _1099;
    assign _5477 = _1386 == _5483;
    assign _5478 = _1376 & _5477;
    assign _5479 = _5478 ? _1391 : _443;
    assign _5474 = _1381 == _5483;
    assign _5475 = _1376 & _5474;
    assign _5480 = _5475 ? _1394 : _5479;
    assign _5471 = _299 == _5483;
    assign _5472 = _1376 & _5471;
    assign _5482 = _5472 ? _1099 : _5480;
    assign _5488 = _285 ? _5487 : _5482;
    assign _223 = _5488;
    always @(posedge _277) begin
        if (_275)
            _443 <= _1099;
        else
            _443 <= _223;
    end
    assign _5502 = 8'b00100111;
    assign _5503 = _280 == _5502;
    assign _5506 = _5503 ? _6252 : _1099;
    assign _5496 = _1386 == _5502;
    assign _5497 = _1376 & _5496;
    assign _5498 = _5497 ? _1391 : _440;
    assign _5493 = _1381 == _5502;
    assign _5494 = _1376 & _5493;
    assign _5499 = _5494 ? _1394 : _5498;
    assign _5490 = _299 == _5502;
    assign _5491 = _1376 & _5490;
    assign _5501 = _5491 ? _1099 : _5499;
    assign _5507 = _285 ? _5506 : _5501;
    assign _224 = _5507;
    always @(posedge _277) begin
        if (_275)
            _440 <= _1099;
        else
            _440 <= _224;
    end
    assign _5521 = 8'b00100110;
    assign _5522 = _280 == _5521;
    assign _5525 = _5522 ? _6252 : _1099;
    assign _5515 = _1386 == _5521;
    assign _5516 = _1376 & _5515;
    assign _5517 = _5516 ? _1391 : _437;
    assign _5512 = _1381 == _5521;
    assign _5513 = _1376 & _5512;
    assign _5518 = _5513 ? _1394 : _5517;
    assign _5509 = _299 == _5521;
    assign _5510 = _1376 & _5509;
    assign _5520 = _5510 ? _1099 : _5518;
    assign _5526 = _285 ? _5525 : _5520;
    assign _225 = _5526;
    always @(posedge _277) begin
        if (_275)
            _437 <= _1099;
        else
            _437 <= _225;
    end
    assign _5540 = 8'b00100101;
    assign _5541 = _280 == _5540;
    assign _5544 = _5541 ? _6252 : _1099;
    assign _5534 = _1386 == _5540;
    assign _5535 = _1376 & _5534;
    assign _5536 = _5535 ? _1391 : _434;
    assign _5531 = _1381 == _5540;
    assign _5532 = _1376 & _5531;
    assign _5537 = _5532 ? _1394 : _5536;
    assign _5528 = _299 == _5540;
    assign _5529 = _1376 & _5528;
    assign _5539 = _5529 ? _1099 : _5537;
    assign _5545 = _285 ? _5544 : _5539;
    assign _226 = _5545;
    always @(posedge _277) begin
        if (_275)
            _434 <= _1099;
        else
            _434 <= _226;
    end
    assign _5559 = 8'b00100100;
    assign _5560 = _280 == _5559;
    assign _5563 = _5560 ? _6252 : _1099;
    assign _5553 = _1386 == _5559;
    assign _5554 = _1376 & _5553;
    assign _5555 = _5554 ? _1391 : _431;
    assign _5550 = _1381 == _5559;
    assign _5551 = _1376 & _5550;
    assign _5556 = _5551 ? _1394 : _5555;
    assign _5547 = _299 == _5559;
    assign _5548 = _1376 & _5547;
    assign _5558 = _5548 ? _1099 : _5556;
    assign _5564 = _285 ? _5563 : _5558;
    assign _227 = _5564;
    always @(posedge _277) begin
        if (_275)
            _431 <= _1099;
        else
            _431 <= _227;
    end
    assign _5578 = 8'b00100011;
    assign _5579 = _280 == _5578;
    assign _5582 = _5579 ? _6252 : _1099;
    assign _5572 = _1386 == _5578;
    assign _5573 = _1376 & _5572;
    assign _5574 = _5573 ? _1391 : _428;
    assign _5569 = _1381 == _5578;
    assign _5570 = _1376 & _5569;
    assign _5575 = _5570 ? _1394 : _5574;
    assign _5566 = _299 == _5578;
    assign _5567 = _1376 & _5566;
    assign _5577 = _5567 ? _1099 : _5575;
    assign _5583 = _285 ? _5582 : _5577;
    assign _228 = _5583;
    always @(posedge _277) begin
        if (_275)
            _428 <= _1099;
        else
            _428 <= _228;
    end
    assign _5597 = 8'b00100010;
    assign _5598 = _280 == _5597;
    assign _5601 = _5598 ? _6252 : _1099;
    assign _5591 = _1386 == _5597;
    assign _5592 = _1376 & _5591;
    assign _5593 = _5592 ? _1391 : _425;
    assign _5588 = _1381 == _5597;
    assign _5589 = _1376 & _5588;
    assign _5594 = _5589 ? _1394 : _5593;
    assign _5585 = _299 == _5597;
    assign _5586 = _1376 & _5585;
    assign _5596 = _5586 ? _1099 : _5594;
    assign _5602 = _285 ? _5601 : _5596;
    assign _229 = _5602;
    always @(posedge _277) begin
        if (_275)
            _425 <= _1099;
        else
            _425 <= _229;
    end
    assign _5616 = 8'b00100001;
    assign _5617 = _280 == _5616;
    assign _5620 = _5617 ? _6252 : _1099;
    assign _5610 = _1386 == _5616;
    assign _5611 = _1376 & _5610;
    assign _5612 = _5611 ? _1391 : _422;
    assign _5607 = _1381 == _5616;
    assign _5608 = _1376 & _5607;
    assign _5613 = _5608 ? _1394 : _5612;
    assign _5604 = _299 == _5616;
    assign _5605 = _1376 & _5604;
    assign _5615 = _5605 ? _1099 : _5613;
    assign _5621 = _285 ? _5620 : _5615;
    assign _230 = _5621;
    always @(posedge _277) begin
        if (_275)
            _422 <= _1099;
        else
            _422 <= _230;
    end
    assign _5635 = 8'b00100000;
    assign _5636 = _280 == _5635;
    assign _5639 = _5636 ? _6252 : _1099;
    assign _5629 = _1386 == _5635;
    assign _5630 = _1376 & _5629;
    assign _5631 = _5630 ? _1391 : _419;
    assign _5626 = _1381 == _5635;
    assign _5627 = _1376 & _5626;
    assign _5632 = _5627 ? _1394 : _5631;
    assign _5623 = _299 == _5635;
    assign _5624 = _1376 & _5623;
    assign _5634 = _5624 ? _1099 : _5632;
    assign _5640 = _285 ? _5639 : _5634;
    assign _231 = _5640;
    always @(posedge _277) begin
        if (_275)
            _419 <= _1099;
        else
            _419 <= _231;
    end
    assign _5654 = 8'b00011111;
    assign _5655 = _280 == _5654;
    assign _5658 = _5655 ? _6252 : _1099;
    assign _5648 = _1386 == _5654;
    assign _5649 = _1376 & _5648;
    assign _5650 = _5649 ? _1391 : _416;
    assign _5645 = _1381 == _5654;
    assign _5646 = _1376 & _5645;
    assign _5651 = _5646 ? _1394 : _5650;
    assign _5642 = _299 == _5654;
    assign _5643 = _1376 & _5642;
    assign _5653 = _5643 ? _1099 : _5651;
    assign _5659 = _285 ? _5658 : _5653;
    assign _232 = _5659;
    always @(posedge _277) begin
        if (_275)
            _416 <= _1099;
        else
            _416 <= _232;
    end
    assign _5673 = 8'b00011110;
    assign _5674 = _280 == _5673;
    assign _5677 = _5674 ? _6252 : _1099;
    assign _5667 = _1386 == _5673;
    assign _5668 = _1376 & _5667;
    assign _5669 = _5668 ? _1391 : _413;
    assign _5664 = _1381 == _5673;
    assign _5665 = _1376 & _5664;
    assign _5670 = _5665 ? _1394 : _5669;
    assign _5661 = _299 == _5673;
    assign _5662 = _1376 & _5661;
    assign _5672 = _5662 ? _1099 : _5670;
    assign _5678 = _285 ? _5677 : _5672;
    assign _233 = _5678;
    always @(posedge _277) begin
        if (_275)
            _413 <= _1099;
        else
            _413 <= _233;
    end
    assign _5692 = 8'b00011101;
    assign _5693 = _280 == _5692;
    assign _5696 = _5693 ? _6252 : _1099;
    assign _5686 = _1386 == _5692;
    assign _5687 = _1376 & _5686;
    assign _5688 = _5687 ? _1391 : _410;
    assign _5683 = _1381 == _5692;
    assign _5684 = _1376 & _5683;
    assign _5689 = _5684 ? _1394 : _5688;
    assign _5680 = _299 == _5692;
    assign _5681 = _1376 & _5680;
    assign _5691 = _5681 ? _1099 : _5689;
    assign _5697 = _285 ? _5696 : _5691;
    assign _234 = _5697;
    always @(posedge _277) begin
        if (_275)
            _410 <= _1099;
        else
            _410 <= _234;
    end
    assign _5711 = 8'b00011100;
    assign _5712 = _280 == _5711;
    assign _5715 = _5712 ? _6252 : _1099;
    assign _5705 = _1386 == _5711;
    assign _5706 = _1376 & _5705;
    assign _5707 = _5706 ? _1391 : _407;
    assign _5702 = _1381 == _5711;
    assign _5703 = _1376 & _5702;
    assign _5708 = _5703 ? _1394 : _5707;
    assign _5699 = _299 == _5711;
    assign _5700 = _1376 & _5699;
    assign _5710 = _5700 ? _1099 : _5708;
    assign _5716 = _285 ? _5715 : _5710;
    assign _235 = _5716;
    always @(posedge _277) begin
        if (_275)
            _407 <= _1099;
        else
            _407 <= _235;
    end
    assign _5730 = 8'b00011011;
    assign _5731 = _280 == _5730;
    assign _5734 = _5731 ? _6252 : _1099;
    assign _5724 = _1386 == _5730;
    assign _5725 = _1376 & _5724;
    assign _5726 = _5725 ? _1391 : _404;
    assign _5721 = _1381 == _5730;
    assign _5722 = _1376 & _5721;
    assign _5727 = _5722 ? _1394 : _5726;
    assign _5718 = _299 == _5730;
    assign _5719 = _1376 & _5718;
    assign _5729 = _5719 ? _1099 : _5727;
    assign _5735 = _285 ? _5734 : _5729;
    assign _236 = _5735;
    always @(posedge _277) begin
        if (_275)
            _404 <= _1099;
        else
            _404 <= _236;
    end
    assign _5749 = 8'b00011010;
    assign _5750 = _280 == _5749;
    assign _5753 = _5750 ? _6252 : _1099;
    assign _5743 = _1386 == _5749;
    assign _5744 = _1376 & _5743;
    assign _5745 = _5744 ? _1391 : _401;
    assign _5740 = _1381 == _5749;
    assign _5741 = _1376 & _5740;
    assign _5746 = _5741 ? _1394 : _5745;
    assign _5737 = _299 == _5749;
    assign _5738 = _1376 & _5737;
    assign _5748 = _5738 ? _1099 : _5746;
    assign _5754 = _285 ? _5753 : _5748;
    assign _237 = _5754;
    always @(posedge _277) begin
        if (_275)
            _401 <= _1099;
        else
            _401 <= _237;
    end
    assign _5768 = 8'b00011001;
    assign _5769 = _280 == _5768;
    assign _5772 = _5769 ? _6252 : _1099;
    assign _5762 = _1386 == _5768;
    assign _5763 = _1376 & _5762;
    assign _5764 = _5763 ? _1391 : _398;
    assign _5759 = _1381 == _5768;
    assign _5760 = _1376 & _5759;
    assign _5765 = _5760 ? _1394 : _5764;
    assign _5756 = _299 == _5768;
    assign _5757 = _1376 & _5756;
    assign _5767 = _5757 ? _1099 : _5765;
    assign _5773 = _285 ? _5772 : _5767;
    assign _238 = _5773;
    always @(posedge _277) begin
        if (_275)
            _398 <= _1099;
        else
            _398 <= _238;
    end
    assign _5787 = 8'b00011000;
    assign _5788 = _280 == _5787;
    assign _5791 = _5788 ? _6252 : _1099;
    assign _5781 = _1386 == _5787;
    assign _5782 = _1376 & _5781;
    assign _5783 = _5782 ? _1391 : _395;
    assign _5778 = _1381 == _5787;
    assign _5779 = _1376 & _5778;
    assign _5784 = _5779 ? _1394 : _5783;
    assign _5775 = _299 == _5787;
    assign _5776 = _1376 & _5775;
    assign _5786 = _5776 ? _1099 : _5784;
    assign _5792 = _285 ? _5791 : _5786;
    assign _239 = _5792;
    always @(posedge _277) begin
        if (_275)
            _395 <= _1099;
        else
            _395 <= _239;
    end
    assign _5806 = 8'b00010111;
    assign _5807 = _280 == _5806;
    assign _5810 = _5807 ? _6252 : _1099;
    assign _5800 = _1386 == _5806;
    assign _5801 = _1376 & _5800;
    assign _5802 = _5801 ? _1391 : _392;
    assign _5797 = _1381 == _5806;
    assign _5798 = _1376 & _5797;
    assign _5803 = _5798 ? _1394 : _5802;
    assign _5794 = _299 == _5806;
    assign _5795 = _1376 & _5794;
    assign _5805 = _5795 ? _1099 : _5803;
    assign _5811 = _285 ? _5810 : _5805;
    assign _240 = _5811;
    always @(posedge _277) begin
        if (_275)
            _392 <= _1099;
        else
            _392 <= _240;
    end
    assign _5825 = 8'b00010110;
    assign _5826 = _280 == _5825;
    assign _5829 = _5826 ? _6252 : _1099;
    assign _5819 = _1386 == _5825;
    assign _5820 = _1376 & _5819;
    assign _5821 = _5820 ? _1391 : _389;
    assign _5816 = _1381 == _5825;
    assign _5817 = _1376 & _5816;
    assign _5822 = _5817 ? _1394 : _5821;
    assign _5813 = _299 == _5825;
    assign _5814 = _1376 & _5813;
    assign _5824 = _5814 ? _1099 : _5822;
    assign _5830 = _285 ? _5829 : _5824;
    assign _241 = _5830;
    always @(posedge _277) begin
        if (_275)
            _389 <= _1099;
        else
            _389 <= _241;
    end
    assign _5844 = 8'b00010101;
    assign _5845 = _280 == _5844;
    assign _5848 = _5845 ? _6252 : _1099;
    assign _5838 = _1386 == _5844;
    assign _5839 = _1376 & _5838;
    assign _5840 = _5839 ? _1391 : _386;
    assign _5835 = _1381 == _5844;
    assign _5836 = _1376 & _5835;
    assign _5841 = _5836 ? _1394 : _5840;
    assign _5832 = _299 == _5844;
    assign _5833 = _1376 & _5832;
    assign _5843 = _5833 ? _1099 : _5841;
    assign _5849 = _285 ? _5848 : _5843;
    assign _242 = _5849;
    always @(posedge _277) begin
        if (_275)
            _386 <= _1099;
        else
            _386 <= _242;
    end
    assign _5863 = 8'b00010100;
    assign _5864 = _280 == _5863;
    assign _5867 = _5864 ? _6252 : _1099;
    assign _5857 = _1386 == _5863;
    assign _5858 = _1376 & _5857;
    assign _5859 = _5858 ? _1391 : _383;
    assign _5854 = _1381 == _5863;
    assign _5855 = _1376 & _5854;
    assign _5860 = _5855 ? _1394 : _5859;
    assign _5851 = _299 == _5863;
    assign _5852 = _1376 & _5851;
    assign _5862 = _5852 ? _1099 : _5860;
    assign _5868 = _285 ? _5867 : _5862;
    assign _243 = _5868;
    always @(posedge _277) begin
        if (_275)
            _383 <= _1099;
        else
            _383 <= _243;
    end
    assign _5882 = 8'b00010011;
    assign _5883 = _280 == _5882;
    assign _5886 = _5883 ? _6252 : _1099;
    assign _5876 = _1386 == _5882;
    assign _5877 = _1376 & _5876;
    assign _5878 = _5877 ? _1391 : _380;
    assign _5873 = _1381 == _5882;
    assign _5874 = _1376 & _5873;
    assign _5879 = _5874 ? _1394 : _5878;
    assign _5870 = _299 == _5882;
    assign _5871 = _1376 & _5870;
    assign _5881 = _5871 ? _1099 : _5879;
    assign _5887 = _285 ? _5886 : _5881;
    assign _244 = _5887;
    always @(posedge _277) begin
        if (_275)
            _380 <= _1099;
        else
            _380 <= _244;
    end
    assign _5901 = 8'b00010010;
    assign _5902 = _280 == _5901;
    assign _5905 = _5902 ? _6252 : _1099;
    assign _5895 = _1386 == _5901;
    assign _5896 = _1376 & _5895;
    assign _5897 = _5896 ? _1391 : _377;
    assign _5892 = _1381 == _5901;
    assign _5893 = _1376 & _5892;
    assign _5898 = _5893 ? _1394 : _5897;
    assign _5889 = _299 == _5901;
    assign _5890 = _1376 & _5889;
    assign _5900 = _5890 ? _1099 : _5898;
    assign _5906 = _285 ? _5905 : _5900;
    assign _245 = _5906;
    always @(posedge _277) begin
        if (_275)
            _377 <= _1099;
        else
            _377 <= _245;
    end
    assign _5920 = 8'b00010001;
    assign _5921 = _280 == _5920;
    assign _5924 = _5921 ? _6252 : _1099;
    assign _5914 = _1386 == _5920;
    assign _5915 = _1376 & _5914;
    assign _5916 = _5915 ? _1391 : _374;
    assign _5911 = _1381 == _5920;
    assign _5912 = _1376 & _5911;
    assign _5917 = _5912 ? _1394 : _5916;
    assign _5908 = _299 == _5920;
    assign _5909 = _1376 & _5908;
    assign _5919 = _5909 ? _1099 : _5917;
    assign _5925 = _285 ? _5924 : _5919;
    assign _246 = _5925;
    always @(posedge _277) begin
        if (_275)
            _374 <= _1099;
        else
            _374 <= _246;
    end
    assign _5939 = 8'b00010000;
    assign _5940 = _280 == _5939;
    assign _5943 = _5940 ? _6252 : _1099;
    assign _5933 = _1386 == _5939;
    assign _5934 = _1376 & _5933;
    assign _5935 = _5934 ? _1391 : _371;
    assign _5930 = _1381 == _5939;
    assign _5931 = _1376 & _5930;
    assign _5936 = _5931 ? _1394 : _5935;
    assign _5927 = _299 == _5939;
    assign _5928 = _1376 & _5927;
    assign _5938 = _5928 ? _1099 : _5936;
    assign _5944 = _285 ? _5943 : _5938;
    assign _247 = _5944;
    always @(posedge _277) begin
        if (_275)
            _371 <= _1099;
        else
            _371 <= _247;
    end
    assign _5958 = 8'b00001111;
    assign _5959 = _280 == _5958;
    assign _5962 = _5959 ? _6252 : _1099;
    assign _5952 = _1386 == _5958;
    assign _5953 = _1376 & _5952;
    assign _5954 = _5953 ? _1391 : _368;
    assign _5949 = _1381 == _5958;
    assign _5950 = _1376 & _5949;
    assign _5955 = _5950 ? _1394 : _5954;
    assign _5946 = _299 == _5958;
    assign _5947 = _1376 & _5946;
    assign _5957 = _5947 ? _1099 : _5955;
    assign _5963 = _285 ? _5962 : _5957;
    assign _248 = _5963;
    always @(posedge _277) begin
        if (_275)
            _368 <= _1099;
        else
            _368 <= _248;
    end
    assign _5977 = 8'b00001110;
    assign _5978 = _280 == _5977;
    assign _5981 = _5978 ? _6252 : _1099;
    assign _5971 = _1386 == _5977;
    assign _5972 = _1376 & _5971;
    assign _5973 = _5972 ? _1391 : _365;
    assign _5968 = _1381 == _5977;
    assign _5969 = _1376 & _5968;
    assign _5974 = _5969 ? _1394 : _5973;
    assign _5965 = _299 == _5977;
    assign _5966 = _1376 & _5965;
    assign _5976 = _5966 ? _1099 : _5974;
    assign _5982 = _285 ? _5981 : _5976;
    assign _249 = _5982;
    always @(posedge _277) begin
        if (_275)
            _365 <= _1099;
        else
            _365 <= _249;
    end
    assign _5996 = 8'b00001101;
    assign _5997 = _280 == _5996;
    assign _6000 = _5997 ? _6252 : _1099;
    assign _5990 = _1386 == _5996;
    assign _5991 = _1376 & _5990;
    assign _5992 = _5991 ? _1391 : _362;
    assign _5987 = _1381 == _5996;
    assign _5988 = _1376 & _5987;
    assign _5993 = _5988 ? _1394 : _5992;
    assign _5984 = _299 == _5996;
    assign _5985 = _1376 & _5984;
    assign _5995 = _5985 ? _1099 : _5993;
    assign _6001 = _285 ? _6000 : _5995;
    assign _250 = _6001;
    always @(posedge _277) begin
        if (_275)
            _362 <= _1099;
        else
            _362 <= _250;
    end
    assign _6015 = 8'b00001100;
    assign _6016 = _280 == _6015;
    assign _6019 = _6016 ? _6252 : _1099;
    assign _6009 = _1386 == _6015;
    assign _6010 = _1376 & _6009;
    assign _6011 = _6010 ? _1391 : _359;
    assign _6006 = _1381 == _6015;
    assign _6007 = _1376 & _6006;
    assign _6012 = _6007 ? _1394 : _6011;
    assign _6003 = _299 == _6015;
    assign _6004 = _1376 & _6003;
    assign _6014 = _6004 ? _1099 : _6012;
    assign _6020 = _285 ? _6019 : _6014;
    assign _251 = _6020;
    always @(posedge _277) begin
        if (_275)
            _359 <= _1099;
        else
            _359 <= _251;
    end
    assign _6034 = 8'b00001011;
    assign _6035 = _280 == _6034;
    assign _6038 = _6035 ? _6252 : _1099;
    assign _6028 = _1386 == _6034;
    assign _6029 = _1376 & _6028;
    assign _6030 = _6029 ? _1391 : _356;
    assign _6025 = _1381 == _6034;
    assign _6026 = _1376 & _6025;
    assign _6031 = _6026 ? _1394 : _6030;
    assign _6022 = _299 == _6034;
    assign _6023 = _1376 & _6022;
    assign _6033 = _6023 ? _1099 : _6031;
    assign _6039 = _285 ? _6038 : _6033;
    assign _252 = _6039;
    always @(posedge _277) begin
        if (_275)
            _356 <= _1099;
        else
            _356 <= _252;
    end
    assign _6053 = 8'b00001010;
    assign _6054 = _280 == _6053;
    assign _6057 = _6054 ? _6252 : _1099;
    assign _6047 = _1386 == _6053;
    assign _6048 = _1376 & _6047;
    assign _6049 = _6048 ? _1391 : _353;
    assign _6044 = _1381 == _6053;
    assign _6045 = _1376 & _6044;
    assign _6050 = _6045 ? _1394 : _6049;
    assign _6041 = _299 == _6053;
    assign _6042 = _1376 & _6041;
    assign _6052 = _6042 ? _1099 : _6050;
    assign _6058 = _285 ? _6057 : _6052;
    assign _253 = _6058;
    always @(posedge _277) begin
        if (_275)
            _353 <= _1099;
        else
            _353 <= _253;
    end
    assign _6072 = 8'b00001001;
    assign _6073 = _280 == _6072;
    assign _6076 = _6073 ? _6252 : _1099;
    assign _6066 = _1386 == _6072;
    assign _6067 = _1376 & _6066;
    assign _6068 = _6067 ? _1391 : _350;
    assign _6063 = _1381 == _6072;
    assign _6064 = _1376 & _6063;
    assign _6069 = _6064 ? _1394 : _6068;
    assign _6060 = _299 == _6072;
    assign _6061 = _1376 & _6060;
    assign _6071 = _6061 ? _1099 : _6069;
    assign _6077 = _285 ? _6076 : _6071;
    assign _254 = _6077;
    always @(posedge _277) begin
        if (_275)
            _350 <= _1099;
        else
            _350 <= _254;
    end
    assign _6091 = 8'b00001000;
    assign _6092 = _280 == _6091;
    assign _6095 = _6092 ? _6252 : _1099;
    assign _6085 = _1386 == _6091;
    assign _6086 = _1376 & _6085;
    assign _6087 = _6086 ? _1391 : _347;
    assign _6082 = _1381 == _6091;
    assign _6083 = _1376 & _6082;
    assign _6088 = _6083 ? _1394 : _6087;
    assign _6079 = _299 == _6091;
    assign _6080 = _1376 & _6079;
    assign _6090 = _6080 ? _1099 : _6088;
    assign _6096 = _285 ? _6095 : _6090;
    assign _255 = _6096;
    always @(posedge _277) begin
        if (_275)
            _347 <= _1099;
        else
            _347 <= _255;
    end
    assign _6110 = 8'b00000111;
    assign _6111 = _280 == _6110;
    assign _6114 = _6111 ? _6252 : _1099;
    assign _6104 = _1386 == _6110;
    assign _6105 = _1376 & _6104;
    assign _6106 = _6105 ? _1391 : _344;
    assign _6101 = _1381 == _6110;
    assign _6102 = _1376 & _6101;
    assign _6107 = _6102 ? _1394 : _6106;
    assign _6098 = _299 == _6110;
    assign _6099 = _1376 & _6098;
    assign _6109 = _6099 ? _1099 : _6107;
    assign _6115 = _285 ? _6114 : _6109;
    assign _256 = _6115;
    always @(posedge _277) begin
        if (_275)
            _344 <= _1099;
        else
            _344 <= _256;
    end
    assign _6129 = 8'b00000110;
    assign _6130 = _280 == _6129;
    assign _6133 = _6130 ? _6252 : _1099;
    assign _6123 = _1386 == _6129;
    assign _6124 = _1376 & _6123;
    assign _6125 = _6124 ? _1391 : _341;
    assign _6120 = _1381 == _6129;
    assign _6121 = _1376 & _6120;
    assign _6126 = _6121 ? _1394 : _6125;
    assign _6117 = _299 == _6129;
    assign _6118 = _1376 & _6117;
    assign _6128 = _6118 ? _1099 : _6126;
    assign _6134 = _285 ? _6133 : _6128;
    assign _257 = _6134;
    always @(posedge _277) begin
        if (_275)
            _341 <= _1099;
        else
            _341 <= _257;
    end
    assign _6148 = 8'b00000101;
    assign _6149 = _280 == _6148;
    assign _6152 = _6149 ? _6252 : _1099;
    assign _6142 = _1386 == _6148;
    assign _6143 = _1376 & _6142;
    assign _6144 = _6143 ? _1391 : _338;
    assign _6139 = _1381 == _6148;
    assign _6140 = _1376 & _6139;
    assign _6145 = _6140 ? _1394 : _6144;
    assign _6136 = _299 == _6148;
    assign _6137 = _1376 & _6136;
    assign _6147 = _6137 ? _1099 : _6145;
    assign _6153 = _285 ? _6152 : _6147;
    assign _258 = _6153;
    always @(posedge _277) begin
        if (_275)
            _338 <= _1099;
        else
            _338 <= _258;
    end
    assign _6167 = 8'b00000100;
    assign _6168 = _280 == _6167;
    assign _6171 = _6168 ? _6252 : _1099;
    assign _6161 = _1386 == _6167;
    assign _6162 = _1376 & _6161;
    assign _6163 = _6162 ? _1391 : _335;
    assign _6158 = _1381 == _6167;
    assign _6159 = _1376 & _6158;
    assign _6164 = _6159 ? _1394 : _6163;
    assign _6155 = _299 == _6167;
    assign _6156 = _1376 & _6155;
    assign _6166 = _6156 ? _1099 : _6164;
    assign _6172 = _285 ? _6171 : _6166;
    assign _259 = _6172;
    always @(posedge _277) begin
        if (_275)
            _335 <= _1099;
        else
            _335 <= _259;
    end
    assign _6186 = 8'b00000011;
    assign _6187 = _280 == _6186;
    assign _6190 = _6187 ? _6252 : _1099;
    assign _6180 = _1386 == _6186;
    assign _6181 = _1376 & _6180;
    assign _6182 = _6181 ? _1391 : _332;
    assign _6177 = _1381 == _6186;
    assign _6178 = _1376 & _6177;
    assign _6183 = _6178 ? _1394 : _6182;
    assign _6174 = _299 == _6186;
    assign _6175 = _1376 & _6174;
    assign _6185 = _6175 ? _1099 : _6183;
    assign _6191 = _285 ? _6190 : _6185;
    assign _260 = _6191;
    always @(posedge _277) begin
        if (_275)
            _332 <= _1099;
        else
            _332 <= _260;
    end
    assign _6205 = 8'b00000010;
    assign _6206 = _280 == _6205;
    assign _6209 = _6206 ? _6252 : _1099;
    assign _6199 = _1386 == _6205;
    assign _6200 = _1376 & _6199;
    assign _6201 = _6200 ? _1391 : _329;
    assign _6196 = _1381 == _6205;
    assign _6197 = _1376 & _6196;
    assign _6202 = _6197 ? _1394 : _6201;
    assign _6193 = _299 == _6205;
    assign _6194 = _1376 & _6193;
    assign _6204 = _6194 ? _1099 : _6202;
    assign _6210 = _285 ? _6209 : _6204;
    assign _261 = _6210;
    always @(posedge _277) begin
        if (_275)
            _329 <= _1099;
        else
            _329 <= _261;
    end
    always @* begin
        case (_1381)
        0:
            _1393 <= _323;
        1:
            _1393 <= _326;
        2:
            _1393 <= _329;
        3:
            _1393 <= _332;
        4:
            _1393 <= _335;
        5:
            _1393 <= _338;
        6:
            _1393 <= _341;
        7:
            _1393 <= _344;
        8:
            _1393 <= _347;
        9:
            _1393 <= _350;
        10:
            _1393 <= _353;
        11:
            _1393 <= _356;
        12:
            _1393 <= _359;
        13:
            _1393 <= _362;
        14:
            _1393 <= _365;
        15:
            _1393 <= _368;
        16:
            _1393 <= _371;
        17:
            _1393 <= _374;
        18:
            _1393 <= _377;
        19:
            _1393 <= _380;
        20:
            _1393 <= _383;
        21:
            _1393 <= _386;
        22:
            _1393 <= _389;
        23:
            _1393 <= _392;
        24:
            _1393 <= _395;
        25:
            _1393 <= _398;
        26:
            _1393 <= _401;
        27:
            _1393 <= _404;
        28:
            _1393 <= _407;
        29:
            _1393 <= _410;
        30:
            _1393 <= _413;
        31:
            _1393 <= _416;
        32:
            _1393 <= _419;
        33:
            _1393 <= _422;
        34:
            _1393 <= _425;
        35:
            _1393 <= _428;
        36:
            _1393 <= _431;
        37:
            _1393 <= _434;
        38:
            _1393 <= _437;
        39:
            _1393 <= _440;
        40:
            _1393 <= _443;
        41:
            _1393 <= _446;
        42:
            _1393 <= _449;
        43:
            _1393 <= _452;
        44:
            _1393 <= _455;
        45:
            _1393 <= _458;
        46:
            _1393 <= _461;
        47:
            _1393 <= _464;
        48:
            _1393 <= _467;
        49:
            _1393 <= _470;
        50:
            _1393 <= _473;
        51:
            _1393 <= _476;
        52:
            _1393 <= _479;
        53:
            _1393 <= _482;
        54:
            _1393 <= _485;
        55:
            _1393 <= _488;
        56:
            _1393 <= _491;
        57:
            _1393 <= _494;
        58:
            _1393 <= _497;
        59:
            _1393 <= _500;
        60:
            _1393 <= _503;
        61:
            _1393 <= _506;
        62:
            _1393 <= _509;
        63:
            _1393 <= _512;
        64:
            _1393 <= _515;
        65:
            _1393 <= _518;
        66:
            _1393 <= _521;
        67:
            _1393 <= _524;
        68:
            _1393 <= _527;
        69:
            _1393 <= _530;
        70:
            _1393 <= _533;
        71:
            _1393 <= _536;
        72:
            _1393 <= _539;
        73:
            _1393 <= _542;
        74:
            _1393 <= _545;
        75:
            _1393 <= _548;
        76:
            _1393 <= _551;
        77:
            _1393 <= _554;
        78:
            _1393 <= _557;
        79:
            _1393 <= _560;
        80:
            _1393 <= _563;
        81:
            _1393 <= _566;
        82:
            _1393 <= _569;
        83:
            _1393 <= _572;
        84:
            _1393 <= _575;
        85:
            _1393 <= _578;
        86:
            _1393 <= _581;
        87:
            _1393 <= _584;
        88:
            _1393 <= _587;
        89:
            _1393 <= _590;
        90:
            _1393 <= _593;
        91:
            _1393 <= _596;
        92:
            _1393 <= _599;
        93:
            _1393 <= _602;
        94:
            _1393 <= _605;
        95:
            _1393 <= _608;
        96:
            _1393 <= _611;
        97:
            _1393 <= _614;
        98:
            _1393 <= _617;
        99:
            _1393 <= _620;
        100:
            _1393 <= _623;
        101:
            _1393 <= _626;
        102:
            _1393 <= _629;
        103:
            _1393 <= _632;
        104:
            _1393 <= _635;
        105:
            _1393 <= _638;
        106:
            _1393 <= _641;
        107:
            _1393 <= _644;
        108:
            _1393 <= _647;
        109:
            _1393 <= _650;
        110:
            _1393 <= _653;
        111:
            _1393 <= _656;
        112:
            _1393 <= _659;
        113:
            _1393 <= _662;
        114:
            _1393 <= _665;
        115:
            _1393 <= _668;
        116:
            _1393 <= _671;
        117:
            _1393 <= _674;
        118:
            _1393 <= _677;
        119:
            _1393 <= _680;
        120:
            _1393 <= _683;
        121:
            _1393 <= _686;
        122:
            _1393 <= _689;
        123:
            _1393 <= _692;
        124:
            _1393 <= _695;
        125:
            _1393 <= _698;
        126:
            _1393 <= _701;
        127:
            _1393 <= _704;
        128:
            _1393 <= _707;
        129:
            _1393 <= _710;
        130:
            _1393 <= _713;
        131:
            _1393 <= _716;
        132:
            _1393 <= _719;
        133:
            _1393 <= _722;
        134:
            _1393 <= _725;
        135:
            _1393 <= _728;
        136:
            _1393 <= _731;
        137:
            _1393 <= _734;
        138:
            _1393 <= _737;
        139:
            _1393 <= _740;
        140:
            _1393 <= _743;
        141:
            _1393 <= _746;
        142:
            _1393 <= _749;
        143:
            _1393 <= _752;
        144:
            _1393 <= _755;
        145:
            _1393 <= _758;
        146:
            _1393 <= _761;
        147:
            _1393 <= _764;
        148:
            _1393 <= _767;
        149:
            _1393 <= _770;
        150:
            _1393 <= _773;
        151:
            _1393 <= _776;
        152:
            _1393 <= _779;
        153:
            _1393 <= _782;
        154:
            _1393 <= _785;
        155:
            _1393 <= _788;
        156:
            _1393 <= _791;
        157:
            _1393 <= _794;
        158:
            _1393 <= _797;
        159:
            _1393 <= _800;
        160:
            _1393 <= _803;
        161:
            _1393 <= _806;
        162:
            _1393 <= _809;
        163:
            _1393 <= _812;
        164:
            _1393 <= _815;
        165:
            _1393 <= _818;
        166:
            _1393 <= _821;
        167:
            _1393 <= _824;
        168:
            _1393 <= _827;
        169:
            _1393 <= _830;
        170:
            _1393 <= _833;
        171:
            _1393 <= _836;
        172:
            _1393 <= _839;
        173:
            _1393 <= _842;
        174:
            _1393 <= _845;
        175:
            _1393 <= _848;
        176:
            _1393 <= _851;
        177:
            _1393 <= _854;
        178:
            _1393 <= _857;
        179:
            _1393 <= _860;
        180:
            _1393 <= _863;
        181:
            _1393 <= _866;
        182:
            _1393 <= _869;
        183:
            _1393 <= _872;
        184:
            _1393 <= _875;
        185:
            _1393 <= _878;
        186:
            _1393 <= _881;
        187:
            _1393 <= _884;
        188:
            _1393 <= _887;
        189:
            _1393 <= _890;
        190:
            _1393 <= _893;
        191:
            _1393 <= _896;
        192:
            _1393 <= _899;
        193:
            _1393 <= _902;
        194:
            _1393 <= _905;
        195:
            _1393 <= _908;
        196:
            _1393 <= _911;
        197:
            _1393 <= _914;
        198:
            _1393 <= _917;
        199:
            _1393 <= _920;
        200:
            _1393 <= _923;
        201:
            _1393 <= _926;
        202:
            _1393 <= _929;
        203:
            _1393 <= _932;
        204:
            _1393 <= _935;
        205:
            _1393 <= _938;
        206:
            _1393 <= _941;
        207:
            _1393 <= _944;
        208:
            _1393 <= _947;
        209:
            _1393 <= _950;
        210:
            _1393 <= _953;
        211:
            _1393 <= _956;
        212:
            _1393 <= _959;
        213:
            _1393 <= _962;
        214:
            _1393 <= _965;
        215:
            _1393 <= _968;
        216:
            _1393 <= _971;
        217:
            _1393 <= _974;
        218:
            _1393 <= _977;
        219:
            _1393 <= _980;
        220:
            _1393 <= _983;
        221:
            _1393 <= _986;
        222:
            _1393 <= _989;
        223:
            _1393 <= _992;
        224:
            _1393 <= _995;
        225:
            _1393 <= _998;
        226:
            _1393 <= _1001;
        227:
            _1393 <= _1004;
        228:
            _1393 <= _1007;
        229:
            _1393 <= _1010;
        230:
            _1393 <= _1013;
        231:
            _1393 <= _1016;
        232:
            _1393 <= _1019;
        233:
            _1393 <= _1022;
        234:
            _1393 <= _1025;
        235:
            _1393 <= _1028;
        236:
            _1393 <= _1031;
        237:
            _1393 <= _1034;
        238:
            _1393 <= _1037;
        239:
            _1393 <= _1040;
        240:
            _1393 <= _1043;
        241:
            _1393 <= _1046;
        242:
            _1393 <= _1049;
        243:
            _1393 <= _1052;
        244:
            _1393 <= _1055;
        245:
            _1393 <= _1058;
        246:
            _1393 <= _1061;
        247:
            _1393 <= _1064;
        248:
            _1393 <= _1067;
        249:
            _1393 <= _1070;
        250:
            _1393 <= _1073;
        251:
            _1393 <= _1076;
        252:
            _1393 <= _1079;
        253:
            _1393 <= _1082;
        254:
            _1393 <= _1085;
        default:
            _1393 <= _1088;
        endcase
    end
    assign _1394 = _1393 + _1114;
    assign _6218 = _1386 == _6224;
    assign _6219 = _1376 & _6218;
    assign _6220 = _6219 ? _1391 : _326;
    assign _6215 = _1381 == _6224;
    assign _6216 = _1376 & _6215;
    assign _6221 = _6216 ? _1394 : _6220;
    assign _6212 = _299 == _6224;
    assign _6213 = _1376 & _6212;
    assign _6223 = _6213 ? _1099 : _6221;
    assign _6229 = _285 ? _6228 : _6223;
    assign _262 = _6229;
    always @(posedge _277) begin
        if (_275)
            _326 <= _1099;
        else
            _326 <= _262;
    end
    always @* begin
        case (_1386)
        0:
            _1390 <= _323;
        1:
            _1390 <= _326;
        2:
            _1390 <= _329;
        3:
            _1390 <= _332;
        4:
            _1390 <= _335;
        5:
            _1390 <= _338;
        6:
            _1390 <= _341;
        7:
            _1390 <= _344;
        8:
            _1390 <= _347;
        9:
            _1390 <= _350;
        10:
            _1390 <= _353;
        11:
            _1390 <= _356;
        12:
            _1390 <= _359;
        13:
            _1390 <= _362;
        14:
            _1390 <= _365;
        15:
            _1390 <= _368;
        16:
            _1390 <= _371;
        17:
            _1390 <= _374;
        18:
            _1390 <= _377;
        19:
            _1390 <= _380;
        20:
            _1390 <= _383;
        21:
            _1390 <= _386;
        22:
            _1390 <= _389;
        23:
            _1390 <= _392;
        24:
            _1390 <= _395;
        25:
            _1390 <= _398;
        26:
            _1390 <= _401;
        27:
            _1390 <= _404;
        28:
            _1390 <= _407;
        29:
            _1390 <= _410;
        30:
            _1390 <= _413;
        31:
            _1390 <= _416;
        32:
            _1390 <= _419;
        33:
            _1390 <= _422;
        34:
            _1390 <= _425;
        35:
            _1390 <= _428;
        36:
            _1390 <= _431;
        37:
            _1390 <= _434;
        38:
            _1390 <= _437;
        39:
            _1390 <= _440;
        40:
            _1390 <= _443;
        41:
            _1390 <= _446;
        42:
            _1390 <= _449;
        43:
            _1390 <= _452;
        44:
            _1390 <= _455;
        45:
            _1390 <= _458;
        46:
            _1390 <= _461;
        47:
            _1390 <= _464;
        48:
            _1390 <= _467;
        49:
            _1390 <= _470;
        50:
            _1390 <= _473;
        51:
            _1390 <= _476;
        52:
            _1390 <= _479;
        53:
            _1390 <= _482;
        54:
            _1390 <= _485;
        55:
            _1390 <= _488;
        56:
            _1390 <= _491;
        57:
            _1390 <= _494;
        58:
            _1390 <= _497;
        59:
            _1390 <= _500;
        60:
            _1390 <= _503;
        61:
            _1390 <= _506;
        62:
            _1390 <= _509;
        63:
            _1390 <= _512;
        64:
            _1390 <= _515;
        65:
            _1390 <= _518;
        66:
            _1390 <= _521;
        67:
            _1390 <= _524;
        68:
            _1390 <= _527;
        69:
            _1390 <= _530;
        70:
            _1390 <= _533;
        71:
            _1390 <= _536;
        72:
            _1390 <= _539;
        73:
            _1390 <= _542;
        74:
            _1390 <= _545;
        75:
            _1390 <= _548;
        76:
            _1390 <= _551;
        77:
            _1390 <= _554;
        78:
            _1390 <= _557;
        79:
            _1390 <= _560;
        80:
            _1390 <= _563;
        81:
            _1390 <= _566;
        82:
            _1390 <= _569;
        83:
            _1390 <= _572;
        84:
            _1390 <= _575;
        85:
            _1390 <= _578;
        86:
            _1390 <= _581;
        87:
            _1390 <= _584;
        88:
            _1390 <= _587;
        89:
            _1390 <= _590;
        90:
            _1390 <= _593;
        91:
            _1390 <= _596;
        92:
            _1390 <= _599;
        93:
            _1390 <= _602;
        94:
            _1390 <= _605;
        95:
            _1390 <= _608;
        96:
            _1390 <= _611;
        97:
            _1390 <= _614;
        98:
            _1390 <= _617;
        99:
            _1390 <= _620;
        100:
            _1390 <= _623;
        101:
            _1390 <= _626;
        102:
            _1390 <= _629;
        103:
            _1390 <= _632;
        104:
            _1390 <= _635;
        105:
            _1390 <= _638;
        106:
            _1390 <= _641;
        107:
            _1390 <= _644;
        108:
            _1390 <= _647;
        109:
            _1390 <= _650;
        110:
            _1390 <= _653;
        111:
            _1390 <= _656;
        112:
            _1390 <= _659;
        113:
            _1390 <= _662;
        114:
            _1390 <= _665;
        115:
            _1390 <= _668;
        116:
            _1390 <= _671;
        117:
            _1390 <= _674;
        118:
            _1390 <= _677;
        119:
            _1390 <= _680;
        120:
            _1390 <= _683;
        121:
            _1390 <= _686;
        122:
            _1390 <= _689;
        123:
            _1390 <= _692;
        124:
            _1390 <= _695;
        125:
            _1390 <= _698;
        126:
            _1390 <= _701;
        127:
            _1390 <= _704;
        128:
            _1390 <= _707;
        129:
            _1390 <= _710;
        130:
            _1390 <= _713;
        131:
            _1390 <= _716;
        132:
            _1390 <= _719;
        133:
            _1390 <= _722;
        134:
            _1390 <= _725;
        135:
            _1390 <= _728;
        136:
            _1390 <= _731;
        137:
            _1390 <= _734;
        138:
            _1390 <= _737;
        139:
            _1390 <= _740;
        140:
            _1390 <= _743;
        141:
            _1390 <= _746;
        142:
            _1390 <= _749;
        143:
            _1390 <= _752;
        144:
            _1390 <= _755;
        145:
            _1390 <= _758;
        146:
            _1390 <= _761;
        147:
            _1390 <= _764;
        148:
            _1390 <= _767;
        149:
            _1390 <= _770;
        150:
            _1390 <= _773;
        151:
            _1390 <= _776;
        152:
            _1390 <= _779;
        153:
            _1390 <= _782;
        154:
            _1390 <= _785;
        155:
            _1390 <= _788;
        156:
            _1390 <= _791;
        157:
            _1390 <= _794;
        158:
            _1390 <= _797;
        159:
            _1390 <= _800;
        160:
            _1390 <= _803;
        161:
            _1390 <= _806;
        162:
            _1390 <= _809;
        163:
            _1390 <= _812;
        164:
            _1390 <= _815;
        165:
            _1390 <= _818;
        166:
            _1390 <= _821;
        167:
            _1390 <= _824;
        168:
            _1390 <= _827;
        169:
            _1390 <= _830;
        170:
            _1390 <= _833;
        171:
            _1390 <= _836;
        172:
            _1390 <= _839;
        173:
            _1390 <= _842;
        174:
            _1390 <= _845;
        175:
            _1390 <= _848;
        176:
            _1390 <= _851;
        177:
            _1390 <= _854;
        178:
            _1390 <= _857;
        179:
            _1390 <= _860;
        180:
            _1390 <= _863;
        181:
            _1390 <= _866;
        182:
            _1390 <= _869;
        183:
            _1390 <= _872;
        184:
            _1390 <= _875;
        185:
            _1390 <= _878;
        186:
            _1390 <= _881;
        187:
            _1390 <= _884;
        188:
            _1390 <= _887;
        189:
            _1390 <= _890;
        190:
            _1390 <= _893;
        191:
            _1390 <= _896;
        192:
            _1390 <= _899;
        193:
            _1390 <= _902;
        194:
            _1390 <= _905;
        195:
            _1390 <= _908;
        196:
            _1390 <= _911;
        197:
            _1390 <= _914;
        198:
            _1390 <= _917;
        199:
            _1390 <= _920;
        200:
            _1390 <= _923;
        201:
            _1390 <= _926;
        202:
            _1390 <= _929;
        203:
            _1390 <= _932;
        204:
            _1390 <= _935;
        205:
            _1390 <= _938;
        206:
            _1390 <= _941;
        207:
            _1390 <= _944;
        208:
            _1390 <= _947;
        209:
            _1390 <= _950;
        210:
            _1390 <= _953;
        211:
            _1390 <= _956;
        212:
            _1390 <= _959;
        213:
            _1390 <= _962;
        214:
            _1390 <= _965;
        215:
            _1390 <= _968;
        216:
            _1390 <= _971;
        217:
            _1390 <= _974;
        218:
            _1390 <= _977;
        219:
            _1390 <= _980;
        220:
            _1390 <= _983;
        221:
            _1390 <= _986;
        222:
            _1390 <= _989;
        223:
            _1390 <= _992;
        224:
            _1390 <= _995;
        225:
            _1390 <= _998;
        226:
            _1390 <= _1001;
        227:
            _1390 <= _1004;
        228:
            _1390 <= _1007;
        229:
            _1390 <= _1010;
        230:
            _1390 <= _1013;
        231:
            _1390 <= _1016;
        232:
            _1390 <= _1019;
        233:
            _1390 <= _1022;
        234:
            _1390 <= _1025;
        235:
            _1390 <= _1028;
        236:
            _1390 <= _1031;
        237:
            _1390 <= _1034;
        238:
            _1390 <= _1037;
        239:
            _1390 <= _1040;
        240:
            _1390 <= _1043;
        241:
            _1390 <= _1046;
        242:
            _1390 <= _1049;
        243:
            _1390 <= _1052;
        244:
            _1390 <= _1055;
        245:
            _1390 <= _1058;
        246:
            _1390 <= _1061;
        247:
            _1390 <= _1064;
        248:
            _1390 <= _1067;
        249:
            _1390 <= _1070;
        250:
            _1390 <= _1073;
        251:
            _1390 <= _1076;
        252:
            _1390 <= _1079;
        253:
            _1390 <= _1082;
        254:
            _1390 <= _1085;
        default:
            _1390 <= _1088;
        endcase
    end
    assign _1391 = _1390 + _1114;
    assign _1386 = _299 + _6224;
    assign _6237 = _1386 == _6243;
    assign _6238 = _1376 & _6237;
    assign _6239 = _6238 ? _1391 : _323;
    assign _1381 = _299 - _6224;
    assign _6234 = _1381 == _6243;
    assign _6235 = _1376 & _6234;
    assign _6240 = _6235 ? _1394 : _6239;
    assign _6231 = _299 == _6243;
    assign _6232 = _1376 & _6231;
    assign _6242 = _6232 ? _1099 : _6240;
    assign _6248 = _285 ? _6247 : _6242;
    assign _263 = _6248;
    always @(posedge _277) begin
        if (_275)
            _323 <= _1099;
        else
            _323 <= _263;
    end
    always @* begin
        case (_299)
        0:
            _1114 <= _323;
        1:
            _1114 <= _326;
        2:
            _1114 <= _329;
        3:
            _1114 <= _332;
        4:
            _1114 <= _335;
        5:
            _1114 <= _338;
        6:
            _1114 <= _341;
        7:
            _1114 <= _344;
        8:
            _1114 <= _347;
        9:
            _1114 <= _350;
        10:
            _1114 <= _353;
        11:
            _1114 <= _356;
        12:
            _1114 <= _359;
        13:
            _1114 <= _362;
        14:
            _1114 <= _365;
        15:
            _1114 <= _368;
        16:
            _1114 <= _371;
        17:
            _1114 <= _374;
        18:
            _1114 <= _377;
        19:
            _1114 <= _380;
        20:
            _1114 <= _383;
        21:
            _1114 <= _386;
        22:
            _1114 <= _389;
        23:
            _1114 <= _392;
        24:
            _1114 <= _395;
        25:
            _1114 <= _398;
        26:
            _1114 <= _401;
        27:
            _1114 <= _404;
        28:
            _1114 <= _407;
        29:
            _1114 <= _410;
        30:
            _1114 <= _413;
        31:
            _1114 <= _416;
        32:
            _1114 <= _419;
        33:
            _1114 <= _422;
        34:
            _1114 <= _425;
        35:
            _1114 <= _428;
        36:
            _1114 <= _431;
        37:
            _1114 <= _434;
        38:
            _1114 <= _437;
        39:
            _1114 <= _440;
        40:
            _1114 <= _443;
        41:
            _1114 <= _446;
        42:
            _1114 <= _449;
        43:
            _1114 <= _452;
        44:
            _1114 <= _455;
        45:
            _1114 <= _458;
        46:
            _1114 <= _461;
        47:
            _1114 <= _464;
        48:
            _1114 <= _467;
        49:
            _1114 <= _470;
        50:
            _1114 <= _473;
        51:
            _1114 <= _476;
        52:
            _1114 <= _479;
        53:
            _1114 <= _482;
        54:
            _1114 <= _485;
        55:
            _1114 <= _488;
        56:
            _1114 <= _491;
        57:
            _1114 <= _494;
        58:
            _1114 <= _497;
        59:
            _1114 <= _500;
        60:
            _1114 <= _503;
        61:
            _1114 <= _506;
        62:
            _1114 <= _509;
        63:
            _1114 <= _512;
        64:
            _1114 <= _515;
        65:
            _1114 <= _518;
        66:
            _1114 <= _521;
        67:
            _1114 <= _524;
        68:
            _1114 <= _527;
        69:
            _1114 <= _530;
        70:
            _1114 <= _533;
        71:
            _1114 <= _536;
        72:
            _1114 <= _539;
        73:
            _1114 <= _542;
        74:
            _1114 <= _545;
        75:
            _1114 <= _548;
        76:
            _1114 <= _551;
        77:
            _1114 <= _554;
        78:
            _1114 <= _557;
        79:
            _1114 <= _560;
        80:
            _1114 <= _563;
        81:
            _1114 <= _566;
        82:
            _1114 <= _569;
        83:
            _1114 <= _572;
        84:
            _1114 <= _575;
        85:
            _1114 <= _578;
        86:
            _1114 <= _581;
        87:
            _1114 <= _584;
        88:
            _1114 <= _587;
        89:
            _1114 <= _590;
        90:
            _1114 <= _593;
        91:
            _1114 <= _596;
        92:
            _1114 <= _599;
        93:
            _1114 <= _602;
        94:
            _1114 <= _605;
        95:
            _1114 <= _608;
        96:
            _1114 <= _611;
        97:
            _1114 <= _614;
        98:
            _1114 <= _617;
        99:
            _1114 <= _620;
        100:
            _1114 <= _623;
        101:
            _1114 <= _626;
        102:
            _1114 <= _629;
        103:
            _1114 <= _632;
        104:
            _1114 <= _635;
        105:
            _1114 <= _638;
        106:
            _1114 <= _641;
        107:
            _1114 <= _644;
        108:
            _1114 <= _647;
        109:
            _1114 <= _650;
        110:
            _1114 <= _653;
        111:
            _1114 <= _656;
        112:
            _1114 <= _659;
        113:
            _1114 <= _662;
        114:
            _1114 <= _665;
        115:
            _1114 <= _668;
        116:
            _1114 <= _671;
        117:
            _1114 <= _674;
        118:
            _1114 <= _677;
        119:
            _1114 <= _680;
        120:
            _1114 <= _683;
        121:
            _1114 <= _686;
        122:
            _1114 <= _689;
        123:
            _1114 <= _692;
        124:
            _1114 <= _695;
        125:
            _1114 <= _698;
        126:
            _1114 <= _701;
        127:
            _1114 <= _704;
        128:
            _1114 <= _707;
        129:
            _1114 <= _710;
        130:
            _1114 <= _713;
        131:
            _1114 <= _716;
        132:
            _1114 <= _719;
        133:
            _1114 <= _722;
        134:
            _1114 <= _725;
        135:
            _1114 <= _728;
        136:
            _1114 <= _731;
        137:
            _1114 <= _734;
        138:
            _1114 <= _737;
        139:
            _1114 <= _740;
        140:
            _1114 <= _743;
        141:
            _1114 <= _746;
        142:
            _1114 <= _749;
        143:
            _1114 <= _752;
        144:
            _1114 <= _755;
        145:
            _1114 <= _758;
        146:
            _1114 <= _761;
        147:
            _1114 <= _764;
        148:
            _1114 <= _767;
        149:
            _1114 <= _770;
        150:
            _1114 <= _773;
        151:
            _1114 <= _776;
        152:
            _1114 <= _779;
        153:
            _1114 <= _782;
        154:
            _1114 <= _785;
        155:
            _1114 <= _788;
        156:
            _1114 <= _791;
        157:
            _1114 <= _794;
        158:
            _1114 <= _797;
        159:
            _1114 <= _800;
        160:
            _1114 <= _803;
        161:
            _1114 <= _806;
        162:
            _1114 <= _809;
        163:
            _1114 <= _812;
        164:
            _1114 <= _815;
        165:
            _1114 <= _818;
        166:
            _1114 <= _821;
        167:
            _1114 <= _824;
        168:
            _1114 <= _827;
        169:
            _1114 <= _830;
        170:
            _1114 <= _833;
        171:
            _1114 <= _836;
        172:
            _1114 <= _839;
        173:
            _1114 <= _842;
        174:
            _1114 <= _845;
        175:
            _1114 <= _848;
        176:
            _1114 <= _851;
        177:
            _1114 <= _854;
        178:
            _1114 <= _857;
        179:
            _1114 <= _860;
        180:
            _1114 <= _863;
        181:
            _1114 <= _866;
        182:
            _1114 <= _869;
        183:
            _1114 <= _872;
        184:
            _1114 <= _875;
        185:
            _1114 <= _878;
        186:
            _1114 <= _881;
        187:
            _1114 <= _884;
        188:
            _1114 <= _887;
        189:
            _1114 <= _890;
        190:
            _1114 <= _893;
        191:
            _1114 <= _896;
        192:
            _1114 <= _899;
        193:
            _1114 <= _902;
        194:
            _1114 <= _905;
        195:
            _1114 <= _908;
        196:
            _1114 <= _911;
        197:
            _1114 <= _914;
        198:
            _1114 <= _917;
        199:
            _1114 <= _920;
        200:
            _1114 <= _923;
        201:
            _1114 <= _926;
        202:
            _1114 <= _929;
        203:
            _1114 <= _932;
        204:
            _1114 <= _935;
        205:
            _1114 <= _938;
        206:
            _1114 <= _941;
        207:
            _1114 <= _944;
        208:
            _1114 <= _947;
        209:
            _1114 <= _950;
        210:
            _1114 <= _953;
        211:
            _1114 <= _956;
        212:
            _1114 <= _959;
        213:
            _1114 <= _962;
        214:
            _1114 <= _965;
        215:
            _1114 <= _968;
        216:
            _1114 <= _971;
        217:
            _1114 <= _974;
        218:
            _1114 <= _977;
        219:
            _1114 <= _980;
        220:
            _1114 <= _983;
        221:
            _1114 <= _986;
        222:
            _1114 <= _989;
        223:
            _1114 <= _992;
        224:
            _1114 <= _995;
        225:
            _1114 <= _998;
        226:
            _1114 <= _1001;
        227:
            _1114 <= _1004;
        228:
            _1114 <= _1007;
        229:
            _1114 <= _1010;
        230:
            _1114 <= _1013;
        231:
            _1114 <= _1016;
        232:
            _1114 <= _1019;
        233:
            _1114 <= _1022;
        234:
            _1114 <= _1025;
        235:
            _1114 <= _1028;
        236:
            _1114 <= _1031;
        237:
            _1114 <= _1034;
        238:
            _1114 <= _1037;
        239:
            _1114 <= _1040;
        240:
            _1114 <= _1043;
        241:
            _1114 <= _1046;
        242:
            _1114 <= _1049;
        243:
            _1114 <= _1052;
        244:
            _1114 <= _1055;
        245:
            _1114 <= _1058;
        246:
            _1114 <= _1061;
        247:
            _1114 <= _1064;
        248:
            _1114 <= _1067;
        249:
            _1114 <= _1070;
        250:
            _1114 <= _1073;
        251:
            _1114 <= _1076;
        252:
            _1114 <= _1079;
        253:
            _1114 <= _1082;
        254:
            _1114 <= _1085;
        default:
            _1114 <= _1088;
        endcase
    end
    assign _1116 = _1114 == _1099;
    assign _1117 = ~ _1116;
    assign _1113 = _293 & _301;
    assign _1118 = _1113 & _1117;
    assign _1376 = _1118 & _1375;
    assign _6254 = _1376 ? _6253 : _6251;
    assign _6256 = _285 ? _1099 : _6254;
    assign _264 = _6256;
    always @(posedge _277) begin
        if (_275)
            _6251 <= _1099;
        else
            _6251 <= _264;
    end
    assign _6258 = _291 == _6257;
    assign _289 = 3'b000;
    assign _1104 = 3'b001;
    assign _6298 = _306 ? _308 : _1104;
    assign _6257 = 3'b100;
    assign _6259 = _285 ? _279 : _315;
    assign _267 = _6259;
    always @(posedge _277) begin
        if (_275)
            _315 <= _6243;
        else
            _315 <= _267;
    end
    assign _6264 = _312 + _6224;
    assign _6265 = _309 ? _6264 : _312;
    assign _305 = 1'b0;
    assign _269 = row_last;
    assign _6260 = _1106 ? _269 : _306;
    assign _6262 = _285 ? _305 : _6260;
    assign _270 = _6262;
    always @(posedge _277) begin
        if (_275)
            _306 <= _305;
        else
            _306 <= _270;
    end
    assign _307 = _303 & _306;
    assign _6267 = _307 ? _6243 : _6265;
    assign _6269 = _285 ? _6243 : _6267;
    assign _271 = _6269;
    always @(posedge _277) begin
        if (_275)
            _312 <= _6243;
        else
            _312 <= _271;
    end
    assign _316 = _312 < _315;
    assign _1096 = ~ _316;
    assign _308 = 3'b011;
    assign _309 = _291 == _308;
    assign _1097 = _309 & _1096;
    assign _6297 = _1097 ? _6257 : _291;
    assign _6280 = _6276 - _6279;
    assign _6272 = _299 + _6205;
    assign _6270 = _293 & _301;
    assign _6273 = _6270 ? _6272 : _299;
    assign _6281 = _1106 ? _6280 : _6273;
    assign _6283 = _285 ? _6243 : _6281;
    assign _272 = _6283;
    always @(posedge _277) begin
        if (_275)
            _299 <= _6243;
        else
            _299 <= _272;
    end
    assign _6285 = _6279 + _6224;
    assign _6286 = _303 ? _6285 : _6279;
    assign _6288 = _285 ? _6243 : _6286;
    assign _273 = _6288;
    always @(posedge _277) begin
        if (_275)
            _6279 <= _6243;
        else
            _6279 <= _273;
    end
    assign vdd = 1'b1;
    assign _275 = clear;
    assign _277 = clock;
    assign _279 = width;
    assign _6290 = _279[7:1];
    assign _6291 = { _305,
                     _6290 };
    assign _6292 = _285 ? _6291 : _6276;
    assign _280 = _6292;
    always @(posedge _277) begin
        if (_275)
            _6276 <= _6243;
        else
            _6276 <= _280;
    end
    assign _6293 = _6276 + _6279;
    assign _6294 = _1106 ? _6293 : _296;
    assign _6296 = _285 ? _6243 : _6294;
    assign _281 = _6296;
    always @(posedge _277) begin
        if (_275)
            _296 <= _6243;
        else
            _296 <= _281;
    end
    assign _300 = _296 < _299;
    assign _301 = ~ _300;
    assign _302 = ~ _301;
    assign _292 = 3'b010;
    assign _293 = _291 == _292;
    assign _303 = _293 & _302;
    assign _6299 = _303 ? _6298 : _6297;
    assign _283 = row_valid;
    assign _1106 = _1105 & _283;
    assign _6300 = _1106 ? _292 : _6299;
    assign _285 = load;
    assign _6301 = _285 ? _1104 : _6300;
    assign _286 = _6301;
    always @(posedge _277) begin
        if (_275)
            _291 <= _289;
        else
            _291 <= _286;
    end
    assign _1105 = _291 == _1104;
    assign ready = _1105;
    assign done_ = _6258;
    assign part1_result = _6251;
    assign part2_result = _1100;
    assign state = _291;

endmodule
